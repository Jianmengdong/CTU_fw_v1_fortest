

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
TvNAk+dzefmJC5/xfGEoXo1v1zzw15yvf2w3I+7pl9weHnOYLTwk2CtA6qQwUdiv+KPlR09XyHxt
UocEiAlS9g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ccd1Kr3IgmbU3Zd5R5UGhugxe9OUvTTk5M/+YDzRXyTvXIMaUxHB5fv7SuuebIYqGrGlL5seA2Sg
zO1i2uQFXVFn4M1DHS2E7BwirWBP5gmU/RaWKyEfTu3E5ZGbc1lvK67CCG8szRwdrvmY+Z8CpiC4
+fKoXg6GREReZgylTmE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
D4OySXRBGdK3bWTwoBJnna9JJTCfjtow8OCB97TMc0CHJtgWscKG0sA6JP+WmQu+g/St8V3dnWCm
Z/oL2u8esW79WhsyQGAkuc2zUGutMTiH5JtlsxfFXreCjsbpfiQ4cOTSVV8RKFLaZCW+eXj7qQwk
WUd+Rk2Kp6kViZmb9GfGDSBc1qKbMuYuGLGiO+UVYNdt7dkYg9aAhJYx3c/Tx4m6BAZTpzEs9xzl
Mg0Plk7PRG/v5PXojT+9MvJ80iSqd3ejpG6kEE1mYBAhD1zmHQfbte6ipINFibjTuluuS5i0pIbf
HaA/nmULSj1xFBTfeEdDhm4CrFUWEdYvrJoOhg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YmbWYAZhC3ayB3FdtHMbSkvV5OWWIi6gmohNfeiL3hZEqSlPd2B43zehv3FM2BA2v3N0HlGO0TL6
neUbRccVG37R0aVoXEjetzHP+ZMpVpr2wNRYoVv9EAzvD7YjPAyiMQMLJO1wmw/LJVkGpP4UCg4g
tgMS7M+LmVgeot1Fmcwa4mDyquYpShDC0ZhYtWL3VmO204ubc1HcI1fEQiMp+tBP7rYU0jIyGMtz
dXGUYS7PdIYkz5ApCjSfCCueqmWeZf9/KXMkoo9udSh2ZyT9uNr+GM8fH8rcz5nZjN4ShPghIUSN
XIZbR6KJ/+WqugC6B6ULpEZUxft3AS1vxij4dA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pRgO0aX5waanQk0eZ4W7Q+LVxiXC+tf9hFRN9nsdM6xbA9apyUI0wd0pRjkzt/X5yvazLViQDSfS
Bm9cP+mYh23I891gOC2bMeto93RQUYlDhWmKA2HAuokJj6wKo/vk9LA0e/rAjHMWD7cTXHkdXPdz
d92x8sSRX6Z5gz0YOJ8hU+X3aLkMrr/d+Rs3UcELF+MTGSf53SzTuIbnaw08EsHUObyFusQxXlt6
ZuByaRiPP1ofEvMk+UCLRZThOA7sR6SIfjXOTF55TQgss4/Mf30sm+t84LW+xNBWIqVfiQ671PZF
CQ8K4qBj3nTT9D0FTUvfHdTmLtywWgV65+5W3A==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
d38DScsESf/yIfST5KEEwSUvjI+Km/dbua2xenGdzq3rgc/diAWKNIN11lcJIPDVBe6fB9J2TqbT
eXC+WnYP2YB9QXYlwKxLW7HOYcLC6Ivx9uoTg503B1azg5yB52W8iAwxelCieuRZ3qo4CxwOJ4w3
kwV+F675PsE0hWvEwTA=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Bf4H+OH1vHHXYQ0B+xvr52Pkbk3t9R17gzpbDdSPXjerF+p1mOwTJrxL3jQRkm9rUtVIgJGiq2/s
crniU3gwf/UiAzOrNxcIp9eKlLwDNsxSMYn+mkUQWlDdifqNNVK+YFJD0ZFE6pzyWAfSd99uwvf2
B/+VXkZFAWz3devN4zOqXGE5+OZKTJNNH2fm+gcI0n7V4lPByrga5xMdlx99MQZZRprmMts+yOHQ
eVL2q0jneXaC7j4j8aSjRtpPAjf6aWk9xkdj2iVGAqs6TlpdNPyA9bKumNf3XCjAnjbNwxHWWAao
tHbBrxiXF1qQUoAzJ9mjy31tCjRX+JQOzKafLw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967856)
`protect data_block
n1T0pdpdBe+K9m76BbkbTkR2VwoSYeK2S7jkOqOMao1KdXJ62rgqV67iHxgdsXwpKYW6jCiQtvjF
+jPHQzE3PI+vqY8+MrsKqHfMOETXZA5QBu8mCr/3NTeLiuD2Fw7R2erxyw8k+JL4Flc9H+sLKnUT
FkM8+5WYr3wNDJH3qMXqUF8XLj9yh8KgkzJ9xKCWweRnJCk8I//GByfXNVoD6F1S9uEQ7SqCOnau
fWrVNiKmL2JP8rZ1Il2ulWNjOZSvGE9foLirF5/GH0MFCBo0BZZ5czZtOYme8oOcNM6h7njEKuZD
FC4oesDCl8JhsUYKpFMLgdwhcOdLPjDR4bcuvv9A5NfW6KA/xVfp/EG0GAgA1ScpSRhaZxYApby5
7IRyFyM4y+zRGssmPv4eoUhBFGXlxOaFlIQLz7tbqu/bSHTXBk5otWInlLSD0f/aaysq551RwVdm
3QDFAKN89B7uY1SLnxlLIRpIJNfsWPoqXDCwxSOAFLek00foaMdAB1LXdQUeMizT4bEYSjtzVw2J
+Qt2h79ZXT4m492BK4JcJGNf7Sx6AMJYK546ptbzDrvUGsKHdXRP2VtCWg38ruTGyJA+sDY4lQ+D
WB9fnAkwEQaAONx3zVf0L4TiyJEg0Jroo+oD55erOKmluLZwQwaixsoIBGDagjZFZaNDr6WiEOp6
55pRYniwxLQkbNKYS6nmKbEXgW0HuQ3ZeyBKCgMFht807u9WA/ObDS/Lz3AJreJVl4k1fkuL6eJW
us+4MjnlfPzJV1wha/15TkIaMefef3KsfGiNQzf+8dVCW6QXD6MmOF61il2+PIwbTkQx8QQjEtol
mjouYFlH/xD9XsSx2dq5MmePDUb1HYmuqHWkA1POMk0+HjLW+4R+2v0tDDrs+oaWCgbiOupBYhXW
/aLd//8Gcce9sk7fC3S0VWBO+wKc/683viKfyxEZqh2//68wyZbwfldUftjsftGCz70m1OnwLnNj
PGiy1eAA6vEx/BOBrrTWNeTjZlm4nvTuRGE/XVO53ZG8g12DMh06pB2bjCUehFNxwPtKEprFqa+T
Wv5y/1cUn6WhwqK7NVdCUxhY5l/09jGnvXMnZJhWux4yV0iuBUBbsJHIQ2IbNedM/MpXalEfgtXh
IdR1mIwDBRzXUz2oHeuTKbLqd4OCIOBIB5eediSB3UvPEArif0Iq7tX/k7yPUHezBs8n2S1q3Xg1
/0THFxE/XigEcDhlcWeXxVvHh9UFq9yrVZZeY7I+aaSnRDGqgUjGbzZ2spJTgB1bOJZ6u1cVBHwo
TGjsDptsimBXrSAiJnIs8b+MQ/k2ggt0G0+tM+rdPiY9nxXcKVbVLvFAtfAcsGiGTvJjidtYOr8m
rtxEhbx/prtQRtapUJgTCOu8tsFN1PFUwPfK6XI3lfwqi8HqTJrJqmGPXozlHYzdKIN2CvMlUJ3Z
RNsuKcCGnl6ccTngW+UdXGqV6StvuYox37NpKi+7XI0GP5WrXh8AAis7tK6reLlvAGFj4Y3vn76F
ef29r0BR7UrDZqFs6TABitVaulXNJGnUAadDsYD1X6lB9kIUpREhS/uCXCdSQPG+kcyoLQRuQx5q
gR4qQ93vFTurmjmIcE5xV8zDJmkTI9BeKeYqRn9c7eywcnMbpQiYXOw4lcDJYMnpJpPcJ3HvOG2q
PfZq/TofVmZAgJPZr4EWh4Jcf3WFKSxqX8abG11lNWLP6uoFvqdbCO2WNobFJZTy6tjah0gKJCXa
SFiAmnJ5emtC8Wqxn1K+9leDA2Rronha/+EQfeZHhkbdINHCLuDwQDmX4j+WF4IZ8fiW/eb5kDpc
12TLXtTjvSJ65Ipw+rnyhR35PgqtG+KxYjWLfaYe5F0/mDFQQEH/Wpp0SntvQGvkEBWTmZDqaRe4
ATDj0o8qZ30bTAAW4HqPN1X2XUxQwq8OaxVVXo9ROzpDcgwVGGEyUy9NHYkZM2BbSe0XiXoYuBSt
61UEygJ/WtH8Qf/RaJcGF4oNF+aTBkO7A3W6d7xDcVFJFxyGV9A+k8+1Eaw+Qsqkqz1zTjThDWe8
G/h6dFniNInCm0yQcEtvRqAJ73m/2I1EjkXFcn2qEyy4lWXBmra/UWJ8wsxiB/jxcKxrtUdcZWRk
2/JVxLvwrDxi9Dp4Q7rPKbyV39EelWXi6vyq6wcc3pEDXV4hXBBCIYLvayi5keiMsm1Gw6eCOZWt
AcGma4Vy96HwFz/y08B54S5ovPoC7+Ko0tRJyfwwpOghR/F7d4zJHzqKqXJ/w52FCUjwjv6aG9CR
hDo4ROYHZZOLAzdRtRvallkZokgxYCtLBYTACihnMnQiEJFTRxsaJi56m1GAKB9HrI3UrZT/sKyC
Z/8OOoSljt8mQpuAI0VDWnpCKRg5zu5f3lla8usPGAVbxDFbRWYnFiyQBPVajyOXB5brYq7NxxfI
t4SuWJUYlxbvcEuXJwvB+1J6UVEWsVQ4nJcLxNUC5IIHUKqw0FoMnDf4kkBWbGaGDg9iS+bKhuy5
OyeOaGFWVZjwHmF0Tag+8Ts0OfeUmgc0PoWesaiiVxWH+uexn6zjIXM1hLyNIcGCy87Lf1zjwH+/
c+PPTwVjgIz1k0j64fd1p5Rk1Zd61qR5S2TBvkJ2IC2ZKsTqnL9gooPeOFW/+O96bIrvNsETaUNl
3RgNd1nd1UKwJWjcIOV6DoOXUW9FM+auGFQs3ea+2W8j9kLDdipxoA06uUfwBfRhONq7wyXsDred
say0b7m82ru9tbuPOxY5xBQWsA6Ajxis38p7aYKogP+98VhwY1v+ZtJ/gJt7iYYYcFOb5x9/vGcw
ukJDLSsYgoevv4zQMkUT+AYwEYiSlCjXIUHrBQ79g5LpDE2m/jANvZ0hgaWKvGJ/ECboC4q8HDbl
gFRJG4O/auLaRlQZhVr1uWLFvY6nBj/YVSkqpXOYjKTLspqfzz8FWwZMCuMLcW2buP0MD6njGDg8
HnixK3cTd0GB7wCi27WATJqdIgJuhoDja1iEPhjBG4xF97A+MsZnR4L4jHQ7WliUhCrEOPFTDwec
E74TjnLD9NThAA8qiy7PuOhzSOJwAy9vLSshb4bWr0kEBuLNyd/23J0UXq/izioH7//7NrXVx/5G
xQdl39fgSu+DUgj1rGAyJxmx5hi3xu0oi4x7Dj5tjHDVkPV43gXgLdPRnE8EdPCuZZw2nLlxEJuk
1eZKvlYE/wr54Ruy0S1+hUFDd2Pi3uQJD63EtUwt0JlOFlTG989BbcSsznJVCfwpHcWYKsAG1Rnt
BwfVmOyD8/YV6zJSkNv1djRdFjbDdNpsz4G9yODZ2uO+qtLVER3lxlANKyMq36dhtDldsYV6QGpv
xUWsLlfU9G71d4IZ2aW49p9xcU8v96M+h36O6+NAdBWskWvGzx+xBDR6h01dpnIyCHGM+f/uRzL+
H2PwwbsZcxC0yhfipt8Y+o8I5bN/PELG5Dq/hL8sFn+13mplPMrzq/THnmO2XyRyA5EMv6uUN+8O
duCToQNPEq86mfWicbK3xZR0Eymf8im1EmdXEfR/6NCEKROhmyV0X12eyB/lxETmSdmsiCS3EfYS
MS1saOY21kR4tLBIY/B7vjSGq/SEuY2l453OVtbQf+kgOkr2/nC60kamYYP0P0EfF/hPRDj1mPZX
Ia2Pwewjt+PkMbSKwEeRGbrsGWG0L0C9uRnFe/5G+XemmcVvezrt3okBDq58NM+ZJsTB89hg170g
SQLC2ko6DJltRCguDdCoIM6fJ5e7KlbNlRS+7lXiOXtGgAr8aHVqt7ECnMWbI1Cf2kvVPiQlK0KO
r234eodKUo5MwxJ/7eKui+U0JnKwHdPD4AxflqtpWyOJfim/pezgLaouQuugN46dc0nIXT3HW07P
b2pZdlOtmrulvNGP49xmiQSq1nA/o52ZTK/zfMcep5btRKKVnLov9TZJjQAYu1NxcuIHYl6Vt52z
S7pdP1G6hLhPmZykgdqd7MDAraRVcR+EVHimvwBGT3UztrlWJOzCLFy0PxJFDRxC4qHJYejVmS1u
9vCDS3Yanlc8+jC3LhPOgQOo/S9386GgrgL1XAJN1fu+bHAo+AiCuyw8hEblrjYECPd9jOMYEJHT
pYbMWrCzruISyA5tNsIiNtqr//61dxMGwVzIMMn8SpXzhyzsFZQLcQdqgHMS9UJmA0quwTfFk9Pt
eJW7SNHojY113jYhvOnqkeIwVd9LPqBpjmZTQP6zAY4Zvfkj7AWraBpcRTY+63E47+QIXcA0cS8h
Hc3R7ClXPd/wFlfphWRIAVzn/tQkMWIQl3of9P0af8Vlse8aFJVHAlnCi+xIe8J0gKL38SpBRlUK
CxuM+ab5MjFDLzJuGovERyY0PU2OOEoyMfl/YXq7Hj5BlhdL38Sv2o42xsKzXDNDDCM4bElIIubZ
jQYhj8FpkTTff6xYrmZcu8enORp9lIwYApgJY/nmtX+k6+diNI4xizLauG0H0jg00csN86J8bWmW
ZBRMGSSR9TCzvmWTdPzWYVZ3x4fx7hW4uKD6sh4a9vQr0RJF7w4WLv+51Li3YcZ2j4BXAUlmllM0
1mI326yLqjskH5pCeGlpk+rVKIy/v4+QA+Rv8mpKrfeeCaror3YoP5xSDlpwPyWESgkWN+6u3gQR
trXXoFK3pAJ9yqgkCmQprrCSPkO0UG0UewktA7LzJ3Dpd0bbly02u2kQjcHy6PvoFmiNE2CMX8Pq
N1wBoGOZ8uMM3piC7bLHxBclWtOteEOQl8P5XuxyGHdXWdwf0NCYCXKpWc952RBCOJm7/GY7HnHn
K1zk99WES+lPFyOUK47FJ8Cr+hlvam5osrknlLNnmd4wOls5gP71u7VLwzE1iG0yBYkE/Z5oNRWb
B+tljAVmpoEDdv/2RHhlYSX64fCWQVmKYDsmFKdH4KvhvxYRgxONcsqm7XoJMxlEGyxmD+1kLk1D
Qq1H+y6Vf+0ebhzYyl5QLpF2IKdMFIMqZNYNxVT3wPqDeK3eY0BUHDcsYw1OZ3ncbOBPzLgcjD4F
dCp5X3eaNUdilsyiKhL1ptkLD+ALsrsUtyRDbPzfl6JpBBNXsfXdpcAc5EswNdx6uNhqfznujAt3
ngt1kwgBvQI/xX5vIesjq59+xm/vYD8/WwODEaifENG6H3axjmeDAaP15ZGUxn/tNUOB1HuV6eJ5
1dw4/iIPNfyiya7sXO9YnZoKL7qbBjgZghy8HPUmeGg3YVvrDtxcir6/8FXRq+eQUN9C2GTgpu0/
gv/VshwOSeHCy6Pf9fYWrw39S9NFc1Kr71x8oWMIeJ4WmNOpgcnDMtByM7YMJ2kQFdYo6/L7zTxs
lTOXMKn2kavNOWH8G5XbQ61MMo20IgPBqnjM6QReM74BaAD27D15Q8/8BbOqAkcsHrNq03QYpsBV
UURH7UxdsZngCN1YG8d6Qx6Ps50Jsv2qXo7+ntB9mrVtUM0URHVhR4/pq1IOAJ1vLz/1Bg9sHBo4
tzrsSMBCBP9nznFy+MQtx5kFnT4qD4qAbd9OeJydRM6GZePjkcG1pjBH6FcQU6UI61ClOfLrNCrN
OiZ+2owCFIWpokpTR6IACCzsS5/mU5cVezhqaQIUL1DdVKr/jbD88OOf/coBEKX+AZ5Nt+VWo9YV
fLUluvkf1uN3vCTW8RE7H73K8zzGJKRpZKZQYWbwl9GYYkXWnuL7JYQ8lADqX3Ipb8Z4F9TlWfPv
j3JotRkvEYfao9UgHbc0fypo9F4GpKO3qH1O8YvcFQa95lZnNZTcLsQrTdpApnga7HoRBJratSk6
gsV68iTBe0aUdTceVAcOxfjts1yqNE2HKG1/Own+DxGZNOY88hgLgnf5w3DYMDPvQlmNvmOJGc9V
v1iTLJwkXfwydglMls9LrV1Dy8qbTXFQjrI1x2JGilf3qQ5TqXcl7IhcLtuRGIUQs01BJNiIgUPZ
I6WCKU6LGL2ZdXGDME36IDyXV0I2ZeBfpGhJ923Nqe4MgIGI1VslPKJ9NiY+lOlHeRLq4d+4eZPe
AIBzEcznVhbGb6pZdRuELlFlDeLL++myeFTP+WmcNiG0qtPY5cSdTdt8O8U4WdYXuGkaDPS/7QrN
3LUxjqk3XZR1WGfkJ7eM3hGT9ggjm7KHjRHuFxujRVk1711NCvKCylc8LCF12J/54daWCXmqZRRr
yO/uf+UTPDKrANNYI9dDkea7qpjzkBQ/kiITqM+guY4Z52bmtfYyes7xUlReAaS+qNu03Dr1zYtl
0aZuRvGc0hxioVhW6ek9ql+U5fi9tp7td81NgeAKdLGQeRkdZWH/WeRGCfX4vCXqvaYUHMZAI6hr
1ZFLn8r42mzVkQe3EMqGzV7QkAt8KO4zb8vw00tEBKaimsOzKXogg4FCesJA2F9fAX31NNsUqERy
i1UHoyFApmIXnB3kQ7HyMhbyZluY5WjSb9RdD13joGPFLLoNhJRL8j2/XbasmIhBH/X2T5zYOnA/
ieh1L8jLY00uIFXTGISiDfWzK6dgduMLUxLtlqRfEfd/2zC98J1suMrkuKzL5RkfROWTZxHnf5Tf
cc2KUIRP6Jr+rad8v3ZJV90E8/z8sB8+MJYwoseTKpH9vN8Oh22Bm5cLm9quDkwR/FIUunLCgIPi
hJ91laJ7O/Dl456zWto5JaL5WTn+KuF2mezY9i1bulST6v7ywDGWeGJBthcjM5pckesjGBazGUTn
ckz296V+WJluUe9ELjR7Enk4EaVztEdZf/Bgi9vF8Dx8T45+2nZwCtlwGgtRPOF5xw70DY6+2GbC
YUhYZk0OC7Jor6ySC5z1lzYs8mE29Ens44N9+53061AtY7hhb9ZrgwHeFzs8Umc5XzrPRZ/eSKG9
7rtqUHuWlNXCy0TjWaHy5I8COURBq6DetTZ2jSFtkc3BFt0yNCACh/gWzX7XldjKg8PjqeovEIca
SXWDP0uzz6GIr9xlobLlJzq/foHTrzPjCiqTeTVcrh9BkMA03HiWIbdaXZClgWpG+Q11861ZdwSG
a1DkTIyLNycDHayUtauEAQRb11zZ8CqVYR2VYC5USTpi8irAhimuyZ0ZtT9GlLpv/S8Sw4qcoCw+
qouV1chtivUytL660reHyXJZBzLKk2pSfTQCsOBgrktuQiwlFjxxeO9fymAMIXlHbPdffQH7qb3a
bVnYH/7EDbImCBJ8guq5sbHmJR/S81vBv1FuogcLMW/Een3GHDP7f/EssaAakdZhH7+Q+WdaH8DF
2UowkOsuvUWd91of1yc+7F4KrgfNiuNpjTN/KYqZzxzBwcy2bAi/LCtmRBezhaVtV+6j1dq6imz0
Xyb0LxTg4OAWDZyky3MekKk2/0vER07A0UeKHhpUfFnZIFWvt6rcIaX9dq01ml+2UPBWV2bTi9ps
gvZYYvrNPtZGuezwZM5GdY5itzYu7aK0QvmoCgtzfbjX8TTDZR60RydUmYg7gHC/+ZQhk95+wTQI
2qFJiUbglfr51DnHzKnF1x7Vt1vsoi9zEzDqIjAlbY7o/1H3CgCdyp3szx1HMMOLmHEKKa+ENkOf
racvdX3timNuokOy/BHoo36bz8MrXlSyL1IWLSIQjCwpuaqblCk+vDY6ZhkE8wMa0ifjkdDN+JS6
rkw+orW8ZXvleG039Qnv51/L4Wt1PQP9oPkOGRSSFQPkzoamKWbSjqK3eRnVPUhAC2QV4cIXVmQc
r8M0TFmwC9JCOK0NckxKu756vEqFQP0Y+et30GdJh4Pt0xi67GLLKSSfJCuc68KDJXL/mo3I3WNY
kSLXK+JfxPunz47/jz+TsYCZ9U+YyGqJjx+OelajOOkiZMnETW3+XIqtDDlFEX3HruzHGLPstSDW
0mADNOCyum/BsTIpRu3b+ckSw6IiCIdxPbjeNxsX6Jd5ppvfmrbNdsFzSKF4OSILCDy7SriYBZ03
fQPiNTgHh0/YaCXqaOYQDchyurHJkQvRP/zhyKl+ER6phIDY7Zn7DW4X/5ZJWCH/kru4uArNt9wY
CeSjBTqwoyxRl/iUvOYxToDmrl7QKf4bblRCiK/AuBmRBhjmGSO32uiHbShWc6uNtVGlGni6jt9y
I6getNH0gAf80HgC217ClosxuL6PAlgEjA303zpVW0r5xDukMoPSr0yyIFgm83Dt3rKimY7PuG6+
sgloMUChUglCcLUPLTifwwIMbBXbQ8uWo5U/XxPY8aPcjIT9AIXhACJfj+TkAAwLv+TKrDcHBPsT
+f8Hkf0qpiDEODKnKtQHSANLJBEg60fjdz9jfxFMhfH+oBLWT1gnYh5VvhBU9atA6db24ww0U2wr
Wj4+UTG9zb3ZcOhPHYlQ91B/zFwZ05EUCWOFBelgz4+GR+HkUl4XUqXySbCZdZ57nFMWmGCkT2I5
PuPELvJxX5Wz1V27P4EW4VI5sGil4l1FAfy54hrHwDB1BAljIr+1eL+sU6JcgmPtvU1B702wuoop
Mqe7yiTmYpJfy0vSlQbMtFc0ULpp6mGuWO7Zn3wwoC5BhP/PQbT9y3iriWuGrNyEgSErxCmgbeEz
YnH8aqGRHpDfqU7o6EeMJje4TtJeTJn5IIDOtUAKPwSfIngHj8c8CW4GKxXZ+LyVYXnr5pOSnGXa
LH9T0UUEnvFwIvkI1x1QmQC5cbsfAMdwLagp05GHRJUbtvzJQXLWSHfREGz3IFOpqS+JpR+uMIuH
faxPm021d1z83FVKLN2PAQAhQcSdZKGBEJmi+NhLf2bEEPrVvV6ywD0Mh5+1u6RlEPctKZm9ZQUy
KCW0q6xxxhSZYhr6rcpAqLnCwtfTplsyDnbya7iboqG00V5TzA2C9OIaIzfk5qPMbTpJDdwhRpZ8
9BOrgzT9gG+Gcq02nZpEOkClsmCHl2iMFt9iHJ8C1zodsod4Tb+13LLhzzTKfUAeAEXtwDo+9UIL
mt4Tp53KrUzkCMmKzYUwYGknBGI61j22toQhioVNRI/fLjfqXpmxa8qelYPRzBQetzon9HTtH2wc
/gFUtpMSFVbSAh7EwCSLEjRxUdKHK3eedKS7N5pGx9r0oSjN00dDE9ygiVYzapXOh8NccOaNgRnX
P8ZWbgnxf00IiswwYE+4HgwqYX/PvTMcAwNyvx8GgntLlRPgtUwBuo0DFI7AicqVNDwbJwx9NLmq
p9j1bNa1BppEjcBPkxudIPyjI4nkzp8MC9KgnL3YZtaGtgdvdWBp4YVn2AycTOfYxZIwkLndUN1G
ZW34AGQOa+q6hSUX82uVMr8Gdt2oRuX/CXD/AQQK4cubBj3o/14/RAQJkzmXzdyfGgIqPLeT3cDI
ZoBKG12VL2YKTXcma3JGnJD+jEcttC5NaHpFWtldrAFnJZNxozTQ39sJD2tB4mYUYOC78wM/YZkm
o8jbf2bG+ekmt8zDGR0gQcRIvy/eSl3EbtCK4U8tWZT6PAYCA1vofPynT+Zp1jBAsdvGracM+keO
4UUOglu7J7m7aQAXBq7ImQuCqNvtFUryleSfoMwiRacYJG4bCgYc0MyxET2qTqg28VsTaF36S0Zh
dmnQZ7x/8VHykI7fP00uW/L5J4d4S2j8cRvpKFdeCgf9mfH2tmnluGZRS4By+7ainKGTN7X7zYvw
4I+hbGqmdrG2D6e3qZe61e7D+yj+mXolx3aUaiAmz+v2e4403w3QJBWYvRPPIcmRr3Tyq3kzRcjN
uY1ai9hq3cMOyw2svKG2LHOd5nmSzjjk5ZP6ZT9MYPb8WUVfs7kn9rCSTiPwTuVESoJFTn8v4HJv
TU7UeWO5XCqjqFRpft+CIUfzFHVGOvadlG4jgQKfdgvj5tz6USfGLqvg2ySgBOa6O0z5Ce4jfgB/
nDK2kUtHWYnPovdQiW/SZlz+X+zNjL1DQiaxJ+JmbJKo8Q2kcjKYaxYrzo19DaqFED0ABmgSpRA2
KAFHt5KE3go0EZ0nJWnOX9ahmPA/iqDRlYnr1UeSAPDO0yC+ZqkEoUsspUNk2x4o1qmRaiCy0g3m
z3vpt6gkfIXZTAKAItaYDpqa5t2Sh/gQfXmlZuJ7teZMQzlQfqz/3WnG2sU8URRtPl5Qm0JjTL7t
2RZGrF5tu2a37ysVlBslwjOaYJsLESQ1yvPveDRuC4gXKj0nlgNLCsD4xIQ2rJfG7AtGLnBs8GI2
BCChXXZpOjqWsq/ycGxPuevb9RfQi/orwrcLsNGYN4Q1sNhak3VBGP//om2wLi4OBfq2t6Mnd/jB
K1aYgl8bRlGr7R/Iuals71fTnGFRyTN9QeCXl61NYWqlJ+pqMSIlFtOMWbCY4I1QxPwJkkfHHOOl
omhsg8oG/QiwwNI60+47rsl04nNFcq4h3cDX4fctmuDjEn1G7YtbMvLv4NY63ldQV374+rYGBQWS
dmtzMfJ4HbiadbEl33ZkoJ7gBn4CqIczFu0CrQhC1N6k5NBcGkzzDd7i6gGNQuftFEAreCAfML45
BoPf5/ZTWdn7+iK9mZRc38QWOTOfU/Oz4ZKK9F8HrUajGQOX+RVJgdcB/8lFlZcHv0w1tdW8dKxl
wFOw2Q1Kaay6mqHxtV4V+aSe/GTHPsbrf+oXY+YLD63k1/uBJjth4l+/75AQnCVsxMMTb3BLjEws
hqz9pcKHvmHche0gVQErGrHa4Ut04vMaRmgzdDHjUg1D/VnWOvNmYnQe7kkIERPDITkC5mefWuXW
pfMZPNhvj2JAmZ3RJ8nCv97Dp/jNyOVI/oODk0gy0jpSfpg4b+R4Wj0pgH+TaURW0oBRLqqGlhFB
rUK12b1X0AWkXrh3n2m76A+mHnslgK+v7XbByxGhW/Pvv/ZOg5om/0zlDlUwweuLm5QkkgQzW8Ix
D/BtBTN0pqc6aFvIuDq740ja1JeJNxqfx1qgGBR9qyXXXL/SP82G4oPVTYIQ/HWFXoO8fkz/NkRY
xkMRgJfvSCO6cm6u45w+haBpTC6PkN174kZ2D40h2UKOh29zJYZaw2iZ2+bjkARVX81jIF4YLI0E
w7tyDSMca4MI3RIxensNwBNL1GLpoejWYQ1Gkjb3lWi7fwoWIRhQsQckjKPZ0MOxP6L162NIZPUN
SJrQ0fO+drr3+mnwwW1KyUtjFNMTwCDaaW21ovZ+4Wb28S1Nx0Pldr62RWG1Z3xmVCmJHr3ebUno
aFyox1lMqpH1jpeeTgzw7eyD4MbzO31jj+T2OXtMxN06hFh21rUEBQdcsAoa0b366Ie+5+/V7nXJ
xaos0Aml1z7wuWVEgBrkGf9dln9QEjjT4d9mRFR+gqXzuI2dQKgRtRU/xy9e4QU2P2DbbvXtnh2p
YvT2A2VfOLzlQi8GBVwh9VMJlVmBJTskey1UV+KTmnIdfwx1063nZh79bG401cNwuoaE0ikzqLSo
p5VNh96B955Hvg9aE1Qw7rXs1Cs5s0XgxZ9p2Maoy9KXveGbtR+WmklRSbefvFkWa4XSq6eX8fv9
S9nJkvg+ZUk5/gftmO/b0zUYHjgFn6veawVy/HbzUJCY7FsptO9DTZ53B+WWUVrGDQxlFzOEdN47
AQGpTPj2nfSN++MmmMQvu9qSbW54YzPHy2lUWhhFhB1OWZstD3D+Xv7+ExZv7DqcZBLX4lFIKo0K
U+QBVl2ww9qxWWpGjWB1KsfGcDJ4HJ2s8BBA4aHXA2zBuGjyAPCHULpI2vfOfgMQtq9dQQniTD8K
6FgkakGl3pECmTyhI1Ezu6S3DHJGvjyTjZQBgxlV4czuTF5LR6qeQT39l+AxZ6y6rI4L+9V/UYTC
LwKBwl93mRuZ2NafyE6OShklh2XT+lLRlrkJGcQ2hcC31Rd6oxbgJkRQ008KsSwRc8MJ/OJ0Ss9G
5Q4nPZfYM9bgyvEWQn1kqc7PZPAcmbkVk7qGPr7lRUh/uH1HxsFhQNzh01mkrFnnKxtNzAEbVBVw
QzbQmiWS5SIKE3+epz7dl/NoFesVODrkR7AyEcG9Xfu3wOqGFT6Ed+V9wNk1Nmwi2spX/BWpqEgN
3h5QGLcKiMzvLSU7fUaSApmAc4cZRAUZbjIBuntWTuQT3fWODq25EDYRiRHksnQsbPhaXFX4tQFY
Ti4doctX+gFS0l0HCBcgykQ+vTD6urT6gfYoeWirpKWrjEA8AZkhuBP4u5gyjHjM8C2LRRd0KJT/
sJDCska2uKX+xoG9IvaDT3HNOm5Bt0d7T5b052SdLfGJiOp8H16WXrdd2xxiiioL5jo29+rduHUy
pczj0TrGBi+IUzjiyHn5pgk6MAeuWAqC5aZ58oG9h/obAtv6q9ctcqD0kk6THJiewqiIwaQsDVhh
B5hBDWYSBpei4Ya+5AGcPlC6nAFwjAWnvDKEq3J4e4SAvwOQvfTEYpSfnQ2ieB1tGA3w2fl+FPAG
z7KWPta90TeM8Pm/cvjceAQe4wPbKzRCNQ7gbkIU+NjlDzpVUisGoC/dyysaisw7c/Rd1IiHZGMo
PmfdmH3aFmlyP/Qq229Rx+d/6jGOhEe9puewQrzyCisJS+Dw2ZxMu8L72WT1ZhtANVuuIS6BZwNd
H3D1KfIHrYiNShzQH3OW190JFqxV7hflBIaGUYvRfp6skBS73GVKXvTsDvGr2ucpYC0pTYBheCrG
M5+3cX4RNrgWgxafpFhETTczOtiRoTfV20hRzr3W0WN+wVODlxFuddS6GqtI0a5SmY0Gov/llKt3
sVXaC7ZrC769sTCxhLXVfh9jhbbRVedvL5DNLdeBE2fwpjlISLrQEPppqfAsrESV704o7fl1sKIg
540RLjmiWVFwpG+qs+kRzkaEr4+JHf9JncIp0gQliZ4OpT2OQAS0Mrcwgb7a/PWACUEpDG0Orp+9
y0jfefckicAsJbDeFM869rG9RIb6YgQWe4n6TzDmHWPQT0Ya79rZp9cdRGPzSpSkx2F++DDsjnvR
bDUX8wdfEenn71WyXeQGru71R99ytSwFmz8bO4m/2SeyTzZMq20Wb2V2jRAAgaZyLgdbNTLROp6K
5iM8DIwY6Hm4/UbhUNBrtchXt+Z7d0KkeV1NRebuSYC3zc35GZMb7Or7pVBMKgH02y5P2Bz9MYLG
W1xEMb1Z7XE1J25Dsojc3oFRIdIKghr/cySw1LFeqEVfdPshWlEzyei1FetB0lM3f9+v+8t4Ixgf
YbwEEZ5F/JBFOmOb6Cs3DD29Yxd9tslJ2qF86ywCkmTPuxwgX8ix2af5TCfVnkAYrmEi+dnyDShk
DmL99CQS8VDQlPQdqFgFenmwY5FqGwLrUify1fMXv0EXWoGQMo7xBpBIDWmd5bTYWaAIcnjIC6Mv
zjL+GhnwPiPimYW8wjN/0mbSq7lGwyvEDQ6y5otGzMFpxqipNOmAlwTK6udYf7GJUynQpmJirAKo
upEhDT7T8vP1LM7ZztqcjE8JYYxmzZO0yLACZh/6bwGTt2XHlDHbuXJqODwmVeNLAzDlGYCEydpd
A/CinUnn/+mXNf9PhtVfYKN8kYLda/+++ycbs+xVVXN4kcqxFpXvFaRUFVomPgfXaHTkItlcy2Zd
Ahr2Uj1CsaLbrdRVo7Y25HHQYiHBzbvrka19sf5I05TcAw4deSF9crserGm0Jf77NneImAYwdWfI
y/OEo16QDCL0BfiUn/MkrO+ynwdUWgDyTPdCwOUtzktywjqzBwIKmkj/obXQOnBtEJ1190tHmKtE
QagO3/6c6+9M9hARiACdhHc5SbihKj9R92SHdNMpIUuF4aLIOUHW8gXGNy8XmSXZfDr1WxAG5aJK
HvpFWPgqrVJaxl7vNkmJDollk9bULLKkkJnLtqPeUE6EfLOrs05NC0r9iJQ+q7udWVqBKD+F2SCu
DypeaQVpn6Uvhka85s4U7Sj30YJJVGjT9+7o3HDzJUcXGmqK6pZb3YBXLzOLzkDj82R9/PA5UIq2
rYfPauqi0H9eKKROVlbwEYGws56Lczs4v3k+WPBoUP6tXGSxnh9rwSFwcwNSLXpmGuo53Gfs0g7s
X0ZV/twRytRBDotUXX40mG+99XGwWVSDx6/NnwKJBaaxInMi/jKdCx+gg+xoq50gGUu/WP5Wy8/L
0z54itNayXo3e+nGuoxOAvSnnEU4bdgOYVPOyTTdy8G/SOWwFyQ/U6r5gWl+yjZ3HgdEM8KoDLlq
vr3vxYgUdr4fH8oquyALlbKtd+0D6KGbQaKZaRTnMDPu8dqK66hkzGyLMZPhv8RGv2mLaRevv8wn
mhvWxFj+ii8XQ48Un7WnpEBigJrEkNZgbTmSxWL12if8MzLhZtt/PMkktVcCyv0DTpBE8h9JJsrC
DCyBZ8ZsofysXJHn5yIvT5AlfNie5u3OCwOjD6EVTw26ndZwGjLdJLwgRn0yBFjhF4gtP9ZHv7mO
kD4x5Bs1Vzd/Lk6ApbuNl5pH8ETha1366ykbNCzFUsyZ1ecXyFbH5uXAjKuUW7zQcJjuouPZ3rWs
+nYuSuteJilDheqlHaTkv+cJRAHMXiWIwhYrYSOTKZoqNNwA8qX2IHVCjAp4kWj2uhC5qkowV1RH
GVjMUln/ZsSsXlgxbC6bAyvMFlYwMavcP+uf+7RzQ4Ks0ii6kdhT3VrWlnF874Yd8uUrxHv8VY8l
ZdhEIbSbS3mTN1HJSf2ZPICMavNnIKU+QrxahVeJNC6hgEEYMg9wjxZLa/Cl8YQlRXzP/Wmk6d8P
WuF+V4XIw2JUiN2cNJUv2hldDezCx1LOURcAYi3k8TL4iTCVs6Gn9dzvuw+siryW/Pmplw090f0k
5R0lYgNIrfW7QHv+VzzaC7niHKJkz+Cp6GkhDbIt0wiLG/FLEKV9/Pz6qQuF3ck3RLZdFFI5TUwQ
jYbjgyA0zQGlVa+jtRYHj5pAPjL6Oq9Ih5e6l6CBj0UJbZ6gDxJh/AkS6aeNZ6QsRWyWsjtUilWl
XR6iar4AQYMKrSvjEjTLhEy2blR3vZ/MauXWWNhMEjQCw6zZA7Amrt0Xv1UtXsYK4yc6iJkKIsMh
lMZwpfzNGHiJAE3/Tvxd1txEy26rbrgh1Ue6yr3kkCDAzH1sgtjJe0EA2zTJE9AUHJxFKbYjhAz7
I5jScfUMjtrQh+nT0nF0APt0Z0ycFQU5ir4lgIpQLe2F4iU2YgqZmAhvdYKitgIOtGw6oIAMUxX8
feEP6Tzlbg58nyhM0HZpBLVM0HzpyQ+scPNAtyTG7Wno9QeYZKUwG6xE3qzn345MUgl4liy5dnQ5
zIc5ShuPTsMxbY5uH0hfd0jeLsBXIq64cWelAjUPlMWgn0niq+ku4k4p7rDZxO7ZGxSmKr7hKQV4
a1ZDFoB8JeSirh7xc9EjikmVAWN0yWfMBquLTurQoy7KoCJAKKHRX/B4u5UCZPkvL2MFbkkPh5rV
DkodOgynezpOlVEABtH3hJzA3MyfCbSm1iW1K/H1ueInGLQJgE4xFdNmMAbksSn4DkRF/WTdVHS3
4hTt2zeK6uRwRWhnAzw7ZANgaaISB28BpO73Zp20rYdH6hwXJU7moxl55o8nTxrwlYLUr9pXse5d
wVYiVx7+T3Y3d0IAuH8sx/HWK7bU9H4yUesOV3kZ9CLv+ei8Hqs552dgnhm4Nc6KciTAfWRlf7n1
5mher9VGi60cLUUSAUC0Qt3CEaKeGLcSn0wzdOrKGcTiSIx7E9wYUtvauQ0MA03UnjCA1PUqSOLx
BeEOK1mkc0kA4lFkveEvnxf29oa9IrRJb8p13DEMOE8BXXNeOqu6cr8GDWZ2PJuJLsXFmEusMgIf
MTqg0D6v4dEvsQOSnqIDTb4DNOJ7F2khhdNDVdmb1dMe90p/Q0Um0NfwcUE3fY8YH5J3hHfUr3f1
c8RA1mY+ERlAb3BT7HoKJJddkLuOw/8SU7K7Fbyu7MshRk5P0abaAyqhJ+NITxvh3nIfHay7+Oz9
as8bh14EVOda5wHi8qNy40asPmvVc1eDvZtJi6H4I0FHhZofkS4gzZoXXiZpQkTjjEv+K7+hbiqh
raH3NVXfYHalZoB/t+Z+a7OFdCmoNu8zukEXnKI0SqvS8fdFrkOtmH89FYTje3BfnX82uA/yUTvy
Cqf48BGc2BxyjwPspYWeSAnfpOV4cbOuLVv131IOHjotfPEA1czoULcbXtvEZrU0yfcVhwrSG3tt
5gCRVpcTxirS1ZTyXAl3vsyDfWvLIxVCfEdcs8jOYQLpObjOjCb/OPCvwJncir165W77eMUhxgCQ
S4M7202V0PIAWiMh397i1ZWkT49/J0RQfqs035pz71cVtgGLbqfJVDDps8hf+iZzgs7qFWKFG2FY
BFUWlBIu5OY76v4V9OzBM0nTZch0npTtK3sdM6F9lCZtDYLA2KqwdHq6Ing88XOeW1L8h1wC2f+Z
nKp/A1+M3x2zCdaGt72UyaJuMnwTiz3zriSDSZAWU0k2eVgnLW4x6eQ63//6iOXF8/U9/1UIubin
I9seNnjVyJpFRaaH3+yxzik6LpRFekeflPFlcurmnyaAvyufnE1VcCCO0CmW2x/VjdYRr55VHlLj
REwVcGIn0MDv/GWX3y2I3aDyrP3xVOhMGFMwawIePVLPVAvHKLehFFPR9GpVewbYPKhHJrwdYwie
cwiDCOgN2AYawvmGc5xdbWimz3QAnOla+hHn9IHwXa/SlUz9U1bY2xzJQIyQJGizJyWT4NddHYRa
VQt1k/rZFneScStTzhKgIfbuEEKPFzA+JONacrf6Q+nl6ztilqMIxI6xamtHYk5rRKf+0HsBjawa
vwaXqKen8gvKWHx7c/dW9XF+x3W+K7Y8whlOiY/oc8BBTVGunV5kd/sF7lqc52AdImfDBs+wdOUy
rFrRyOgwyYgISl04o+gFm6jRWP+rzD2syKznm6f/mB5tHEjeZak4h+59DKXmXlVul8DWZ0CgJ4Lt
xvjvrcE83GH4lAaLvkfUuE2q42++Iw06rvsEedoHOew60/IEzW4vzF/jhntqtSfkvBnZ0PXw6LCT
6AMeGzkyV6AipXLrlCVAUh0HLpxvP0NfjtnoqFAXYOe9kBjWL5vayPOjLaLYxVMoSHX3+hY4DJzT
cXQYB/g5bOHjOfswEec6hQDBBWNqHGi8Vg3TAS3joIEm+J4bpsym4gcRsje2IiUw46PFioUudlvE
sOLKDNFZJgNJtMFQ+qGcR+r+gqLBfNF8NBlFY5HERpmFIEfpGfy5f2Ss1wgt1SnP7FCZhOgvhaeD
8Px9S2X3C9eKlHReKwRNauk+v7uh1uDSszPZWdmsBdrbzbJ3qaWe2KXEqt20FeFPDs+VGodDPAMA
O8aBFKOVP6e21RBKtuF+X0NJ8/2qjLjBLELble5amKiOoetW8KvHkq4r4czEq5AVo3a7slqxSAHw
XryqXwevlglNSKPU3pkOCAV+ajSKibm3oPkUN+UstmnzcfW2Ztix0gwT8mMApk779m9qzMpoPSCj
/lZMOFf3m6jc93fdYJNuF+EliWzJTLawWD26E1BqORLgaDUXj6XXZm1hwXQxb25yNcLDFM2+1Qam
wmRN40soGm3EKdzXwnwLMAZq5xHnPGglbLEpXHPqFdENCnLHBAhUdimfJG1DRaI16a4ueryt6GcM
77wCr58Ft9OukLbtU4BW4WHN8dNNqPQ+rVu0El3ou7/d68y72lkRC+TcNUzJm/OEkT+Hz993upi+
qSCESlQqB6B5Hme8DwWe3xIIm2xivnciKgvyC/ox4G576FFWKpnELmDJ7FY22c5CXroYtPfl6zmI
KH+KU4lwc1dSS5rW2ijhZCwFjifc1Z9miX8AQRDRTgdEv/BugYZb/RHiwhao50mq3kuGwxOYGVEw
KnSFJ+wt8NAGNVSBK8/rgcl61edu5/9k9EfHAnw+nqT55wllxAQDBqRrI5MKn0zSefYJJE/X69eI
l7b1fQaYvChGqyZurmAAgQGQ7W/E9XgIz7N7LyuA4AcZJ2GUB5zJTB2vvr7nb9X+AqOrrmJ4dqZ9
fortZ1o2jM/uXzEPs4Dm8QtNk8G9ACR4QW2i6fsahJ0tHdmhOo4Kaf+1mH5NHa1KrlBwYgzprRqH
epF87EtGQAIkUVaOZEG3sXsPH6POw3gwKriVr4alouzxT4PJ9LTUU6gwSkyePc3qLW/5jRBZkIFh
aEESS40dzw8Jl6h/Anp1evCG1stcVWuloOy2c1Ac1T7D9kCqe+cHdsrF325zNJ8ZBfE3Wg9833ur
luOGEjufqO3UF+9hw1Wj+HBKpG2ilIoaU/+Qu3X01zKasfGpATXtP0cFB0iY87Xjh8zw2JdLqH2I
Cy3uQcx1CXSAV27F76bDocoCDMmt8tiZoJPy1j6BPVu9oVOVFkP85l4KucN0ExS6NdbRWl9YZqXW
rBCghMrZjEszgE3IKbDOhv4kJJHiIgFJi7xhUT2a09iAv+eUESLQ4RbzLQlILvX0YQ2zySahCRkF
5YHYFsCZ2WEzSnAUFZZX+EHUAsRr7GQ3HbbVSlt/YdI+M0V+YVR+MjiHyugP719ul3uNG5VFJwAX
sUywFXoeRfRGvb7bvxZ47RPNaHy8yFldo3IoJLOUTRlRebbVyVgsT5FDEfS3kh0GsYdhQKREzLz+
U2ES02KbiL9JnCOO27MYPp6XKqFM+AA3egVcKuATSWS8pZiDq9ZjoU0sgHiygwmVCbYkH7Eff7Ma
rP44G/AblUmoEnlIlOwAqwxQCdbIVC4Q/U+uqcZrWtwSg/DQWNAGU+pUnd+Cap8AFYAPYiGZLrt6
OVOJBcU6vdwWelIGxvmPR85HE+UNJrOA/kGNY7KcFKp4Unx2lKFxiMtAxCeZNHwavaqX58w9Xwsw
fD2/pxKtgF/eqDnv55FjhB0cgW/49WEL9XLFmy3gLXdczz+VhrrTvUniHxsFIpQTLYuxH6xmrF/R
iR8NI6Q3SYjEPbL0CDu6mf7Wzlyvda5Dgk93kCQrQavg8zL8wIZ8BYfN1/k2PgCoKxiOFy2Nf0lN
BW3l/1HbW1yEx5+NL518ToSYXiyZ33/kUXqYdujcWq+hltPxl2JYQLe+bzpM2tIqH5dwUJlOAJXe
nmCtMToJT9KfF8lbI5srWfVl+jWVtdKAAAQvO6I0YLre5OjSpwD0d5E1YdLVAUBjotZkw0uI70Ou
1iQoEJHyVPTm+jycG4mc0OU3DV1Z2SSdpa2fG0dHwjaBSm6un0ltWbtUBBViM8/WDdpMmE+D39Fa
1kUMWjykVYVWgrZrXI81APFVU2AWsLO8l6StjXleXDCfhfVJG4Ja+stJ46mwNkPWbsA6YJC7vB+O
kkDl4GXWWylWObi8rYYIj4OT3CGp9Ev9R3h1ReJXSxXOq05rocEvyDzginTFHSNFgMeTUOXwUu2N
4FAxwk7DnyoWUAclcOb0f/jesG3XJIZdjrP4o9MzA2g4o/d7Hf70+ClsvmOmFHeHzgvH/4wnlk6g
TiXZHuGxWvDYCw5HMAB1W9adu3A6jD7OB8kZ3ZB90bwLlpKk7pnLdD1+03Utk6OU9Fn92gonYywj
aVxgu3Xt8rwzQFKfKD5TXL3Ye+Nj39efYFdrFl/qEdgZx6kPxVrHO72sx2ZpNS3uRQKFP/h/evNu
SCWgQsPV8BdIk8rzI8wRTZv14gMehnoevl4arYkJ5JGGy4rf7R+9EEXPHG9xIolKrJexAGy5CEpq
MUsVjzgBO4NUBIS/j46oTAA72RlmwA/Hx5QNWY5U4wxnCL3xbwC9PtM3qAU4YdEjoUDucyMVfWiq
zC3nL+ecJBebWFhCTkkcRtrKcDB6rYizvV+QMmoXra4w24zmuHixJz3AdcnVQaBeBCi4voVJVZpd
0BiYgoejAZwCjfEz4KT2qVDptIrRUZrRZ8AggcEVUK21wI5i/X7g7cIGPGl+9HQCV+0jRjp68GcL
G0kEU6V3+QDwkw9co+plr+WrU98qdPYNld5xRheD6rxhllweg57bNmgxBFQWfqB5TphWRtntyeP8
5kl4z5PBkPFk+61vBbkspnPpQoLoBEnaa/ECeS8bJkELybrxFbbWjFnpu95phavN4E8rg+Uk06mw
QMJxtIlcuCzuzn+0MWVI7JFHneW5sPxX9TaBG/V9gIDccs1w4p9/onwTl+YaXS+yJVI4GqmzI1/G
kmITQCtBOR7K2nmK14wDjPeineCY2fakOMKC19D6xCt8/Bn9Oub3CPsjaBsR/jhZt+/esJXuU1TD
9TTYse286QiOxLMxYeYAm/02fqPeVzQHT2C1JDZDSnA5VH8tPCXqNxpRFa4cqjxNeuu86ZENxDzL
RrM37DWB0mQHKICtKddpNK8wxCnKluOAACoXscAxl/WQxlAfnEcMz9cq70YzGxEO+hsUhpO7zXLt
DelrA8diC1GDECnnn5z3eMxwZSVT12qz4cDZ7DaiuO9o4Ve0SgXgnFlhvim77zDTapq4uAQ7aOvU
OaLIcDj7M13bUbrTob7V2gUpQH3RySPbYLLMtVRdlHzts7pBp3wXU2RzPyHqUqQJ9PihFpTbLVBk
3tW6EiYdBaV5r9liQSsjyXzCQKtWpNJbM8Sa5Q1A2QgBOWOTOFkTGgupvjEZET2vnWqN9z0DlHn9
zC0qdxJgOb+l41EnlKqqFYJkR0vhUAED1JcgXPLbVrF3WIcs2PZbmBS6n6hKg+lrCCI96V49Qzlf
taO9IY/91I9WL4Z2HwaKP0BF6fFsEPVtoxgb9SGivE/i2ICPbqr8je7d5iM6wQN8JVu62UBwjvkJ
OKM1Nwrl5mHxizLfCEe0Y+jPOzbJlsgI6Oc8wb3fgBxIUwycQQ4vfsCcPIJ97cFK6Qiy/CEW+Tit
bkZV3VnzzDi2ADna7xsdIX8JU+gRVz/IEt/8ZscrJjZeXWeA4RmqC66EzltsdgIFFuppUc9R5tT7
P21nZFTcOVx3KmK1W35BGXHm+KouWop90VihWnC4L09jkQ0vwqHNkWEP/HaL/ZYv7UrjSAt7t3ZM
/MMqWvl/KNhXk+yoUrYH/K+L8GgICoDkPJOZ9Bvexupw5xlXTUqlj4dqn7aDkl6jjkibRl3viNBh
IvSI7C6DSdH9tvF+m3izFM+qinJfgx/mtNvByEVb6Cr3jdT9P+2skEFSlEPQZw86gy3Jcu72bXVd
kkxMOVTC28KrfCBFRuCX7epThRA/Wzrx5HwTSwXUMn74ynzF/1ZJXbAvtQaszCrkbqMW94Fty5Ga
EVxBQ4+aCYNVOLG79PPYVO/cT7A1fMo5hZ4HkTAKtVXidcRW0W97SbYWlUphRh67ebqZ18RlPUFS
0j00wl6NEB4pdWXFUJeNiCG7B6SJOmdAgrrG2xa4GWopP9xWmFw2MuR8i4XtPdkwrnzSPxu7moUf
pp0+z62cJ3fhR4wjmJL6v1qiIqjimi8mw4s3cT9B5siOurDZ9sxVEGh9YnTxUBc8X83XGYyp65/q
9bVpNnuE+Ppum5/rca1Na2UoCnZYZV9L0VDUdpTTTGSg14fpSXli6kDTEHE2lgfW3AgWN/8ySokG
V4p1MzdFGack5PgZWQpuAvHhMW+o9SUq3RNDHWREcUloV3txHqTLwzjQCfhsvMXOUdjqvtgTW8w4
uk4bMP9Jxs2MF/97x0hEIt32hS0mt93DGhJW+2PEKoKudx2utHbxpT80wvqpdcMvumwTNfgVw5u+
esklZNSUb+0ELJNT4JuOcTco0VJOu7WZjxzO2r1nBX+TTDK//FTHDHwJDPpGp5Syc6Fftzl6JKXl
u7tcfpW3/mxJI3E94RiyGEDjFPOeGmdbQYL6LJynFgxncRTJq0buYqG0APK26tfK5i45KQikSApU
T7uBx0eHnUm2A0Mj6sd0PlJxftqjhbn+WiB3KOArATMsY+kcerf0vKARiv2shQhyGXxvZSSHmc12
micBve32sIB/03+w6wuifhJ+70xIwERzf64Uvm8QlBoXi+u8/MwSjJk8QFOBdDneAutweSgTAJFL
GUb/L+hyCiWTdXkSFU73A6si7cLqE3rVnyKYN1uTl5zGeZ12Ndxkx+LfXdVGBljnj0a7RkCmRlsI
tpkyiVsdF48hhZy10nWOXs81BpWX9uA5m9DJL+9mAclXgJVwEy66gtMxbYo2H/j9Z4iV+nTEI57x
8uVEtCPmXQxGj/juKOkRQHOYKOsN5ZmHkI86AxMIMIyGA1wFOweWqD9ceNFjKb7Sj7dLKWyamsrt
7eXGyQYhLgIRi8HISEzp9BvDhEKYesxGviObB4Ws/bvSpdBB66jXC754azyvOnvVp7SWdrUX7FnX
x5Htu458fWikfIqISW1d+r0eKc6ezlheKw8BNeol3TRuMP8ngyVWbL1/OmFW7cc17prF9XA3fPou
CqrrP1y7Bc45sy6tjSv/BkPdN/kbmb1qrSlVJp8ahd1Bh5nPiPG1snGX7THxDH2F0IRuh1ztZ4tR
SIY2eO+eMFlIKs+BpjGiaNU/opJ1mFQ4FrNAUiBmX8JeClWv2j7lzfKKhGWb8KJpiFJFgpvcLe33
WeHtcloGpZNkMiKuPQEb+Ab7A2tWjTEPgQxmM3VLBemjlNtHQwJuOGwWTqjk9DiDTDDkYyTKocfI
RJVgDJIHGboe0pYAAEo2KpwW9YlywRmN1HsbBGPChT5NPkH8dIKZVfMLZ1Icr+SDOGyxc6zX/BL0
MYEopUUyH130w92A7FFZLxhkuaU5kHAVw0ZKYAkE5dqhHCTFhFJQ6h9a1LsRSk1ZhM/9hXys4ORC
mdTLJGp0JkDtMTj87Qamv4udE5rfyc/i0sCrRdBi8pjZsx7kqDb6Drg6vrhuywKU8UgXC75uU54h
E7e0xy1bQ8qECE5MsihuR7RobUcEok2G8luvJveyEKVrhQDdYgsqSDtA77DS0+1j3MeQQfv0qwso
FhPG3ALDNt3mrhNHNxtQR7yZMtypRTmV97IiW4CrElUTyrKEJ/j8Gbmetevpm7OzWFeIfRs8FGvL
u7h25QbebkI+KztWPnTca+3a5jRH2oOZXoSAuzoDLye7Up+K0kRACWDzi2xq5FvDeOrI93m7CA2x
PqsyftZaC5YRs2dfIYxeGUnNtyW76ggKuNoyrdGWd/qCvVDDX/mK6ff3qXH7ivgjXinSmFiaopdx
HfufZTetRxqkHSnTxjEZPaDIPLJVOqMdXkzjBLgJont8daX6OsnJV5tM4roNgxvfhgV+3qm2rJCT
BF79BOvUcJa8dE9byXeQKsbEMFr1aRgoKTqed+EQkp1Sh2hg/ORJeJs7yWh1cfYtsz65edFQjfu7
GWBlGyaGyG3gdFy6nFV3VAo1NetoDrpmhUFJJP181i2M0xR7xLDaetyAqhCfYhYzScYMm6wrdvig
87yhei+i143vwLq89RFX32NehgvNeKl6uJ/b/vnB6hsd2z7JqXtr/1yAnMTIm3tMAH/IbGnQ6Vx3
Pxx0PW2c7DtuBXHIB6GFL5wRbPNZ90MGcc2DVxrAayiVgH8uaVAmYW7cw3WSNKmWZG+RlVTMCX63
5wlMAkBXU5gr1Tt88y64w76ocNm4DT6GUwCGxP+DnDCFHXNscWvbdHIe5JS/rweVUj+U2DQbfzTR
yVb1TRfqUVNwnvyQAXiDn1TIUclXEgV6PE5yycYOyvBi1cqAh1cRg0j0Tg/k7+lQJCvlZ/zoj7Ve
PMq2SQ0ynFt9PMeznxAVM1MUi4VrCJgph0+rXTzu4X5uF5s1WTSxG4QBpIem7XX3d0Bgr/F0lIHF
TwQYLv2IDQtoy0jJ1RhaiQmude/P9VSINUwiDWqm//gi6Soa27F9djhlCi22GQIBKgymhXNHQdwM
hDqQdgA8ktFqvOsdP6xzmkZWINtK0CaRtMbxKmQXhqE6qXwOSjN8Wgko7ev9GQjJqU0N3MSfloNc
YryXD+ce+DncBLMFUv+iGRJCgsE54eg6yt3C9CSNUNTZh6TIV0yxAwVA3e45kHADtfBoI432rYdR
sNTR5RMwneuUNSL6Qyx0ch14J/izeB9cSOQymCRFjiiytXrQRF/pD8LpwW4lVG5E4tl75zZBl0En
WP3eIxlOx69UC4ApCKvnHRX7d/1udNTl8CPRAdDrcgyM2MuCb2Am02EMRrV7rb0BfM5k4KpKnfrA
oLtGIEdGR4cG3P0KTHoK7JRvOmpGLAI/bLZ+fx+whjKMFQamBsBavUZ8pT4g7UNbk9Kd9YPrDD22
GlkhPGL2o/lnzXr0GrDlmo9crv8xjtthOmFuVC7ZGQ9fd40R9dgsB9NEYS0sRACC7rgoQm+6wSWx
dC1wjoPTNtt3gzBtY2IN4emzuc7Ck+7SHY88ACtW6wWnnC1Yvrbz/pLkkBKcix43/Sdfq83yg962
b0xxH2SK6enUrOMQqrh6XcDV2u2QIjzk2tl1HzIKxTzdldpM2DZrltjZNhletcpk7d3YEWflMvge
/cYm32M3MfRzRDUJHsplhpVERRxmrE9jBjiJmjdWfLZ2PsHyQ+dZ13dfBr34AjrYhL29eos3vrsX
Dhj2xnzAJc9XC+6hPwVGmv1NgBj2W8ufmeT56pxU8M87vILK+gv/O5KCoFBNqdp/I4Y7DbinTiFx
zDrxV6ElMcNE7m785o34zU2Ev2ouAEBzxuf/h5B4HaOQDGlATRTkqx5g220kFFS0NA9tuL8IE/D/
xzKQ+yaEGRMAIMLKcI7RIyoDk3Kck4Vg5xlhq0d99y/KTHIvCHJUk4ENDF4ZJ4HtDaGQUi5mB3wa
bz48CBgTBLRXBFuJWJ+rn4Hcz00qiw647HBgF4DGOHyJyMj+h8aerOFvH+sEjohf05gIq5zSsaVw
vprRxwEK/Wzx2JiNu7eHpXHuC5CP3Cv3NVoqBDSLJeNeknNfMfc/xIb53LoM5oS9dJgeXOz9sKg3
pJqaZRs0iJrTyq9XLpO7UqeEkbWFGV5EcSN+lDGWEoPYG4NkvgC6CDFdmyeERxbllFCAMXXFOJ5h
bDB02+b1588c+32bwe6ErOLHsmm74RBUrcl9GjE8+l1NH8gLKk/N+dm4K0SdktuJT6R9aThkOsiL
LR2YLNlBthsA8PlfOn0fWN9Zo2PEfl5BCvujonvCv5tTV5P5r+sICuLo9woLhUtq/FI2sSiLmdJ0
HRstMC7ZmNhuFGivoEApGEcU2nEwwi6yeKedYpRhbCeCLTFEZ/LzGoasJuyERXY3aEPz8vDmWuM2
UJeV0HMjRNdK0iliBTxqXZvxzmgVYgwNoHqFGIPVWrPUo9qAcNIaAIupFnGieTLo+xds1x63xAa1
1s4hvqFTlNsXSkvuy3Gw/4zCMicYOhcGcx9JAt1wgDIHUuMySrEcxHx2Ts6X4kcvbiKOAyiggBmW
Ce0zOBGrqaIb0yn49CKU8zNXs4IHw9G9MUEKgJcn3dI7wn6mEgv+TppxlvRcrhcM4t+1YanO4HpC
lEsIKdogN3s6j869l2WwPTgz1seuYbktSKsyOgHtxk7wTSzPsAz22SRBxATb3zNWRjWKgbVrYXoj
woo5xDfjPq/DMfkMDZuKLacF/Ke32Rh48YUWXEfxpnSPOmW/ym6mUgusrHFz7LXpJ8Pa5bgdO/sR
LTtld6TolKZmGj+t/bM9We1FHMddp8jNttkc9rbMWlmbG++rN1zCmwne6tXdd1TThSC6B/fVM3jv
Ge1cHc3zGgoVleVLTKS/pbxsa2U6NOlkbEG1FYpj0btb1+Gng03o1nb9JICs2p+Nr8my2x2ihMjk
rQwn0XwEImA+mcvp2c7eboM5akEoybMzrRpT0/TuKRg4EGWo9V5Br84dy/Pp+yfPxm6z77TphKTh
BhWHkUwB4NpXFnwdKE6ThYgON3mqI+vOeHRfE48t5cKgJyNN6WnFar6ECHPiqZfNl0CvlFw1nfey
7qnIgGPp0S15eCxBrWuyaEJCXs12lf0jaIfjUGRKHMN/5iV3SBRa456K6zKOuHI8fycobylgsu8Q
vj1ZE4JcouWh051rnxqBUOY3D+AjIcPINX6bXzp6/mkx0jUMZt0aeBkqgQotSdBzULoNSH6K9jbp
A63ZNeK0B9EA1w8jHty5tiXS20Z0eQ/D7QhDIBN+V2e3Ld14lxbVtVU7Q5bSdjIuobLzX9noL/1g
t9QIvJDCEI2PI1erq2xkJUEmdrzeSOzLg3wmWDoQ5L6ltlxVn2mUYnb7AfZgE8/O1Ibjhf6dKedT
16y1iZ8UMJQH5FA1nw8SpvRneZu6+8PpvZlXD7pne6ZIrrqa1HTJPXzlNk8Mu8i14BNogydAcJQ9
QylvQEnCWot+HhjFjBA3oDtgNbNENqP/sJet6uE7Azxpzkb/AyRVii/EJxAtVfbQw2GjFaGYMktd
0gqWvbFMyVLgA9d7tbVbiHBuDUL4cFBkUtml272lMxKtxGXSpaX8jOJCY+y5/+3dnENroyJKvda2
PpWvOk1meiw8vAuQ4ZIPxJ3PI5A2C0G65swCqFMqVWgwxgf+adI5HXNq919fDMGYhoagGnTP1ERq
98yJTSADcpyiEcRBx4UExd7IuRG3NMS4ZqaxJTcW7Z3L+OdEl5NSaiyTwohhZmSBEpBaSfEAcybU
TUUGSMVpgPVc6+HEMWF+p1jFsg2JuDM+RFWThNrz4kY3bMuG0SCKi0Xx+evbnhNUjpZt+enBwJwu
Y+mqG2xwwB+y/cA03Nf+lIuZH4F3J6+haV/Iko9Ps2V7HG9QFZ58XcXN4yF0X9UPkC3gOxHztn2j
1IybK4+u5WAymS0PED1vcmPKH0C21b7ebrZ7lqxWvvjnH/Hh1BaDQ3kF9OxmP3kqW7CFebmcl5tF
sQs1XlqFvsBqBZ+x+1SaaVvsGntRrJ3yKYFNzRZNyJOPZJhAvRWmtr7muRPupwr+McfNWmFmRAjU
9ktoHMMIRQL84eqsqZUnCEavkIIhqMSjmqfVf3E7Ivxlypb3r/wPyRy/wfF+2FeEBJ1heRnYqfxY
z8gHgW6Xks9JG1MBoHDRj1e0FkAuzjb3dfiP0Gwrjh674VsY+QaS/8SR/4NR4/mWY3/IcQKsPol4
4W3uV2w2sYJRj5qeIywRROr/uAlnRO9VElrwmgpO+LlfskYWZSmfSB3KY6pfWE73kQVvciALNMY3
glygqpLztqORo/q6WBdBKm45RocaKEjMSwLCy6qTjoTkSMVSd6fxAxwrYkGovAJZGYEsF44G1Tib
sAQ5A5qPkOiRYj/OqlbfHE6GxYAeL6Xhonkif5YhPPHx9KcC0PCwyMbTrrBlUWcg4FsJbbZ/Qkw9
lNJ8oQukVIvbzDQu7XjugDJHF02KANUkvFLeKY6AmoCB3y8Bu+RiHouI+FC/MfktU5f+ZFLdUWPp
t8doE39DHAz/J6yginhLdFld8u6i4dS9CQSsWxxnGBy8Z1wXtYRmv4XVT5XcaMmhZpZnAVz/ZSbX
YPhFy/jIxyK/Z4bwDeS3AfqZgFnf7awbnZmvCCruicNcJqij3gH+aDo6/9ceJ8oU+oTrGFrBrGSE
/YZyCzXK8I9E2qA6bPobQFBHMUR0oXoQ21tmwlg8Yz7TW8Kbo02IDykyN96VxCQJTCzVy84JcEtx
FTk3AyRVZD7BDvw59nMZ3CyeYKq7+u3Yj1jsFeLt8ZQ3t516kGUypf1WZvxLLTO6bTPGJGrHHPcI
d9ffO76yENY2fSNZO2qxJJKmRrMeP7MQ+Mttca6dNdKUALRh3w+HxsiL8HY0bwH4PhVW4jJq16uQ
+yCZ3u3uqqPcN4Z+lSEuHalNLnhQUZ83IiAb6iMNvk3FESdQvzGpmD4sS+ZevXUibTV5Ggd+xaeE
EcAGZ9lUEkXHC/UgBjtRREDVy4qEasg9XpRO1DP/lK6ARo1h1kMlso9Oex1SGe9K34JuiFr0a4z8
vzIy6zetsXcIFYQIp9NxMQHLpQJY+Z1QvV/8Xg62H+4cSy65oJOU1RK5ULaM3vsVVRyilnq7E7pH
/sxfNxzrajXMhdDFsvtlEdNn6KtzUd7wmlSliJCkOMrzjh8A3vua0LWwH5AWH+LHztuuT04EgmQ/
rdL0MUSwFUWRVthIhkjMnPlLHhYRQ8svBnbzGdo3qYmmWeCHEGxmHlYgIZgDC/z3MzL5k95kgSf7
yOf5ea+g+UJuX+MYLzSmaYQ7vIExR1nPxu5vQAtQqVmyh5nfxr0Sja5S1KnbWMqjhDI393gEeGtB
dbEWk7Fvjyf+V/8+YfwC6VZgPaf/LsTRADuTxqaEbfgM7hrDHzFJ7FkH86muHz6k4zdh5bn4J56K
XMoKfhAUYhazyOWYKNffnXk1PaDPlSj94mdepQ4aQIrF4du6WdyytTvk//1WJxZqW7L2nRHp7J5W
XFA12BEI7Nv9Q27vLKrXOggEaA7KhEBwxA6ymjAHhJjOP9XfclNPz9TPCCKgPdnlWYYCL9e07Ou4
BSt4ub+Dm1yeS0lrf1jUTKoIlrhupl8QqQRUptYd7ov7KleqItWKbMpp3GuybLs3MZF+7WoQTeXw
g56qwAimdE6mhUk+6g92D7oGsIQTShWN/GBCmAgF7CSuHlHILS5EIs6LVkPtJc+AKDt1A/oQJG/y
8bGbaqO4ahLtHIu9hdFXS269Q9CKFGz3dV6Yiq4kFhBhDh9BB4r3hFcUOQzPE5nMROrHarFWQr8x
x/VQODVH8UyRJpOmo+Ix3mUmmpkWvL5bbJt6bDU2hntRqpitW/3geBAheAhnO3jv4ll1HVmhp+FM
zwCl6Tw66rLnhgMHbEKAhICU84C9/ruQ11P7KRXi/soVVIvCKIDVR/BPmwSyp63iGEbjVbXVNmR3
rDl1JWfU//juRE767QnjQ6meKu8gTddUoa8GLwmY+8S62UfT2W2/clDPZlia6yU7+XQabarNNBew
HW5kF0EiABhw+/9/eM1co6H6qTWZisqpbK15OSz2jE7oyEe9TktZpo5onNYEJvSTa25le432t7+8
Gqux4S0dRir6o4A/MSBfRJ/LzhJNCNzqirOQmXj7uMSc8DgX6kqDrLdukTiqKsD1I/QOgwX1s/9e
tuNW/GKNENrGVotk6X/j0HfIs8tjb7/vSKhIQDQRaK6iMGCYcF3Wd7Ihi5Wl2074igFwaVBwyaOT
n9vtrSr6oA4cxHB3LSkNQq650XkZPHjOImEUAv5TMW2lWV04CLJ8PXKcY1RTAzZTvI+lii87NdT6
hwXRkD2NqstY//pg1jn+d+hPPz6VB/Lx2cBQ+wokJrhLd4kMHX0apM52VA/I6ypTIrf59K/YeL1k
bAsW+uxi2wVnRW44S78sKBQUMOK2+1eSywxE8+1qh6HjfW4woYNwvt3hqMTxyqLbRqNMBg1IKTer
Y65D9Lpn5T3sQJgSYzbzAfAVNMbe+sUVDhQtaemKMi4E3xusMIoapWp4Tx/tsQVonSPFHwpnPpUj
VbE1dCESmcCLkShNvKlAxs+Z2t0S/K0DYeTmM9hbum3k+AafXviEETDmGpmgXCzqcFcJoa32ab3o
SM63jJ0dH1FHeMwkyq2xCsS6gmDTIrfeKb+leQFlE2caGv7FRgdg22cZixF/tglB8qo7hxvqMjFU
rLpLBaaLa8hFII+y2DmNFch1tfdkyma6VBC7+5JwaD9mJLyoGVOw0Oegxxe1W5qYBHFWAC6cinYk
JanUDA1N81Lu4k8n+jQVn+KCmDaTvWOXi/QGdzgJAhRIhxvlDGv3+sjS/5D2t60vMag5dK/asAM9
tUl2GY7Pq5DU6ZAp0a1yQ0GjXipjjiPR0fdrwn9mLNQ3DqdTpoHif4PBiE6pPcB4UG60GesXUWUD
JIsXCbf20da0tFHrgqAX86Dujhzsb1pPB+Rz0RYOWTsLXGCK5Syk+V5JEC6qofRnY4pAImf3SMnV
ZG5Ocwt1/wuZV+k1Ek8bmbjn9tVtxonh4yBsSLdq3URLb05RyhsQifJzpFYwEBAJBANWPywruITZ
U4WkZYpTUjT3zNb1PVVjW3CKZLRdY4w8KjuW5w9NlyRxkzWQ4yxNqVLYha5x2TKac8WC0wTo5v8L
/rEDYbpxZv4zUw5Noicv66EiYAjWvaTUQa+JV9S/TYJ8IRO3ml+alYKqcs+y0/KyWpQz/2YxUSIy
RDa6usLID4PJv5PrbEaNC9K3s00SK7tYOpkn39chU+oCmDg8MFqmY5yLXLm3D+OURS3MnX9nfJ5T
sNWvBShuJXdNBYZENCm0g+XtxRjtopGvdJDOGKQLFNmiRjtzIdlDmlOYYFursCMc5ZHxju6TgK51
ylpVA11mW1Ohvt6GRPs6y1N5SZS4v8mOW08+wHjL8qgMRpu7Y2sRTE0l1el+n2ZrWcG3l3M/EocD
k+yA0pS+KEHCCorPa01vTsaoSEDeWGCotTT/d/GxKO3GxlhnGEh2Qcl+kpx79iAQbgLVwbBRu/3k
EOjuVNT6PkWdG0kXsK2+fcCaAWtgpZGg4tJvS5T/bWy9B/c76kSlxfpxLWBObBuCQgq2UbTEs/o1
WyOB6jTAkCSAZjHZWwgzt2YiM4qo1+6kXrLYFTalmHuNZBy5bfhH8uNsrr30/LOyyIHEqCDS3Q1h
GHSFoYyT22MyMbA/yDHaotD9uaKidbJlkZVOZhOfuHsBUurebDLdTnzb7hJo9sxXiJ2yzHbk92yS
ZUK4xs+lY63Y8qlILKxdaGQfDRE4Zf4Ofue9Rz527q7wLG2evSU66xWN/scmePBmMoDT2iwWjhWi
YuAQZuYWwA9YkFnkJlg0NN3LdI+lxLYuJrDr47TYJbTlNw1Y2MHZSPqCUkRWkI7s3WlH/MvPZl1A
laX0zAM4wZcwQSvFhwDj3A9qLkHnm+jToYcTdjNj7Wd0Tt+3SBr88FyulKCgkzj/UB5idzoNCgi2
jTOv7YnZfCyuO56bHnL3GJaz0y8WVQDAETri8EtQBzyakjpE0Zolll8j9wcOhPnQU+UTatPeJT9M
QwO1EqOAInZyDLmTMQ9BKib65j66ZmkR9X0sOh3zBe7lvIEiFKBPweRXwe2t8X8ggKLHlRfQ5swW
RODrE74dLovij4mR0/hVF3Iyg37Fi6AUo0kZKRCoYQtAjyBd5rHhl0FzfbOauIOP1J9mhaxY8dTH
0dyA61/N3qoJHO2i0t0T7OWsPs4qOwA+cXnqe2Fyq/QCUpAcAo4GLvFal3S/s1MfIGupx+mDY8+C
Qp/ZjJXet899aCQj51h+S/8Oram7LOTPtsbipr/1Cuv+extfrXCbBJ/dY21qf5pj6w+jbkj8ePVM
sRRWNbDWkS+o0XAtuAUwdoNd0eAVueOnOLxaVu7VAcmHNBqORcYp/pd6Ftm9yqSa4Fnh6VpwJ4Jo
6LibY/2ftUYOrTRA5tK1F+A4plYO5k3nXXnwV4R5TtkEe4zVq6lbq8eQppoRi1CX+rth3SoEA5g2
XDX8X7MM8JVP/80R/fM4S261D+WzrRYk6j9AzVlJqHMNDSoWVyfIquDBO9jQPdQILASdMyO+xqLB
3WaiFQE9GPpvCSCCHEnl5oJs6/b4AXGctAPEZ7Q/0UyoVFm3W4oEMV+PVxX/qX62eoCLI0RWz+8H
I1MT535IZ72g9x30c62jdaz4bVdErfOtbdYC4wMdu251j8UezJWa85/ldaWA+EAXdys/0D+g2/SV
Bkdg2UN9dkMZ+YsX+Eb46F4r/YeBnHxUJojcmmXEIHV3cZiOydW4kFIR/c8f6eUXtu2X+Me6y7Ty
vrMOKw8VFapXl/PbAqMZKUy2HULaoYE0p2f0FlBtgxHLFH/lZa/TcinCnxwQF1z7O5Oby5zMZNto
zlvfMowUpaXhO4iqklPU+bEj8IB9r1IPvrNqgF9BiBCSJMvjKZUgY7VusXhmwXCOu6YFjxtiIb2y
7vUTzFqMpQqsx8WmFYv0SBsGZTAPbxQNq8Y5cgdA9GRIiWVDsN8h0eUtZ9NcYl+Y5WOLTpg/WlRF
+8E5Yb/irVTv+iuoSU9d0p+Fth6AMLnSOs1qBG7UEVqFrDXIwczCGuaSx8JiWV5tWS8E3bpTBiMG
JFURuvyZaxSBF8CKAMC4NR6zXMkRigWcuzHLVv7jTtKW5xm1fdvWxhS7OUC5nPY66ayLooTjpWk3
b0SGytPcF6W90EnbOb3yITJtzpy70/7bT8vPxF2xdxixOxLTl8Yb4eERAR8wNxWWYIFZAK5jHHBY
ZFAUnI+k0rEXDdcrJ53Z8wwpm9Tqk0yXxev83bFAXQEzeoFAA2DyzQJHHVaHxu0dRLtGHl1+Rn6e
GpOMArc0QhnuqZub6VAkeQPCA2ovucY4FbMiNxhzgXROOH1E456BvdOnKbz+iiKqmb1LqAlcMidS
SOS8FTvMhuac2vmI7chnmhSkopM27NA5rmCTRMl6KXZH7TX1+HmOpvYma60SykNTdkd11S9fkgdu
M8qi0HifPP8fsTb0G11FMJKROyZ6RX/xbVzL99fI37AH9oP5RoiQA7Q8YpYJpIknwdOMUTxOYRnE
FNiI6/GMT7H3VnmvTf0WoAj+dL+PGKAKX04Ouf7iRMvclX/QwkeIoFtSU53kgC/tTUSpBMOws5MV
gJKmbSy5tkBBcvXo8+rR3ICS/54xcyUKG3G6+9tIMQZgkUMMYkVnEnQ9yVIwhD1Gy1a7123oW2uO
RZ5fLYTtuNFuHoZZ9fM5iwtVUUYmmvdjV5OLe62hAO+ooPElJEKnPaQCYHulmU28HtbIE8yQKWmM
qzq7SWHciFi1rjtTcUpJzNzKMN3IKsskpLKUsclhUGApZ8WdmXMJSmSPnMgLVlRko1jNi6uAEmoe
wtMaEr0dswPyKDVVCh/BBdnbnGqLYvXjiELviFcA1g/K2Zveh9z95CCPRFN2Y9pFDJIdEpR5CMT+
H0nmMFd4+7WXpvJOOzezcL6J/TF4MQHWNercIljWWxMdNqCznbcXIZOd4+sDh+J0dhKsjstVsusu
njlLGNEiv8wiPIgiTWxDrwkTeJpRwk3h7+tDwOhzK2hzzqGp9qyBXhT2bF0Kf0p8mqVuQVh/U3jI
nbCQlkIIzRcGmP6GHVasSrgqYpgeh+gCI2y3uiDwrxAl74JomfOr++MAfLnv/Q9OwO3txm4633o6
OuNA85KLc6VQomF/IG7BZ1+QqQpv6Hzq19ITQZRqDBvY0gBFBYEtCCHDKIPX2Xlsk0q+fd/VGc3J
0TbVwmASlZkSrbo2wRcp6/f2lTaYSiHt6Tg+lYKYEpbXLWSWHx2tA584jhGEhlamWBc2fRcSrOiR
pvuVM1HNneMh4vM2wF71NOeviCAt2xbeVjHBoWy26NmFvpEFGEym0GDYIeU9JgqVzh7J1qN+dBtX
7PR5U/HY28ygTxakXVbI3F4OGHZybsNSTDbDlXipEvsj4vMZ/s5uWUuUdh+Haqb0rCWz+lsRgGmH
1wLynON1X8jFxEdyZNj9uHBA/ivH6SrQ/IPNDyLsNym1QVPzaAdZG62rVMoeBXVMDUcwKHXy4fzq
yflJuzEr8RT/GZ2Wyg9dNxWGGXn9GZPLWN3TuK7tQX9t+WpTJsxgtI2Z9TQdkFlD4XAsyim2GrPh
uU9L07Cu44vAhsM6UM8DhyvNNdx9UkU2zumReKuKP19FSb4xif03H7bVGVTcWogUcb03n+SszxGf
nKNBwTvN6GOXi0VOOfvoo3PJ0tX+DRpzme+2UaidCDW8/JzJCpMiqNnqnFh0nL/5KDywPlT2V27A
3sYDsrO8bTSCwINR8s1auCGGa+tA6t4S6/RezhZChS6q1498dvh0MB70bPvs7p6KxtJFVgDpIJQe
VMvXXSDsO/Ig1Rkkz1XmReUF4pcvHHBKdPbXc2GWFiCX7DnZU88BBVcN4H1q+Kx8S4gJu4lu9tNi
RPCdpjY1rPU0t4aXyQeInsJ+jvvCrQEyCri8BtVI7bp7eTKZ2fHONsHkRFPw/tGVqynRiSJH6oz/
ciW6K6rFBtSmmoFaWSYgi4n4QIDWKu1VVOczxiyz2K09HsJpnBUivQzRTPU/JfPRR6rhsTjKPdVZ
foZXxDoI30eDg0CKt/BJGIpSYh0BjEV3Vy2W4S2Lm0SpjEXihRiiTBQG1u3rB/8Mvv0zPNF3E2zZ
UCtRT+cRNZNg8eL36Kk9+A7OG48Gfj7VkArA4V/VMZqVxalmLfcrPHzdnBe/7MfbmwGd8lNcX2Xo
ZPB63iVQLTuOdJQDbouQ7yAGUsYf4cDvp25EKL2OoEgVXTmd4P4oQBkyOE7jJKXQWxZpYG9f9sF7
o+qClxeCEMR8+i5vOQORzKFP+w83MFrRnPibcN7WtCBdq1zk11Ly5XxpHKhEUVaRg7V3/TOqecc2
ejNXunN4oG4kwcD33JXC/C+NfDP54WUITCjz4eySFh0yxrv0VGAOdjZEfi5B3AOccw2SSwoNYj9r
Bj7xsGAbBUXv9cBlGhel2XVzBJhI0eUppfjl6eXuPOKYnyh2VpHgfXJIUZnNdW2DZb0aQiaNj8Ei
PDxsia3H3IjllBiZ9ZtwBa+bU7ZOSy0r9sq4ZK+7X/Q+OUbhohkZkA912Jbd86aQEpdHaPLHzOaQ
8uxXzrGn8OnuggUCmyJUPfw4oCTfVAgLlpGadL5fwfXSLtOBT1TaQIkLa8i5IkLLIp5+ACa4KyhD
J+d2dVTwjx5j0W8/nihRmQz4KRWsdJIsl4dZajdBtWJStrdrzjhTCaeqd1hj6K1HoYrr/q4Uh1zF
hwid5YR6QrjKzzPkME5ZUCv7Ykd1N8+mbb5OeLdtFkuDQRK28BK9zmwYpjBo57S3n6aEWDIYE9t7
83P6yb3oDsaAZpgumvVghKMcE2mCxKrvBUyJjcKG/bfiedbndKUrwigZjY1vWGoAGw77MdUiB9so
VJjw+tjQzicS8KDucSj7XnVO7BLDmBdWaIzYEumscb/VdeJfcUzfhWaQLnr9TqPNjDLFzZKEe1YH
2MCR3ueiCmdQuoyYVEqjZI+JyXzGh9BG8fKsC7Y4LBF+AXW9QayR/SM5j8c5VPRjrfv2gMF+EUC1
P9l8WhEJ/hzLVhVHpzDCyOEkNhBR3IXqMuKK8CDl5hNwOxohfi6i/YWE6uNfrVuVvJDZv6kqDxGk
YBgl2rG1/BvQQuEU8f73GbL9QQW0TA7opML73+7TXJk6lH/5eL881LrDAe0ZujupU0tX6Bf78Vgu
oMHpHMjax6Lk6m5fTq9mQDmIpjoZk5x3e1hUozZLsQx3IjFzXCq9VIqtoUscpwwfpOiqODOq4cEM
mJkOQNlYJPTlEk0UceJFnd7wqRz0tr5Rgt3pvO/bGEmpzQi/0K9Q+D8g+R2yhQ0OTHQiGfjRt+zv
Ley2axBYhCa5nufDS4bJuSeJIFap0YoMBn6RgylDW4ahD+tmoeqXMv8Mvvhchhp9EUpJ/4sBJIPo
HNVo9qT9s0h3FYH/+5ARuCKJrM6HQt30xLEPLnaDtXcyFxFAfL87RtGgQtl2DzzSUSVYQ5AIuiVs
erP44qlcwKQ9/IzlzXvMw4kgNlxTrLKdcgUpxOwzY0aqZUxoY7FJR7WS/+JR2pzYg9STGVdCWbBV
vL6uLcTeQPI6y7lRGAH/ixcTIDucHDDr84COa86Q3PtFhAhPi/3yRuZdWDCI4E9f0uFtlOsmnkXF
NVzKC3peP/WRoTBbsHQEP+rJ5TnTtoWCj3S/Rvf1ZKwdmbqhuhbSV7CxosYEDelU9wDd3Sdm1LNZ
11r+7HJg3uY+HOvdTZkscYRBX86byjmx8OrLowmrE0GS25BN2k3rDaiwSqdiDn1HaapgTlw7j9Id
CB2S2/sgtaQ5+YFWWKa++M0Eok2WbVzjAwKA8RbGgDKjLo0vCSWpDoQHhqcchL5XOVO+tUXqIogy
Zs0Drqiqt8FlLGXp8MgANQF1OeO88uvrIuYfwDIJr4GOiyypjH+sPieUOqgp+zWeKAzOf98LiB64
5Q5cGew0q5WSA2954tvspX3CPyG+UQC19Wv8e2r1TaDpa43CNFQZmswx+bw071bW+kSZrSQ8YgoG
JSteQTq39oFPG0opZI7Lkyn6iG+kjJZsXbFVaxgJj38tawFdIwQg0ccDufZcDnb/43Dorcnc8s2v
qfc0s3+zSdy//7t76zjMji4VpAOzt4USjyzQiVfAAMsr8+KkYtYCBT1P9ayHy0ucU6r6Rm5RU6j7
4RXCjhdZEHMlPgBcjE6Xi8mJ17zkpsZ8lmOw/fkV9h9CJKSLYNcY9swsuQI8Vct6z4lZIqQtnY30
zFicL7ik7o3MTXq9OyefdTIDV0MjzPJijH+/Hcsb3wF93AvQkhjqQxPyVS4TlQCIwUKe9OQynA/a
C35wj6u94XnI5vkqa9i8sPzb/ESS0EOZ0KPyslz3HS6u0N//HshEnFYAmHy/3iSfQBKsPlfhcvJj
NT9MOUDSEVPYp91+DEIbmwB1S9EHYyZEad7vsCVmXn9mUm3t6cJpsCB4puGum+hoCOCx0ybL6fQd
SGCeTu/HCUDlTTpJq7oaVSH1FzQbmRYpF9kQlodjUO5uPDTmon5MhMhLPmxgKV3UJz32QciEq8XO
UX3LtLxW4lF3wlbOj1XlQYQ3ukFRikuTTcNBBWJsE0wkNxLFRBWmYuov+c1ugxTrHCM5xHz1oEvp
X/9b3XepNJ8CSjnWD4dyF6JpFl+UgiCk3WLbq6YuQgcGpn9PV9+Tg+8nk2g4U1JfdSlJqZl8Pzh4
/CcMxGHN6PCZf81X72KYrrf6gYkjUPYYwC6/RKi9S+1KOWYkp6m2s8ekiX0fGyWtzxiFyzO3UCNl
az3Pc+gOZMwVkVm87YyFrcRy2BIziOXYbYJ4vogyg54Aca0r3syfyQzeBKhFRzU7ByDgXC2OAZEH
ZsvdggWG3JK62gRNG9l8WpoRwKwuFRLhFLn4hmxEcRV0xCTvbFLvIf1qy2btC2Qn0DcY/ONjx7k9
H61/Rfq9fgShI3ZhBGLwFhuZnNkUAeX96Fs+8KZZZiVkoxEhadJ4sXIu//5J0bvQ4C3BHQiB87Rw
br2SgL+suR0Qi7w0ASCsB4hSvAxe+5uTECPDeqw0kv31NAslnZ/BIJLTVX3U+K8Ze5zM1QcdQdzF
1gBWC3VEMYPfblgH1o5s2dmrB5xJjJJ4ubh7v61Clc7+/OrxmOA27U4Vq5I7VX/ApzGmmgFtuLbp
egirWo+2QBNnRwOANkv52wSOTUfxurR2Q8i1e6x9WPP1cXzcbjn1itxaYpSBwyyRXzBcg/WT51Kb
EoCiGIHdFgaaqgc/l9ZJvqg8lUiJoioT4IQdF8jawQdZIEsHJdD5CChD7TpBpyT7Jhhmzcplq+xp
28PfbzIl87ncmblwtUNvXOZVV34iUO2k8Vc2dBbw4Mw5mYDyiLtiJhBp2dqoIfPj72sHB41n7izz
t3HYawcOLldMFberfEHGzSNOeS8YjsyOGUhH1yEXWdroURMIW2UlmXBtCIPUFAMoN05DbyaKOaZS
ubRx3BM5jEGcHRgu9cK4RfSPlky3h1HO4bkNZR0NSB0ZVF0Qae5MjAq0d4Mt2SJ6HSXYeb1kJCKj
V/cZbmOXzgelwtHGNQtRZqAK1DAxD1oGGj6NsFECG00ahpkrDTNrAKaQj7BOMWr/x/mCTpWnrRzF
iDgyDTqn0iPFBSDzgVBynO8X1cCjgkK7sGAkkybpyFSo+5zBnnhhtXmSPOwwX503U/Uhhr8XmOzQ
XqCAmnEhjVmwpomp7u9fk+cbUs1+W0uuLPiheP6jdQ7UJbkRjSfKtmw2nQWCQhiMLHFN8D9mOcuc
ARKlF37nv1Stte4D9hn2ui5xCg3VwXRY0dcBKX7jRsWTdQ40XM3mfTmY3a+sSjI4LQXpNDOIJdgP
mCkGf3tLzV75/UJRy3Fb2ABWXgohJpz1/N4H3a5M1f71q3CrlDNPRV1OzW5ltTRoWqJ0nx2oSGvq
ugfjMhrqj7nx3FOExcJsAb0HEc5jWUHAcSSlLhrkkaBkTOizl9yrJTmKepr+/GWbtrz3j4JtQNzx
tfGZcpizzuwK0DwX+fL5oyPEYbSdwLrxmuf4iVOKs6mvxBwYgFWTjFv9APZYMS5r621teqG6iddq
XaG8u+r9V9TpJmJObZGww2VgAIPAOzSBWBhZxHJnxI+cKopYDY0/G7o6h/eKLUxYgJW+x3kzLR9q
YXgQ+Goa+P77WokZfcdprBx+C6kOJobYCKETJhB4AgSappYMUGWZwLznnuHgkK+rO4Pr6CxCo6sw
P1Z9yYNOl0cuZ8f7xN15gG8fnU9DK1KYC6YWkXZpNGDIi7jFXA+ZuBgPoafGhxSTW9s2/mBPqI9P
2h4Fx6XQTGg9XBsKB0n7tlH5PCa/XQyQ1KObwFblbmYm1dfF7F6VHIdZMKwSeYzUHMIHhWZvKTQM
6uVuUlosgzLRLpZl6nm+iK44drSR2ANp5Tx1W0XK/FWi6fDzd1LDmjlZvoFfI8b9AMlx6Z3hvyEv
MGg2rY2oukg1CvtV78qfEyqcemg/Xn9oFMbTUBZuOJksglRhJ0YysI59pZrdUBC9Rt/7fOUDYg3e
Yi5+7CQrJzTMt05lKAW1sdIAUY7Xx8NzWRib0OmNuwzVdgOEg1bOhnCfRmKofERkaHYtilnLIGGr
163uh/QCjWe55DWK1b0R08tYWnujc9jGLSLEsqkY31FEywaljASV5PBJLKgX5TjkVHOrjaxo4zVu
6NJ8D7JhNWdZUAgKajXKnUkG42aWCkmhnIgPKPUbgD6rcifST5YWkHncQZdbdFwUvnB5KIYcWI9t
U272E6dyLK+ajSDyFtpZiu90wFn1mHY0sWTxokhXmLzI6PQlNdlro6pfezoW8OBQwNmolEC3lOmA
GWJNrpEik3RHaBGFub8NquMyr6/VlctCFkw8tu0ijc+hZ/Hm7ufCXwRbl1i0efB6GINFXetSXzp2
dq7JCo6L+vXqqDhyzGZ9bHhEjhdv6ZGJFegjX4DsL8bASd+Atp1+WEwmqlDNo4OF3ipUqPSn5LTb
s8wiEJX47LFEMQtZ1jVg4gUA30hqOy0Xrh/ls9H8C5wiEXB53wyd+/Wt0mdRk7dXgaPFhiBCgyOH
TVPPpeePbPvzqmmkF4ponEPoB428rTZfJ0nJLHiHQxmApfNs8Z2kF8fdCk9Hwj4cVYhqIs6lGok7
516Cn1jWEHLv0ZHmFF8N+0XE8AZODk/x0hF3+nYvDCdAwnYnYKddlrNww1pAQT/I1EBLgRE9JuUk
bpJqqwAP4UFi1gPWQ63N9V3E07LBI6D+tWy+XqK9r65SSfObbUhcqMXYIYSQY96ruDiPk+0MteQ5
lT6EARM2/jYawvtxJOiTigLOyqEQ8tq6M1KIjDdzAykF5nqWilLWQoS4boIxy1m6dhnCz5HmAuYX
v38vEzdsKzj48bKf/ql9dQxOx2Im8A8HaOOwxnvdxYWASrieNP1Ni8RL035+/r7ygddHj2XWlijs
64Uh2ph3nfinGCapY5D/Zemtvo4DbX45+iJRP19i1+QPOu8OMX0k27sLphwFeRH0w+1QL8uLJhq4
zB84UX+TRxpjM686LtbqOshM/oZtdzgNTdVGYbH44z5bjKrs0FBnnfNsOXRicJLv8XWSKpuSMHfg
/txGdlJ/mHk2Ep8c/e9mEpWDfQIZVpROqAwuc6jrYIoSGLL9QIc5amt7jW+7xmgxltHx2KiFmhNw
W1gZlgp8MHb9dZIRYVHpjle85C1mEO0I6L2Yzj/wkKUdQytJPYQzdEo9/q+hM9YBm0bqhIEC+V+B
4jQzqbjuUuonW2dplECZFcbMc1VXLNz1YS+rZhe31j5/R/dY1pdFHilUGtkl3PYlu9UbZAH59MO5
LamELMqvxHSvWgwv/apCaG+iphD0binLmtTqyNcARy2zL6uXTywQBkDnRswE8vpwFX27mZhAzYnX
RwqgBEPlpyDmWf2TjwYquffb6JTRWo/SG19+bQ2/UChYIdcXPBP9Key6lOJZ8SLriXoISiLrbdFx
Cw2ZYztLffEk5LmY71LgzvJbxoQw2QzzF9pWH1n/bRFec/D6njKGz9LE7pZ0xN5D27q3zSvvkX4t
LGkY5dPgFwOdMAgQ3ENCr/YQPGjrvp4UNkUeMsRXGOQtk+SiJXCrQwk7e3xFIwNOTVucvSuf3OqP
uJ3XhJC4VvhtciHic1190LLnEfkygJJZlhWpGtUQElxNeH/Rz8TPXyBA3WEFIGGsPT8RPZjm+Gjq
3Nn8B1gsbg6HHBwI2kR0Ba2rZTwrlK4dQZiIFzL0d8Hby3jYHEuQOJjz5SzhLbo2yfzxfvPF6D2l
Hlk+ugcV1PNpaX2cV+wc2LtgcgArNdttyEL7dn+CYVXgIvcUn/qDL1cb/DiuL5612ce6FyHoKZfB
cvSM2cRxzL+3AvbFvwZa9U0HzDxsljFvhceM+pwi1Bojd/6SOKW5Qc0QcoCvb9UGR3vk8vO8suvy
DS6/4j1ypt/hqwCSnMHWEHxpSlTc1iK3Wa5GQqPJ2traTrSLC9Hy1Zxd0C9EYFANQgPSttS0H7Wl
SaQPS6UTmh2xTZdu6DQMKqAID65FyGzZi2zAOO6aRSDJteCio9ucQJUc+RCPhElINv4cvHoWgJ35
WnsyKYezE8KRmeOkJPg5BPaD6blT/8qQIk8C71Y3DUk/I/4Xslj7S2EoFVA2NF7BwvZL8shDkxmo
3PqxIwmS6gH6IE8q0SCJky9LsG/pVDO1pSTmRYx144ZBOZ+do/HvOFlS1vYVk4q2uHEQWOr0pcNU
CKTo9iObngpdM4Ze51jbJstNUHlwv06aImPB3ZFYOpnithALMv9Vhza7A++xNOktXpnhpsXJdqkn
XHd5VqUOV3bPlSDobKHQkE2klWzi60M6fK3vrdam7d6Sc5I5uyfmNA2V98BSA0+XyTJhUqyLbmLM
G84Hf+vM7uddTYEapJpj1K6+3rJnkZSwAFT8M/SlHX1kWay0QzRf2HmrvQ/pYU2Pug1oDfN76WSp
DjcwAJHQ0HYsLkP/M8itwiBwy8Ya2Ax36TQeEuL3cI8qL9ultPafU7pzRoG21TgtyxY3LqjOUSng
lMQwyHaNJIroYS20ctvm25JWtLGkRqLesVFIRJtZpe0by0dFI8t5YAGLp7HKn12p1f/h0i/rSAOu
vWEzDWVYP6mQm5YvfA5lkIqMo5WN6Zh+ZVAOSnOju3xowA/gWvjLIhrPeyJgl33DRsfMrfuujoux
2oUd7Jzv7WAakl+vBQWXCZgbtCUKIV3L9ow/8UI5a+6P6fS4gs3UIhIpIavf6n/ana2eSR7nppCz
eGwW/OHwfHTgzD00hdI027Tflwyhx55xLdWXTqb5XexklZnoEaylXAXjChD+pindoy8X/y+dwdAA
SkpW+RChVPReWUWwAAKHtZQxp68Zm7/tncIgpef+ojpoGrAQa+md+FDz2Ic/fhFiAw4dHwV+d69Y
qCu5lkrc6gNwb5XlOcDw3PlqwviSWz2IN7KWbIurQs5q7gGi1VogVE6+QlKKNRj9dehOB7SPDThp
wDkZ7tU8xEIu86Ood7f1bcTL897jKEqfHSC4nmKyRPsvbvckrf8PYKF0zUu3Aa6D3TfYIBRr3NU8
Ka+HtE00uMormj4bgVpNH4GU0Nb/Ap9BE1QZpIIGA4AzBisgJR1TIX4IQA1K+qulYXAgpeC/QL7x
UahYIHWi1WE5VDK7l4GYqj1DQPZZxBEe2KCZQgWZcmUzh+d23KtPgV63h0lLjdsRgGQBhHAcOPi6
4qeLl0+lilTCRH/Dgr4gaxUJr2wkl0ts73wTdI/YS1+9u7wmtLVjwqEGMEBMSqoYWfhhnrJ+uBdx
qaesyPD2EXcfpMITaCgu+rlDBBoz0yyNFw71iP2Fm2gPLiAhF3Kx8VraqR3dQfs3pCE5pW6w84q7
sPPxxXTW/tu2Ot+c0bPpMUBcLBoBLERej1vbIs2UjJi2qEIH7SZWPeIdBAsy51DNzp5vd2J/Q3wI
JnmgRoWSye1HxLaa+4nYHTDJ6JANzI8eWpoYjz5P7VsDPZtFY4wcNqWL7WaWu3g4OaoPYHGY/Ik9
xZeUJtD60nCZ59xuBxWRymQQSjSLlXcpELNDwEE/SuwXAXuTHhdtL89rjWDQMdxyRxebDWuGHNJE
DEb8S/fp7Lz35x22Zfk8r3jCBgjEQ2aP7YcUj8t/O0g9vv5OAGqrywWzhBCHAJzk4cBVRjmCtaBP
W0vr6SWhcqFfk017zIFp/0tcRx+i85NhzZzyNbOC/d2raN78iJY0yWgQy6ErYCq3+ps41g4kYm4j
YNvd1uaHAsy99VZCyR0u10JZwG5pGAUZF0r01BQlUJSGp+E5oicfXO5s2tv4ggCpEY9hgXo1K4Lg
p+AhYtL7Ix++rxnpBCJav13SWJEuz4aq/gryOVuOwPWRfPHsDP/Q3AiJU9nszR77TKC/205QZlUo
ByyeJofbKOXUFfAUwN1AaatVDkzSALOIW12HWOp5M6ZG4RygZQQcZpIRWBNCgmBunGR1UUGJuiuX
w8awGQu7viPUyQyK626Mjfmei6uMP68/bVs7TiqLtjvtk4SvvtTCfuwJPB9yk9TNmEsFl6hstT6S
DFkjXqcTG9RR0Na7zOw2faM1onC1RxF+rbd8Ed1wowHqo/MNblEGXpGrWCTcAA3w/9/sM/m4hqxe
RU1wjZG+7chSWe20ut9KABzZ23Une0djYM2FpoDAiaUarunIdSksq2tH0fowoGRFrjrkPbm3U/xR
A3djznWiHDHmfsK2SMHMX+oU4cAbtt2sA9F0mkhwEr7mXn6WbTlGP1HH1u44bb67PaylTMem4cAl
iamYGVecz2a0Uj4msp8PzoXPWjeQFna5E1YX83PI4EFiDgn26U2ajf7asvlKbZIpXmn7f96Dq7tq
FH85mQcECmocgvhI/WYFj7bMYbW6jfEhIIF/zLL3M1R5pDewM2rRBbNDIolZG+DqGVjKxmKXp31K
TpL2ChypWjTJLuUFOid+zpNKChlnqq4l6hqfhWU1H2ajKaiBV2aZwTOUsMjn1r1K3HPAd/zNuRUE
l45jgjSLkEsP+EKzKwMtfMN/3r2/47BLmsmv/FPs2uha6hYYPbDoXvMHF507yPR2QC28j1wPoWUG
q8hExkACkoqVR3cya3GrvPQjicZ4uH+JuGGAJcOJ+YgVJqk/jOlaIIkfy0S9Wbcr9HpGAiHyKyD0
U/MCZJHX4EX0Q5kuhAjkHKu+43oiV9xMCAZ22hCxvsCzQnuL7MbdCXYPsFDJ4zPIp8dbvh8oVmCf
I3hd4gOofZJ70ecdugfgXZN6ch56ggntGXnK1S0TUyV5dvqKYvc793SrwoYFighvzDfP4lW32v0z
xkdWLVD9DdAbYSfC1rXGGAbtQ/ckWVj9oorLJ74M7VV7NiYWjeFuQQdCHZN6K/PlzLR72mCpotPf
smTfFxrRqy95GLXltLhRscdD7w3+aWCPZkaS9kiDdRik0KTaFy7P4LIMYIoxs+kqnOo6mPbt/SDv
bf2FSlqIcu6lQ02cdO5wjYT9nqn8eQDIK/bm1QsVWF38wLpGRZOZAeBXCRcBaF+ZEtIm8nccAFhm
x6Ra6/7+2pgAsVrNw6+Td53z+FB+lT3RN8nDmldpPuydLuaOjfEjIyycBcE6JRsEPu0L5cmqcCdZ
js33JPcgCZDp0pykKyeBdw3hE3Kj8KX8oL5fj1oSQ9a3Kx4M6Uk+79pEiDYu+u3obn2banlFlUDW
R4QNTtDoOoJXA/+mprexGN3+J7hLSme9+etgISZkEZwOgNVXS2d/xe/YqQzkWX+tjkXgvyMj33yR
5wd0JoeP1lmDqrv8i1hVp0Qf25F6zWWURBFqLM5TqOAIqrL9O3IB9LiBNyWWfmJ0XUXBfHscga/E
ZNLeSHnOevn1XrqJahEjyZmoIj9+zGs1fCo6rHRPglW54Xp0o18+unfFOrOZ6oLIr/s3nOaIBMzA
F7M20dzrax/lUGKOPcswdSszb1VeVfXoEeY9aHw8K9+VgzooEZuQ3BlckPiGthGf1G35aFIkDAhD
jW7S3CZYkjS3toZxI+8HtJzsrcFpLLSWjyUlrLGCTPzsLVRayJVUtl/Meeaup10vCGAR3JvhPcpq
lFjMGDDjDk3l19XZy2SLQfPKkb8D6oPmrud4bADxeuvx3mmG7D0PxxH7SdNvlCdaxSKYB1uO/WLM
PfDmqovJJIe14lZvgeCWzkV3b1oU3BmG38xgpnfmrZ5agJ9DpaEeieN9OTKRMUZTGHoJvIAc1Mry
spfymLSI8lc7ajq8/Z34v1dD8etvTZ/f0gYqnTjuyToNT+IDIzF/02SD90whQmQ7S1cXYaCq8CDh
FD0UYd5/UKMaNqGhFdut/VtK0+hE4jSZEpa5vYagl/u4J/0PmzmK2ZNGsa8Sr/L1agQhdvWdC4kX
Jg7mJXVq6VCwwNb63+5hYwsJyD7tYy3oeRQ6fYhxiUopL/63aVQw096W9l8pAXyqiEUoTzNrQ7Zt
6lgbKfe2GB759oq7Jum/rt9jFdP0/3Cn5kEB7UgvLtsRErxtq7YC0hlsRsFNxYU7AfJTPN2qCoQv
qmWw6vU1QQSPijcWdSHw0ebMrw8Q7nlZJyn+VnC3xzli4kL4Pi9P1zK6y/s525T9bC9HgQebBkCn
izH9CGDnOfCP/6Do2TCzrMhJXafnrdn9QqPUttFqevXk4nB2XpbA22dPOHRgCM3rLMH/0cCS8wNu
6EQJto55Wt8WPSSb3n+r2KScAYh8OcZ7lhsHRxmEc7HHk3QrC63RWWDRYp2qjJuMtY+KJZyxcXRa
2JRxzNIynksJ4+YoT8KK1lPujLoGVOJ796pllsieHyFzIpqU0rJg4zeisrdIwM4UmqRzQzXAXEa9
Jd/gmjoEW7i6a5hMPI8WfUHu0R2tKtMa1soZkyqH0uFSOhMNyTaPpvxm6Y1ardWllztxgQISgaDC
PM32yk58Ef9N2y9Dg/O/eyQCFH3Ui1AS9VuKayJ+9DRMj8uhj97HJ35sxS4PYUOkpN8OgIbI2h0R
qgtXgccIYP3kCSwIfNkVNgsGjTDEBU/itEUny+A9+kE6JyHv6zk74MSBcuBn3UbpedTVqxzu/eDa
xpFw591ptXc7CP46EMCeGMZ7n/CSO7vo7F6LRd+9WvM177bX6rqJpFdO08jLpjltn9ckiEdcU5rp
HfSudU7iUnNF7iPm9s7rO23Ho7r07wafXz5RiSaZWsF8KJel6nRcRaeXt9PMKnoIpBxFrJJBBLPo
+F64Vp9C7sb+WskOxT+NykS10DNn+DkQy9w24Z1roKTfS/E8C1sncTdZEKObDNXLS6S/aJwQpQFG
W6zKf+Zh7kkpcPrUzkvHb2BaRE732/+WOMCdYH/Z9s+fgbT3obeGWQX4iPd/Od48VTBsfxQeUST0
m4YKpDdDfAn1n6WsY4o+I4ycIznFXZn8NIS5Jkdqcf1k9Dn3aGy4WlNkVT/qsVxGzgD/mHbGN2vT
fZKyCipGUX+T/UMmoPVhmCNxdRFeCkUVV+4mAW2jQYuheUeSBCl7Qk2Tz9qIDzHwywEEWApnhG6t
GB/HeKnMCm25t2fzenFY948+Cw+rXbw8kMKhO+/R/0mSU7XlePaPnYUJ5PRcCxNr2t88EToyhnc3
u+clSrzvgHBSlQL6H6EepoCIelxKWn6saP3bNtJhGCvdVWaCP1TGKBr3QRuw8uLxvgDl21gCG4Sa
0mGcz8xjpHSVkMfwzqyLsJyT03jdV8E0YvrCwKkL2WlLLv6IwvNbwVb4NT0mdMFMtDsNICMyBBYa
zJaLxYtzeG3c95cuuUqiiGRTn/XqPUbeWkXqQL9USSVTxi0M5OU6o4OJiuMjV2kNJfIUhV188qiD
fC5ie3RQ8nd0vQB06ImfTvt+xrQz5wcidZJtAmywlCv+S5r8URu+trjNTm8eDDE3H0BbjlB4EpnJ
9qFbIF0Qju+EK9IIoCL62ahbeld64lxlkfcpOC7WeN2tiCiGHun7dxeqzrwMxFTFJyA9zJopyW84
BnPLBvcUJZP1sbxoZMcN5WlIKsAXCBHeybN4KdYRynnFSHj40UX1hrNDGA/wjNAHKEnXdluAwjgK
01mzKSp5kxuFQ8PfUcce4Rh9H5P4ODXnx7wOUdboysBJl3uHiIDx81RgVGXWXTakY1RV1V0hdVmj
Q37uye/u8Deu19JIE6NuhaAjIbkBvsvnLGg/uaNYabV44BHjDiHIZebd2cpNb8XZBQ1JF2Bo5AQp
yXKOCm9NMZJnm5k9Vq09yY5Z/V4bp+I730dWqco/vnBLynvXHIPd91UqfzzwT/hxxqNlHb25NRyj
mVy+UzHmYKC2gI6KM4mSmCS2kAgP2647j3SjhRBjzFrRpYXtMALkjzNoNIIgIvv6LAPctKovpITe
Jxm8jS+WPlzXNGo26CeZL2RgaADnuIm5m5xGxJ9P6gfXxoAnARxhaD5mJ+4Td+EWIvuabi9hjMPA
r6X5PMpgUv2tf/+b2PDR6VyU7tHOPn2/o+XW04pVmWXcJ2cIHtpuvWbnxETxaWZ3Fsx1/b0NZvow
pWmYD+sSahKa0XG+1Z0wVdxunrD+MTxXvzL5cOIQoQLSASbpQu4a5G63ad7H0Wd7ZlRhSUasr8uO
QVVdigEtmE9pYkcird7sU8W8omPXp97o0b2f6xAprtbAWh+2ppgFoK9NtD8dWfUKPtjU99BwhIig
fYAvrpD4XvD9yR5RwZnDper1QLtVkI2DyRXe+HzJ1Ay7wovtDblMk+yRrPna7tYaJqPuREnGYtou
an4Jo9lV28ZdPLQGn8jGLTdiIV3YqpZI56Q6H0NBtj6bPtHUaJN/nqVr2iUQyVSkIVrZrIXqZn1W
bDpbxQ1Kdg0qfoQv8Og8khM3Me5TDiZ+0k9Iwid2IKaAL2OZZ28sw88+pRO4HyWb63S594vw2N+e
CJLYD+p3RwkRupkWNTXN/URqkSm1m6VdXYZ1yZHUhczR6D/69DcIHIzp3riulxD4Fps6yeJpzXFO
CIIDPgMMnl18BDKvY67KIDMiHyip/JD3Pb/Z//cPBomun3zcVGMCpeWRWz2T/mDcmSh4AHewuAWJ
7rLQDXpn6DlZSxRWQJ6nwAg+YG+rmKIe8T6ps5UIuhWsxEoXcCpzglSq2h5tXl3v10xnYJeNaIdH
5MliQ0P5FSy9Lz+IyrJloZhjNLmLRV4E+NlI4NxFUioHLpchN8Y3jVw4RC0IQVyfSAHoj9pG0owC
+xVfxuixHkj9q/gBQfk4wbHvyqKYbDr1srx92ebcQeqXIxxeVbesV70mLhIsv+c9CxsluohnrMqK
n8iFX/TqvBp+3xjbjOi1CcnuvXDP4eh+Ff4WyMNkAQgKEfFP7mEcwzdwvX/dCTFhuABA7zUdJwLD
puQA/XNgqObDCG7lKb5NruHohm/Lj1FxpMaQdVOf5CcqefS2H/6ayeAK7SnJkifU6lfIjUzOg4UN
TUbVb5ALJ72EGyO2GG54UO/YGejWa9DkggrD63pA3E2tQcuTr4EhwRbPo6WU6o1IaBSujK+Nki78
TeTyTARkIhmn8E2w5CzzogaJ3zMpHCZ/iHE9HB891Vf1SUDNAsolbJaUg1yRC2YAT7ONiSzhUW6D
pw38I3u6XnVuns59tYXGhGi0N0f2zenvMCS80ipKj9aoDTOHgc0i5mdlMTPSt7NFzLXcdUYYeis6
8MBSQJrM24q7WRzwIjqaqcebFH1taPID+SZlrItNf1DNDk3AQgdgiTB4vZe0V9jgCWFLT2TJWij6
TTRhoBPG+mrV3os4gcp9tF49bAUeJmTV0C6aERbQ+AmCHr0rZtgYd/HxjZ5OpObVwVKRJ2+KG0df
hDW9UYz0znvGTSvYluxqSoGR3MvHiN92R7wzgPvnCaG9vvOZ/rQztcePR16JdDsxoO6y2eoPv5fg
I/QRmTE1WgyThnXNorg+E4q17OwYQ0bVkPF74Lv8pCMtBWPiJStS3b6rjFCTf7BBwLX+0Il0nkge
v5O3I+xOd5sAlBncsS0AyCTJs4Pt2onUHssRPgPd8Xm1yuW3I+i/4SjC9dU9+ZUHf5DxBqsDsASm
HRcl/WLm3JcacTBL3ff8VbuBVG4TDHaKegnoAnJDM/b4rFhyDZjKgO6jINX0ZNQ3XK+KWoplLwJa
8S/cIpkTrBT95pYcvt2pKdM5J2qqQ6Di/3k0NrMvYyUsech8jnNZoh8NoHfo7oVTnr7J1Mgpl74q
BmQy9CC/nhZ/UEjgaULuhwNMgbJzs0xjhHqZb44aY0oSO3Xd6bJwXFhGW8w535y91NfhH0DaL373
aCZb8diqgoBG1mH0GNv/RM7f1buxsDwTxuwzpsW1lSvOJVH9jJnNmiCufX+LvODlz2Fl12UhfxeB
nUPG+LTX30vSs8Kau23g7khtFEToVjIw5nnQl142vHay/nloaqpFZ1kacmxvG5VQJ/R9tbS4ioo7
Fhmzne16ZYFL0toWKwHxFZH2qHq9W0vi5tk9UhU+5na/Nm2b6f38y1b8R8qS7o26raUBSeRGNBzN
LHS5+Kru4iPR1nHF3xNtvGRIma7nI/sE/lCSFkEi6KPQMO5dpK3sPasYZ+OYAVxNwT1DGhBnPA/f
9J7NLHhDnR1+fCl3p3c0mfQ01jCOCUJRu06t59XOxZGCUoZxEhqUTZ7agG0nXswckz6qrol2LsbH
PywUaInUAH2B9GSvSbM/liOoGWTPrygTkmVaeYpQQb9/qISt1DJuJo9nf+L9MIVbxzOzQQHPJpAe
MbXMieM8MVdYSQfe99dPhXFv7QzZ9EQs3GBrpjxnVKLaH1q9ghth1a0Fs2Dgt4HRvqePvdWcOxMK
N6/X8q/dH55eqKcaDemPhKdjdUZAbjFpnNnNbgL8mB2oZVZsanXGeVMZwmAYdOTEWn4wKZqU7dyE
2XrgRRzUzyr0tEo2kM0SLnCvm/JhLbcOweAL6my9IQfanjhr8j427jDLFFSzuw1IP4dta3pRoixu
USaBs9npapKg3S0LS8b7EGq2GcWbujR0cBB+Z+nPhCLW8IaKixeYuiLmuJYJFlsRXj/OYZYCIN+N
N6MRo0kKh42p1oicHia8pb4o856PgAfhkNi9PxxR7IGeCscnC/lSeI6QB40D+TRWOaPPd5QVv/Ru
YGqslibgonkS+HrkFqfRhWlVcKpiGGdl8/1eMSOR8xNMrY88FpyxyoCWqQcYAHQK0Bb/GfcwMEPK
KbIr+i42cSiiqHYg8bOb63ulOq6ujfrMmETiv0QgttarHTdbUYWeV8lqPD5P1yzvH0UlkNE7EhO6
hDaJZyco/XkTXecBCCD+oWa1WTi8gtz4pxTjoYregKIHTK9kpgVk8el877kKEfOLMSLegje1uCy9
nU/S3B1lUSgGtFMCkpaBzqLibcKREkoqZMn1i4HegMqy0Qlvj3PnjByVYAdXd9WiVdVimnb+8hvG
s90Uz2AFpBQQmJAmsm6yYFjz/ZgbNPgNIyNEyFx8IkLtrUcmVClPjjYFI9ENWMFtwb1xyraBniXo
8dzHn9brrff6qkjSd8pFdu88209GyyfI9RuthajSMV3HaJ/rnkVL7RuL/kdH/ZfTr78IUEkNuX/i
ug6iLEUwHn6e2UGARyiwEdoW+vGXJzoR+hFHeLIVwNAhhnHGDDLe0zCV+KiLdxvyrJRfPljXkVtn
Ib54dNR3HCZzZ4Ge79cZ6vda9K6gtU4s6Uue/pF5euzhD2scavBjMT4RQp0hIr5ctj9DAiFTO50+
GE9f978HkQqJzocBCwEXlb+Z6Ci8cHqNcU4Av08dNvXK836bdtuCR4fvrS2tQtLf5LzxmU8oPNoe
OOz/0EuXVpRT73ZdC0lpw8KUWqMP/xNkbJf8TtlN5R4PxrLatrTY+82oYAxAd82IieVOY3Ngi4eE
ZIQoDzPxNBTZzVDfHrrBxHxmSrJ3L9kzGVN4j7RprHcLeUagzfg9sWaNL5wRtOXL3cXV+VdZXi87
qzZaU3RN/n9LJ680ouCO19vmlXrkHxGQbdE/Z1fonvAgm9+6uGkOOtnPhimEZFXH11oVRS6N/KH9
9YWPjothoL2sipd5o5xcI09gEUkc8x5Rz5b4VBxWEO5OOtw28xmVoij19RfGHXadJ+W8/GYY8V1n
LonrrGt4SqpMKdJnMIzU0RonXfqQ5dEPQVthooLHT6iSEsMRuOQOi/kVUhAoCOA6LSXFrG4Jl8hY
5f5be18hxu2iPrrOzYbZRfdQe3KiQeBqYnbk6J6Nl4PLDRus7oB3lBAd4PBoVYIC9hvVDKPhb93m
tQt0TDXXGtjM+7VEQkbWyPFeTj/0S4JVB9V9Lxs/c/b7MVhQLMl0mej/S0YsuYUbmP6aIjnOUkhy
HP3gC3yEbnT6zzTPUXOeCHpvyxbUxkC5yuCfjMgT5ORqOevZ/6769SNwgsYGjB4PRDWvUhxruxM/
H0gsYBuqnaGpneBEmifpMjaFSsQdp4KsyNd44lbKsKxUXMejZkNUSSNezKi8eoYEWeXi4wKLKcuU
/BFJMCJpMnRkDCCf6zYEgorYVdW29ga8YWtrciesrmKjfGOQ8Tif2V83/HyRVsNoYSc0syi/AynC
QPX1CM2gj1cLZDM1no81kzyI9Aq+YIzqp3rV/ZpwEzGMYhr/6nzOFu6DpQRkM0d7HMRxkNCEaF82
f3NYGTmNg3kD8yxfkqK0QOgzX4hRfv20cYNgv3d9d0YlmgmM4hXUd2J23XLsS9eeHFZjn5vIVDzG
ZoKdrzbULP3JnAuIFvlbTeIrUIbHz6DyDfE1CxxFobynZCTXW/XSWdzl4iZoAmEpo39VJla33gE6
6gW+oWiUfjSFclJ13cw5cdaSGXkN1i6m5LkRnTngQKP70d4iOAE7jvxt+J28Eukym2jg/dIQpLdJ
Lj0pn8zY5HWp8XYsd22K37gCrbjlZSLRze8xLNtNkhqHEhrmkquh+Gq5CGH4K/CzsEtWFVd6JCho
PZOo8Zn+QhxHmpzesMKoRgucqrv1hizZ1IpXSoVLg9kyPiSX1S28fh/ZtCgoRWgoNSVp3WB2Y7fs
2wvnbc6odqTtywrhLAaKpEmrcpprxL7uKpGZuN0XEVGMIN2ELKPsoqL7yBFsaMg1BNeAGVw8mHDC
lDDgwsfOpcsuvhL9zcb3zvLwEk3U9hBlkonOO08Kha9eu4BiCoAHFUSHHBgbnJZk0z9cqcbhbzj7
i8IkWrZkcOYJjsyo999dr8Ov98uvXfnGLYeWAsjBoitNgfzwwICWBPhxsFSCbJqL5pLXrDzIBex6
PVMYjD7Amxk5c1+Iy3RRdIzrDLk1DdgOO+CfZVjjYMEhD+P2/A1fyRU2W7o/HcxcmLO3p2F1kkgG
0gMViwSxmFi90/b2TCKV2qmINyVqMMPpPOur9dreVdVTVWzYKtRRglox5QXz0TpFTmC0WVryF2Mt
8+MJOSoyAf4h/rLxkMtKlOeQJSS7gySqkp8L4tQ0dmNlOL/MAClD0Ipgalxt61lqGZvwFebPODyy
1AFsDNby0syh0T9cZvr2PYLfmxk7osZB9ZnWVsC3leO26IU8GhvHQvvTRjoaL7xI8xixWrOmSegT
VIbDjVRjELlp9a4fgREagk57zt8gsHt0lmYwlbKHsWEc4sAYwA1VvZqserJ+VwT026fhkFGSwxKG
23LlgDp1OxATagaeyK4dBJMznW11p34JzE0+7MVZHjutTOEfvkkPMaBjHzhI5732w/kcs7mDs9e4
5pNAlL3gfopjjeeYF2lGzzg0gHMw2r+Pugt543mvhzSKx/OwHPUWiOvlY0GbhmgMCl6kvVr6fux2
6rNQC6M8MR+tpEsAKD7xl9yWrkJMIex0MZAj3aj4398Xietk5/V9Rhg3HyDG70SByeni0Eaa2fAw
gN7X2IwYVmGsZkC0A0daB040LWddXZAGMShZKrwwFLqL2i3DyyATylgAzsO6w7PO1meVl81Yl+5V
p5coYqjmON9gzb5+LkMNvqK/kg5nDHsVmH2RZ+TP8kq0eMfk33glysaNiU7iDhMR8ey+9noVr25N
C4OXAVWaAGDSG4auOMbr56cyEjP/uO4iQCvVcLAEdzyzLS3Eh/vQsKu1R6pQoIpGfdGAl2/XUT47
l2svdpZmj/is0PWmDnIA75479vLdpmz6xs+VKYB4BV3UxT84XV54lvvhZWjWOTvDOL3d9JLBo6RM
jayhZTnMOjgr87c528EvixugFxZyhe8oAr6Ne4Bir3alc/vAdERvEwKsMZyEhV6tidx7vgSnJwVU
/VcKxA5eV109sOY9OkHoMb0Wbm4eF5De+vrNRZ50v/C6XIYpx8tAs0ltAEENtZg31se2WfPYt17f
PiaA+rGVkFvrbCe2mChMw2hd60Swn2BrO0OE1kOAsRln0Yc3sFDLtwMropyw83BuhayoZtTtQD8N
PgtpKmcU0tnFecfSIeFiFsZsRz+J4sqrQJnEJX0rh/q/guBZOPnA3qr64gX8Be0/EATHq7aP0lKy
TCzlXAnydTB8IivfGBzvrHTBaUlrQOk94g9y0DqzySJeqRvbPX23tW9mp7Ck3BGJPV5UPLC8XvbN
EMewMqTXJ/e8NWsFIZfhXTPlLHcFoEJyd3Cmh80AJmaIX9nzvtWQzkWqVCv/QcV10uplhVP5AFUK
FsuFC+PGklIyli4G+YU3WLhdaSc83Wy3DHe3nrngHYjsIC9gmOkIJRWDP8NhgH9l3GUYT0bGzyH+
A8GXVIBWZSqg9ASpyKbrGgow5fHG60+mCcSZCH6yZ5fibh3GttIkXJZgmCAfCfya5fp4dceMFZpp
txKLGxlRg+/c5C4Yxl4A4FkWLgnuboT6e7mzcY1bUBYGwLoHYCXOA/D2gqgO3U38mfGNQY9dE1AQ
p44sSNEDEmTpF0BiwrgH2Hnyk5P2w7iVMMSHMZ9CRbNA92V4i7VyoQ5wVdfLfHwKd48SucsWa4TX
z3TC7F4K5wsz+KxzpbOePzq3SZE0IioZ9FIvyOXZ/j9uAXuikVM2wo6tGT0e8Eo13YqaM8kA9oyI
f4aodHfYuooCiGTLNnh6sXibvwHd7bPsx1o//mjU4uLrTCqjpLE9X17twasP95oHX0mWrnVWhp/C
AgYW50FRFnD2NSzgEPNpS16q82Q38iawiywEyhuORqQPAwPkQZhNSZ/QBy8S3DuV/ikQoz6S8a33
ylXOSc2iAhxpp0ghDOEdlfZFGb0cMbLwCq//d2yAQRfRtl+QJzY6QrFIMxviTN89UN0yJ6JQ5Tyi
6vsOkwAsN3Ww8CePi856mXujHy4EKIZHd4DU9VwqT5GLpBBAK//lElKdi0zAYB7vh/Lw3Bq4ojPU
wO4FRr9f55ydOqqyMCC9EvrdHgfILRJ9MGQpOJUpqKYBqLJK10ZPwLts1NqDNOvX08tVkFdjWxq8
+wzgge0H/VBfN3ilzPo5QhiTW4lilk+/JStmn7v5qhqzFsrwxGLjue1Gz11bcRCOxHkg8h97yKRm
U26cHSkbfdNzzmlzanjNkUaNBhHEXsuXPcIZAeDG9C4ZpCL2JhPIRYWhgab+I2TyQDsd5LuPpmcq
gI9Yb1VKmtFrTPMAqHvp/kPmRFOv039WCAZummUjLZLO1+xxBULoR9a8w2gwX4+/u1TasVk2qhSM
JTGVYQ3XrO+iYjp1hFnVYtyS0BCOabjwNvl6icNDb9BKHee6NIRcIkQ3yG0sI2VLZOwNJAfL7PJm
S18sQUneeLAPPkEx/m1NORMd++dUGgs4/QXUwKVNCUAfIVoHZ9NMWkY5qyRnAMV5hRzYtvjlalxS
wCYIum2brSVDZ4S/XwGa9NAEopxhFiM7EJp7m1yEuwa4NqEwd3J7U/huMro4M5mhBfsNlBWyG+QN
8XSiBLZz737qdu5qPTNo/uJ6xbC/nNieIq5U/vpZa93LCWX3OvNQoD9Msmqog93xWhbhvRLEsATx
PnyPwIdTnhEXFguW6sHmYENf2EUHF41lB+BJWmxXwO0yphYegRlf3gMRAJ2WP6/RIF49MP3CrajP
m5Es3k7wZX/3lFn+r8vUgzvfwTPiwIWWfAl2X3MgS9rfcB82hUz9yEE/8pcleADYiBuiDG6XX/QU
MIzVeuRtjARQw6TzMTNTBFPCsE75lyD5AmPS5OFxuqNdn1y1ep6F5UjF55A7AMi5VvpHoJsf2m9n
CixVIuGG+hWXw2W8J9a9EDe2D3AUoG8Teo13P7w7Tyx2AFwIUm+xORUwkzvv91UW9jC+hkiC3NT6
AFp3ZkONI/475EEdNYydL+lqXt8fpnDEUaDJmriE+hEnm4tKuG2VrL/SIp1b8NEJqJls/FbJs9OL
mEUmNrrzFZotLMEDTxnt4S+m0f3QHaITy2ci8IO7I3huB/PB+99r/OgcVyX3ZzX2EapAAldjQL3e
07HDfdpKaAMNJVd1Rgp1+6jEbPk5oRXY7v9EQHOT0V592Qapm1MwnYDD+kQkrE5IfwEGweXoX1jY
iazLqAy6z+2aNP8q9baA3XauF8SYfAxHZeeWDc+SCamqHMJB2SoNZcVlZPuZz01im8ZpaH/KxISF
/WlahmeBtmQ/FIRs+gKSsgw22d3NaWF14sg4AguZ0MOWjOXKvu0LvuDM9bnxsLw++tAii1OHNqix
111XOu5AwGPEhLffTekNSZW/QFseJvGbVwChg2OGjUF6DFzHDPxfgcvt2hyPyRNJfrPyXANsE9ss
ROQXCc/UbBiHW9oOXsehHs4twaK8ZM/vDrOPX7t7ZJ10h41hbYIOb4ntVOdSaQU3dfzwsQ/C/lOj
z0jZhVdUzL1xuYPqeR1JTk5jWPPnu9EJzjo97MJ17oxrZkPVjDPQmUgO11XYcAQHK69DpxX5NL2l
mMU8pEkc6aK3UTR7b/duYf/bu3uJWHnoAd5CfJJ56jAfxW0MeQPBQHiN/IFNJeyJ2sB3MgjVdodH
xmVQ/heHisyq99iOZFBPljrPFZVuaUGo0kZpUKCX487N0DeJkSh2o+8X0gVkQc9b32G9fvLMbhHN
iCwFkfyk7UlBcLgRYJDghcaPTjOfsu9RV/kIVWfxDaQkXv1zcJBkcSUr4nNPfM+dLryNZ+X0XT0X
OyQcWYSf8hmfGuHTzZD8Rkm6FF8ujsNG/ykydiXE7zzJZS91iuaLQhEPtwHWJeV0WQnBHOPPBCWh
o0kVQW2h/awrwR8CT294f1nLdTRQBXQwavmYAbvJBkWAo/j7WOw/nNzjQ6204Pkdo7MsDZaIdXlU
jOnuoc3YcbWmpr3hj9i/6dxZJwzgKNhBv4URq48cUCTyq5SUJ7c5Y7YO/vUw5NrnBFcNA0KpG1UR
PP7IVuly3NpoH3c11TaNgEjcRckwTzsAR6SF3OxG99Rq+jpTfSlaCN3nVESeRwsZhiS6CfuUgUC9
7lJBmw9+nWRaYuusPD5fpL2UeLQrL2cJiV0ljVQkJLMd96NNo7/1cElKiu+OaRfe2DfYZV5qcSfe
Awa/Yl5nUxh8tTr5TcuS478kK3haO0IwRAFSYU7YqxIdcQN7T9TRrs8bD1LREOkxeqSeVFuJtpUS
azcj6EnMSYQcNTUvG9JvjGB1kFD5fE1ytobmZVO4h87aTxaqdWIPx/LyZhfrn4z2DIUuiuhHFTaD
/RXGBM5dos0q6Z/6S14nnuNPJSzeozPE9Uhr/zgmRJ2Q68jwf9xz1xE7q33GBv7iuOA8yyUydgKN
04mmGHQyAr+ESddRTE8bQvfJdXu0zaM6E/1XxUxzSwfws2NPYfXSDU0hTY811oYqVler8MIKi/h9
ZMHmTbIk0uZRnqbaWk0bZn7bqs129e1wM+lIZXRX1mw6aq5kL9yiu/F3z7so1XhFwPU8AjoMgdHr
rEvc3Yeb5xmkiN4uSgShh6QMknLoH2vK8fYhRIJsMKVQlWcZ0duAZ7Q2xrTGFnD6tQHDnlhqoE6Y
jhc9ax9Q2yd+KmZXIwa+CCvICGWUSUqwWD/yowMBRoJE7K1+REU0oP+kfh/T52p/ZGzaIh6xf1h9
Gpf5V3aF3QlQuM3jcExZ2X+lDnqcYKm9sH9Reo2RW0KnZOM8jzzHaWCNgEHqIK1s1lubHASq/C/w
rVKSm1ivTSvPeQBiQi05UtJwdjoQScb4QZ00G+raRgU8JbIuGFKOT1LJK9hOB/boDLuYDa56+/jN
6THPCC7/wNKl1Eoodp3U5agvZS+zsONRyVUyCdBUE3ZtFYfsfPyftjRTn68Ut9ZI7RUXQu5AZxtI
YYQIoyxYvWOAUdJP/4W+6v2H2cdyxFShLhZSVLrrJ/UTcuZFY848QIZqjylWaMTEtJ3PRziuFnUm
BsdFFG2FsovtZO9Ev4BRcyW07G3EiNkN+xA/WkrDAwG1nSbX1sxCZ+CsHz1vHZuca8KKAbU2vHv4
tb+5n8eiRhzLRjdS+MjocrQU4ssECzlXxDFbmHI73CI6tqzSZv5NEc4jxifiIjP1yK7YirNRkWtm
K4u1d1x0zvrf1Qill3t91Y2Abevp+GrbtHmT/6a6l3JiEe5XmKwRU377YQjY1H7dJukddztuzTdp
GtFxjYq6UzX5UQT9p9n4C3qtogEAZRaGmkHVjqkGU2Wyil+YRVzPEaOHXMhJZBVAz/9p3wqW/8jL
gOkfVxHM428+oK5Kzxv1AyRQMj3vQV0GA4qlpZFYecjVDQMJXbhzTxWY8MiVQpjagzydkR1H8jlf
We4KQcz4R8KkRRwZGFQ7RE7Ye5J8PCCRPu6PEEOxeU3D9U410O1ObhMvGmO/EGsISY14PMBkGcC/
UJCxMmu1A1NrrPA4Efk7fr/sFkukdNWCZDX6h4UHD1sE9eQpsVqhjqaJnt8GurbkfFmw2oujXsCm
34isER5JZ1eAnd3caVx+Hk7nj3RmhNRrLOqZlODNvvFVFdbWghOhStjMH4MJZD9IAvqGv9NpLCVp
TqKgkBlaBkB0y4EdIL818GmZD4uAMxJn5zFKOv3D60XAfINV8Nr71tgZ0e3FH9VOJdpwDWFQYCWv
fZm8gRxugZYsWo15G9pEncWdpQQBZdqUkJtLVPr6LHNv3lr++D2+FBDLmHg5JHsyk83VkdzfrB1a
05x83EfV8PpJY9oxKl8ybDMWwom6/5UAuJyzCRdnBJK7keRWJc1VdveDhtjc55gJJGgBYS5eLee3
fNnkl2vAYPC1GJ4kbl7f/4o/6NqUObEMWXR4wkojaO6cgXc1WTdei0rPHdY/4Uzv6T5OOctMwDDk
+sqX3JssN3NCaAxKpjfstm4Y8QLeg3oWtZD41piIt8Zn50a7teYdK8/B62hTocbFkagJT1Z6YWBB
9M+qQAlTCMlFDzQckR03I9zHBPITQMwVwrGDjJQvFleJEMRAlCO6J1/2uMpkNPXzbYaridEfnPIB
B8Ad4gbqJgV3NNUpGTzBz61uHMRiqdWiS7lnbkC4HxdLvgvfSrtJ5Qa7nG4BWRMTCOk5IL1zzsaC
CLY03PuX7ngWjRo8FAtmUJPxJN7d8Q3DxZ0B7ePkpmjpo7DGv/1c0+tfPli5VEht28gH8Ho68ba7
4WNwa9+QL9M9nzCz5Ld5YHD7ANfP/B+DhbKL3SjKi++eJmamVxPwoJ5KhUHSFeD50RToKdqx5yXU
ouM3tdAv4XudrCTyj1lQvB5WnrQJEZevu4gcmSuo//2yUGhi2VvP5OkKMjhij0clgdhrsq4XGUZQ
fkxKhr3k6Ae7g7nC7O0v9FfGXvYi6PHptrhBY2GQw+QNfCcxLIvhQKiG3P5kenoaA+bz90DLZCli
XE3asGvH959yCVsO0+iSzhAQiM3JQFOGgtVt3hNiRQ+R6uKtNBywYPQJqMxJUQaw1uuYMwBouRTC
qi1goj+7fd2rjSVRB0NAUOLKMZn1P5e1qutAoaxhUT36Q6zfCdQOO6ebufsbvyscQiUP2xKwPuHk
DVqVsp2x2jZMQaafmqfmyWxTqJm7CBb8Ba3u4LvFSnlJP9YKHLp3TQlD0s+0r+L6pQb3SigGYTt/
AhY3EfWPEde9pYVG3aK2x3u2EAbJ8uxn3L0mqXsmuVbdR0mseLk7Nhgz/bNnR8+fTWWYg3KX9U7n
fI+uU0vpBzq/vwbcTpb9WLu0wsHiFQouqbaOteVxHafyOPrYATjSJ83nq8ZGiTmnTf9gG6cZ/gH/
c/ENT2zNAU7+Y8+Kut76MX83ijGL/KQnjx0nGt5Da7SS0kWrblaW9iUOllCeIutIehGbf8xe+wMg
jn8jyUcvTxzBaVq5lfoTITg9PJhiO2JfNoTxOCXhMbC40ItoWIoUiiPG+RtLXglz/DBKsAaNwtKN
G2bjaGAS7K5mnS4WtCA5s+xPmbvMqmosxtp79zZW3IeKD5NSaTYEj3QElbmW3380NP5SfWU0VE1/
EgpDHARUqNm3M1JBMlYU4F6VEOSpZ3q8pc6A6W2qv5KIJLqIl4Ho8nGR++JkK0JyX9+A7k3uZUnh
aNOlRqzVN2Yx4TFcBmoKqGeSK0THLfqWFeoIUBPIpGRkx5x4HORMPCiVT01yLgNUZuAqNWxCCMyq
4HWIBF9NFqWaGj1oMmwGh/Z+cKzFmCo4FCnLFt0b+6iwh3r79hx/49h7njZ9KdL8PGcSXaI2Rr0m
9O7+6mYizJPk9T+JEaeBo3YxR+cRuzOYuzPK2bYwsok5ZVc6vH8lMcJD8QRQjGANJMR5+z4tLZ03
hQZvgGVSnrNlFm+rq7IMGRT8O+rNEMtJ2zMgyXtrQHW+sZbZyV9sPMEAR0T9usCSFA54Zp/lLitS
WS2okRqQGZ8mdWHYgazVfRT+VrHP0FcSmMggmN59p60CJAknNK/29SN/88ZCKHxxkxlpCSYsCA4t
z70ySrbn1S3KdcFmfZnEt9EICTpGay1+EfTlvDu2K0Pyjk+l18D9NRpm8CfocPL3socy/2iLzP4+
aycDCIkiZB7Hw6+NmM/tGDBA442vryb+SGJqxSQw5HFyNq9kURqas6uhqDptySKppnUtKYUPzl3j
9Ss7Hc+v0p4Tl26Yt6wM1ns/Evw072OHmhCP72sGCy90MIlguPyEdhovzFRGSxLPAJuLYDZ9JsTn
rfHmqF2jLzF0lJqQAuh142SSYHKN073uuI1OqIQb6ShR8+8VJaoCDOXCXRkIsm1SDTK01qmjkYTQ
ToN7VL+PeGdlhAgVde5kk4AhOfhrZ46ul0l/Y3vh1typjdDyDKfw+ydhhxKs9PZsqSCYsvrqyzeb
SDdGpjTJQS2f6CnNVjGfTTJZbx38A6Pnch6D9VLQSAc1fXvjSHDTcxxfi9JXliphwCgZ44czcHUY
xh4EpZr2KJ2n0ZA6b7oTEUR5MBJ85iC+d6BxqSW+52m7mAeOQ/7V1bnXE3PQvQrSHJUbgEPjtpqG
6iu9D8giF06QgQn7EJvm6ToZqnYCF0kgCh4Y2VY8R4rG8zrQd3CT143e0TntMv6qmO9iCVcZb3gL
KvHaL8bVfYiqkgnKs8EPnwpkePzS60O7Qn92DICUtbmQdWyJSwyBYe4pInyqrOvrwD2LC4emdJqF
xvVL6hk2mTeE8wtzimfi6yyyLvKDtMlN542HneVW35RKhU3NrTZhVh8Qc1t0WR14U3OY+3j1MCF4
CCZT/0dZpSuvkijbQ0v6bFo2xnjOb6enKbbI3TfaH+21ry//aHEQkI2gEhPW/1wPCgcPjlWx2p6H
Fe8WscNkPi3+GCe5OQjml9zk79FvGeQHSg4u/XsnxvS6U7BRgS0wddyU2npVpThy7fDG1p57mLGz
uFoj1uZ+mopsLijEkpA4iIuP0gQg2NW/O3LVuX92xDC7GMLWW0v5DpMq5q5v24est2wcRIedyV30
xhPBgfoYpJBQgkLjLvKzeiUOhHEYoJVvRO+Z8jYzQXO3GGX0qvyVQHNP5V5Tvy9Fyb1pDX86hP66
87dOBZXKoFDCMa5jX/QCJ1bD6FIWj18X22EnIPC+/e6ANkKcCJ8Jrmz8shJidahW82PmibWscfRG
TSWMnWndH4F3Tjc9dywDYjSUJqLlpc2UvelOWv6XkyHOYAsbtdd7GT+3U+cMUHbSQMLfeGI96HNZ
eDWdhbMJzw6lyOSz40vezzjT5Eh65h4JmFqL74T3xsKrnM9baN5acn7pTR19/NvF7rmkHq0aKkXi
hS3Ff4702dxqx0PFYnv/UI0rEbEaA0YxqXEP0/pFaSkWN6USr1uVZD5K6r+pO+0G1nSYmEEbEGaH
fj1XJte7wQFN72F1ozG6LShpbCa7h6S3SexnyuP8UDstne4YUmgGxJDPqULTJG+iu5kUW/krTKn0
42dgW6Qc1xFSqVPARvric9N5GcnxjjBI7R39wFkVnm5wEY55Ot45LpWc+s8dGYFF8cyML+tALNRa
TMRTRm6hb/YbsXFMK/wdfD9ujs0hXivcpa6OR+ASk+kHsfBwhJ49f+Vi120/hNGuNnGs6BDeI0Kb
SyJSfrrcMsEh6pRTWOKUsrVexCMyjRvRTvqDWfa117Re4LHfUdlbcBhrFLFcoRAD66XHgwhVqCsL
JhSPN59/ze2nd4DCZECukVIIjoAE30OvUrkzrCHRqOM5s27i86n0axRKsThUv0bHi7kMg8OiuBAF
BliyJA/NgWAdajZK3m8RoDN4CCX7eKyAKKTFGaiMA7kf9dhPqXg2cXBiJUiz+q0R3qak99sCZo2u
nt/jS9arH4DgoXdWCs9smCOxUPjPZgQSWfDvziLsoijkZdi7QLK0iA2jK4bh8a10l2Jcpbc4cjsl
kbN6B+34V/zL7YWGlAi8DSGBiIGJ/MIKUGl9d6ol39P3xUNzrZAY/Tdw4Efcm/TXQHSWi8nlO8l0
QrTBllxicXJ3JtlKr9+aoamdbv9ZGn/u0YbGhTMWIIRKPw3E9m61hNB4bTxSWDehDVrRL9JVhJWt
eM4GMW2blxkmwDzZbn13ONyc1EsBH+DO16P4QdsvIJeNWCh6LTHTLOzQtGsRResL9dlh99sL5mKu
JkecrmbcZEZWK0trDPeSEu1y7UMwUxJ3hIUFwjNg464W+fTLLD2g+qsYGXlzc0XIXl+DdwMqjb7N
G0CPiHQ3BuqsVOp8UdGhelngPXBmaBy0xY2VGC1QlrG8H4V5IF5e41TQDXXnD6A1Axuxq0kXddWo
hqc56BjKYYlEUU7KGADSFdDeCBKwuWkqiX7YdW+lxfE9JJMbYjnd4p55TR9iKxieQf/tfXwVj+oT
53y7cAyks3AugdP+pbkKn23s6gJfI/StA8UwwS0WVPLa3P5RgrQkluAqfmXFfRcqkSugkPAb1m8m
EXtGUxp4MWyezXf4Um5HaKV2ZdDSEpHHq3APrzNshFfrU3lFQTHm+3eJBcFA8OaX4S4jvuT3/w7q
sAs6q812Y3fvrhwYVd+J1mBes3ltwHPBfNcqUnfyRw4zCGkHHzxij6WFBN1RBKzm6+y4s2TVtkAY
bUXbAGG1TwWx/lA9RvLhr3cTy9WyHY7RI535u0cNFseeYT9rCvzUYHUcukCwX6QuOmidC7oeFTzA
8KM/gp9v7HzA4IgtZtsBig7jY4oRq9prrlObnhqQgNQTyAIhJtitMc8VGL2kDcmOyP0+aMF2iyAM
TqzL4DwbnFsl6l2R5+7nuCfsEMXjtelhzL5Fa/Mzf5QcZ/MI77rXDfBWgt95/8shZDdmoje/uBRp
8ADmGGUZJqV+lUX6bcMsasGHbP8A/h1/H2+AnXTKioPRr/T/QFjVL5acwQI5XEMsUQkbYRwEQWIz
CxdagW8XOon7be3Wj1QMqu/W8rFmqNrUFIawWjhlLVd9qBAOY2VCkUM3NX3fWW+ivA4w0AH9Yqeb
nv9yaqyhd7uPKs0G+C6seJwR+s4E84XopOL1/u2By6/pY0FCY14IumZG4VmcTygo2FDHTyMlUTpa
vtDDdwRDGU+RCqleyzN2tE0NEGlexkD6FVSwplhHVf89+wlSp5TfspCowHpTvf4Ia/+3b2MHxpUy
E3+QdFhiw1G7w1iIzz7tYy4Q0S6tEdlPcEBbGxdfFBuOQJJj2y38i3mSe8kuZGvKF8nKDZY76eaw
7oYwNh/Rai4bIi0eHGs2GV47mUFf5kH3cgxpU15R6CiTVlvkjoE/Q1Ca/5hO2ox/jolFDkOQjhMi
Kb1634SJmPQO6IRZ2yKpFYValtJIRs98dPEsykU4aPNP8VHAHdZkOy58LK/VfnaRLaWuEmh+mvqp
xx5TktLzG8Lm1rVVpVx4NfvEl3aOy02DnlCVkuQBZTmbGNtRbIgZ2yD1QvsYN4pxc8AyD1ZUvWlG
VoP0r3zX20ugZH0tF0MuP0VcopBq0/bTHPOMqmxuObg2w75mFLNR4W2lSU6uF8lkq83MqPxvuIZY
3WigsIQuizS2ZiNZ+XSTrPKkyKo8krpmbOae1EeKjv5XHX50V5dKLEKtwx27BpDcsoUJTKMWct4s
luhWxtw3Hm3F92Mam+fAqFKisNIWaSvvDyLxU89ZvWZBvPclN+LouVIZ9/ZaJmxa4z7Szv6tcur1
BoF0ootSVt3JbPJ9lOqjctjvs+7D+U+QbMT0iLRFHyLtOvs0e1VqpurIEugNGBWJ+T16D50UYu+o
7ZtRbOs7Qyc4jILiVxak5Jz3oijKhXIla449TfO7zdQykEOWun7ehOJWGgUbC8x9cD1viOopBi6Z
wQnbUpgRn4YTF51rattw4J5f1gXpOSa9EdI3uCP3dNUh6K9I7BYPbBL7MHah2B9ZIhnw1mlTc5ap
GLTmSJLC3x0/BKRN7DGAwTQXFUcTXhaxyVJ/PjRpMbJ5vjfQppRbhxUz0RzBimA5KZQA1axRkyiM
jxcs6hpQOB5ScRhHjmDFGGPeHZiPg5FaCZ/1fBAjjSlCMdyDesQRAzzPCf9pd3cBBOYKMEAndSQb
a8/vninZKsgrHQYUPelPjw56V1BwIcJt+OtZzqJ1Zx2uQWmpRkwgOXm12ga65bP5+fCmhkbgY8di
g0YhMY/coMxbANAWQKJPHcJIjnEmzCb4taPJKSIsZMWlPvmAdDPWEQAVo+Oxo28dLLyimqbHzPBp
TBtkZwmhOBaxD7khh7nqndCOKAcSCaLyUe0CSN1zWr8z4PyrSYywcQyZPsT8PDteSjJdXu1NMs+f
acooGFoHd1MDxM5WMCZctr1UKU7WLPUiHGdTPEIXUyLBvhts0k/oQwkhmiv/0VaeQXbYGscDj0PO
ts7cIoCrDhPeBtOfGGwPxz6gjLVrXAyosCGBP0TK2fEVpWAQSk0XhG6BfYw0physKowWmdYZiSWy
4+vzXkuE2r8MCS7ahsjaCiy0g20Dczzr42IQNMWgoh1Lf/KBa+b42/aukNZ+vB61kvlSUBdG0hkf
z8T1MhA/VGfiMKO05kJzB5tdL6QVDhgRrxW14guyuzl3QeXlzVb274wdQE+xNpFLhUywctnN0Kew
0QobXWZE7wr88o+ZyOBI+xM0pN7tNUPLGoO56tR8snZTC73i8zjzvV5W1oxyfS8rsCkif4JRxCft
yAJVNzesw1oBM3r5SM6j+Ao0X2SiyyyFF9LdM9LPDyD8L6+e0aqjgzFY9N+2bxoeJoz5X6Yjh+ZX
y9ETJRwbGhsJDXTRfkSaYhbe/kKaD/EaCaMC2HDBVFiuAcxmmNlI7WAikkaGZONlp+lhP4YpZV2s
8jSTuOyyMkbYR/bfkCNTAmUyr9dDSqzau0YRewoL6po3aPOSweeGiZ72l9jTSDdjFU70YSheauq7
arv1rHa2h9n0kNa7O0DjFAEj43ROqkxjYwFk0ondtHZqZ5KifnYw//Ezl7Demlx5qoauDkIKTvMa
kbhmKiK1SicVyDTAKkbsrUPRqqa97LXktWvCQeGk5o8E+A4Tnlf93r99+ga+REYINNLQcGRoy//n
Ee/R/GjfiDZWbXFQHLBKYaxn2PONQIgezQacJwPpA/kNle5WapO+je4cEH1/kIw5n/YIu/0Io230
HkDGrsE6Fufz16EnXysrWkx7AeNn/b0yXNqBXPYHyGd2O9EOPY4xWSWuzcfgT1lScNltX9peN3yG
yLoNPoZGtI9wgCJB51S9VVp/u64vWcR+iQaRR83fEZSB8xIJvWkUZDWrAGXgDYrbMRdeFHVqXb2H
bfU7FZhleyWnZUvcw9n/nyBcdZ8KTEFgCcwXuiL0/ojFEN1IzjZ675lM4amcCps2lcA6rWB1bRQ8
Ra3yXt1FzXghlWlAXaJLrJNTMeYcxbLLGUiAlDFHjNfijPCKCzKYAvG/CT2apX8fLUe3/ljCjdOU
MRdV2J6lXUngcpkF9TRPD7EkwV4qcDSHyYoftkb3C1G55OQl7KyQi21hIN32coPS9FPVBNByxBOV
YhEW6eTi3wxr+PhRNiHRlCS8+QsEY7gUbq3c2jcPGCsx149EzspgeoWIzKUTDQC5kMRM2UEDJtGk
czvcCk1H7dym1094MWG+Lb4a/nffkWiqpRpBIm/GCqFtbM6X3qs/LFhc39T8qBU7zmQVcJf1BNDJ
hI/VoXRAbxjIXnC37dw0jgh/s/99hb8zSBQ0gKxZMYP5+aWTn9xJYr4nnyPXEIws4en2LIBbHzc0
AHcb3ggWx5F9Of6LZTux+0sOsZSnMr6BJi7RTVZGGOs+ed0dCgPKajRO1p+cPVm5UTcrfx/To4Au
3IRkkpwBryPnSZSZRO96DBrGjrkC+WC7L+/x/m5xXi2Q9KwEJRara3+UtJwfXjTA8WZzy0rRVlxd
6QnD4mLA6v714Lw/PK5WsDD3HeLPLKxZrxcOwMhSRSnrBiAuJ6mrWDNPR1+8UWS9LB3O12v/zgnd
yVESExrGcne5XOkKKLjNvq1xOfdWiXCJ3WbDO+L6WICqq4NQuWiWTZ45sx6IxU8k8talNT5Hk1aT
LsZJ4n9Ry713MqJgNWlal5dceHnF1iB7NrvukfBy9rPNGc6OLkrxWHKwrNrWUK20FFjsUOnRJIxL
rjnPx0fyUvpJAyWcVJXYL+C2mPFPJgd0Cu4B6yTCExd1jA8FV4dOcT7SQf9LjqB1uizdXI5nrZvi
CKarQZsI/1LXYMGY3Nl4HXz+6zJwURJPbF3l3MkNsr4p6CxSEwMtJfgSdCaDB9kash7UXnt6w/Xf
r51ZmRHS+s+vUwZ4UwfVb6x4Yk4s6dvUcTF2t8jRZT24rOqiLA9O0kebp9HTB6mWugq4JBhX7anD
ge+1RlhKsWBimue7aO+JMe2TElwkATT1lEN0jwVbXXWXffpI12oQaxNQ6Uz6sCrLAnVQ4X0K9rvy
9JdHR+9tutdOMk/hGIkLHpZuiy9uzyuJjaOrhuTQFS/5K7Lp8X8ndgBwanDQe5dXIbclvwQJ9Svw
UW2gi8OCvLOj4iAs5p9PI6PW4Q0Qv2Ky1Jq0DODmtEGWBEFAigBnA2pKfNqFSYNPPI4545gFrBWr
BAfUazQ1HT6WOD2BVmN8tninrhSXUO1Ziy12nR2eSD0t3QkNwDUE3m0vPT7dWUToGHnaJFmfYN0K
BVKATElxov333jQTnZRlEECMo8delzqt1nec0CoOpD6NAuQL7nFoL1wGwkFj8SUxWGOmpwDiKnCX
G7xx+WGtoAP7DUL8Ou+sdF9vZYGGxp8QKIYziuXCd2K6ZVNbkc5TzpQV4TZrQCcbQL2nqM5Y8vRi
573/og5eqpTMQJvHWbPOHWEF1EcqKYPK6vjsMLxX65lIIoLgx0cnvGMJoSN5+cnVqV2h1/vMx+Db
cel/u4sl3nLiO/x+bpm1usm1zx0cjShxdh5tR5DnA2FADP8jW0S1FAGLtREO0XgTrIlLdvppWSXq
hk25MVkHVSjabUpwL6tUyN1DXg7+4glAL2jhW6m91ITgx/V/bt0PR/JBR9ydWmcVO7LtBPAX+5zh
J2RKyzPfS/c/EcodUNLXsFdsJvk2tHNA3r7zQJ5D4ZEfExuIC0W6bDNOOB5hZTPMcespyQpeZXV0
qqbDV5pYuVfo3AzeACulfmc8jL4c4NG5nKbYouHXuoHly0RJjNqJ3l7BwBmx/eZU0D2K65NoAs7I
+hZZd2AgKLB8wIRK5oN46vqA1kbjdTRumQbA6cOgDJaFvwVD2R058y1auvA/me57yIi5DGv58ORP
Eab9FWLHmxKsmVWuW/5RV/xftewmpy4Uda7UoAgwpgAMjtsH9YSXBh96gt5PAq7y2S/ub09TW5z/
CS+qf8/MfXkeRtCgsfDUDbGpnIffcj9HY67Sm0VaVhE0cblnqNYWMZwTXBDHdgPniqQ/QdYyYKn4
72/39WQBPxjklOa53SoVzyyFjArqQVQPX2aU6/Im5d3zlEH22P0U9ksWHOIXRmMoeXzSb9myuhxd
vcsrH/9LVVeNR1vk8aKcPD9sMjZ6ngTxOTdIuJW3HDW9F9QOxm5tmYrs00JgUiT5dU4gK4uCO3jK
QgcpFbehgTuCu4w4DyASCeCWc291HzDbHTUy13tpLzIWMYn7wlvOyRQXj+yLnVoY4aMuwherhmZw
olmj/57yin7mQpBHdfJqSzyCGrAC4FB4om7wAL/yhDX+qRp64Ugy4z2W/Hm/fYDqgAEEg7NptJk7
CvkZU0SY1T3UdYrCwFT+61n4Ch/+Rn8zdu8l6nZHu/kGyA9RFG5UgjA0uxNaeJft0INXSWYN5kaw
nlHyQcuvSyF7DLhy9X3xeM1jQfQPz4hZRpzZ1DCOv0lEEwPOe165S6dD47FO1xkS25FqDDhEBrmC
rCIbz9Tr5xJHFBqLjL3fpko8ezs+JG+OZ1XXa+535AeDM2knuOIPrC4ap9Bn4UdCvzHeO5YFkDJB
6iNe72pPRdmyU4T61BNOTBuP68jg27ty8jLCwUpYRM3a3ehPLLfgW3fvGUr9gqhi5Er5MR8YiHLH
y1AubUdhN4Nxu2adF2mSICndDOSrHHW1X7rx1jmhrojQTFLn+zh1LxrmNom4qwCWQnOoqvy7tsRb
wOLMcmJjIpHACVmHkGch8PcYKJHYQ0Wpj9qxilzEknS0lRy0xSrlDFmbzy3Pqsgu4AMVuNsEoCpE
QOApw3NDqI2C8yoftXVdVSNUaYN+CJ70fs89n7WFEakLwySzXTW4rZmu8eDHX2Sl+V8Yziwooga4
3X5847RxXGJjo2Qpx1Y26XggOvJILKGtByWEFZGAr2XwA3wQroKeotlxFM5JasV8asb6bt0dkai+
YKQadzYRzoDLKP5aObHv+q06qoZUNmf7tJgaYSdSMISMY26D1OgsrbEKw8qHbM1mYbtOkhJTpELN
sQ/6NqPGONyQmGpEvMAY4tEVsDaBOhrfQPyqWhFUQj8jxL0C4NxzbyzZ24AWN/1Zxkx0eZG8DMIS
cZWNGEqWzW6+DbNfWu9kkPEnPKAxcNTfflorbtn2tRI0rpciw3qlKrrFEGCZdYAWxhofZd3cTDuX
SR14rUJa6SKbazQ1iZ5HN8U43Tci+RxWhEWbD9re1vu3v7E1jU0aPhE+AMCSD5x0tLYbHkD0Aj8n
Nn2S83aREhGUg35PI5vWPCrZIrW0NMwpO9Ulrp1J0iXGkwVc7v6Mrb81z5rv3w090ytoiQyoSPJt
ep4JQvrDjAxAn6wa4CzADpr5gRfiBkGrQOxL9xdiD+qxqBX1/XJjVbcQgiHAT6KILpdnkbNGgCpU
akMnEw4vl2r0JQk6q7iS5Xoj6YaFCZUa9j1VH/ssFXfriFIYuJpiZpBsHCOYu8DvedVy005E96aV
cEZEKJS7MiHJ37a3V0lHF2vI1hWmMmw9HuJIIjXE4ROdlBV1pyOKBKD0ps0DTR3NChNTNP5lRdZ9
6sUgL1vYe0Wk1AsTGsn4LxQoiR67ap+Ip0UjHBDZxcxtWXk7i4rHmnS7sWvt1abrX+VJCKNo370z
bEWq9h0BVDvj8F/nZm0XEZwdDmW2hyBYQFihmGgLZs32nSzEngVw99qDNHdzu4T1hqjpKqb56gPb
fs355JV23AYb/sT0Sk+U4OUrWD4WHASQuwqZcRuLasd4xh8QpOOybebU0zCmhNcgawtXQD+ZHbrw
6HxEJYRVoGjOj5vEs5Lo7DtVGv1F8YzefW6AAdIN/2n1lAE9kbxgkcMdP+4tTFlUN3X/iUhpUK/q
ZgBpSxoarRbjOYpXxMjtDMgiCFpABg6fj/J85ByxzFHamQBuw0gpHSDbLosqn/EIUDZXfUuOX5GA
Liip9J7GqjhMe4q7v4536z9nRx9PJqucgm4beKlOSguw2qCUEfal2FzgS6RRy43K6ZLWP9z+W2I/
CUaHsTlm/kuOirIRi8N9RWxdH7RNG/e2h9eskl91w+9c9bSapBGnWmaT7Ga7k0Dbq18GaEPk8vGu
DqIWCMjPwSIEMXKuQDwA4vv8Bko5xU3lacAJhmpqwwKVv34UvI20h0s30JDrsvZ9h+KJkiFosgUx
6sAjW2W0SXX8iF9LIvjRDVZ5tJCFInRGN7z5eGPe/TBj1OQ8LPJjEVy6hmATLxA4Rkl8byFfxbRq
gG6W5SXbD5hj+gI6aC6yM0A2KO84JnE5jBr7YcJcBaHGwM7mcRGzK58Pl7L0u033ebIfzQHDfn57
jm4pIuC+eL8BaXGQo9wP4ugiFhYvEtjJwNCzRhqEQzkTdgh/oxCvI5rXRjf5siruhhJgX4R0sawD
Htq9kq2EqZz2rgQ+74qbGYAcc3PADiLAGY5/TZomikzT/H8SNJSlCTi/nOLGBUgbRyy7QeLFTEZM
sobBguOvAP243H6o8NtqTN/VmiciYuR/ooB3p1T9kEQDs7MG5rMlRt+0VsMyerDzaT0iiBZTqroR
YHGGjcFbkQEuPkyGURfB8fthZ4dbC3VQZo1gD8T6o4QYgn72w8Bv470ZnvALNa1zxhLkL3jRIsM/
ojDZNkrrWKreOJnunD7EBLRzkIpwJAR0yFh27MYkXXcWvWEXWL3/zMnYyN+T2UzzWSR9uZM4K+2R
/L/gYwYlwcLmFF3kZ/nLhOsDAvmPuLqoUUW9kZC6xH15dtIbt54tID9gYe4DjPgCUn3GDLD2VJjQ
ql+NevuVd9dWwBgi5K/kkHbirlHbXepCTZFOnQZAYLPMCsxiaUVMZkhdkgMn2e4vOmw2KNGoIlj3
UKUzuhr1Dk3KCSMsafOrTlfJqCos4XPWNPJG/hCYz2zg2CtTqNRbG4G33QEIm2OYsqkxVYjB0ial
Fsa6ptM5tejjgorim41gXpIukZ+q3Oj+12sGZ+PtIHJZorNsdEfob3gXwqROiBY0ZPPuBuFeP6pd
qJXZWZePDhF07EAkAyRtuIUPIEY+KUAyLG0E1SRumb5aJdKcXLO6ZLaSrkvYbBU+zrCExW3i0PVb
DJWUTOTw+mpDMU06zgajDg19f+TKm/tal6gY8U5Oc+f34jDVuqKMlfpcxU7HgdfsTxGtAFk5tPp7
YMZZV1h2y0USR49jTqX6/96qFSoBdJ1OaahLpWCW/alGOtVGf5JetGxDyXSgN4iONvFrVzeiCejx
J5HYbW8hCb2xydbep2wvUFldtXyU2FHJSmhMwtjbf5qDAbBKMpG1V0jvi/RvlkC3goeW9QgB81FJ
OJzeRifrUhnX3DHONzLQMW7qnTpUDNTGP9aGaRDUu0lDW5A6jO4Ze4nYPPYQk9TWWjgj2/BYobt5
irYO+R41UC1qUXtDs4TJCWd/djuTERwsVU2jUDJzxkt7dvCNfo+miUlKh5mL4BeBVtPpe3QNC/0U
MoFRxD8m1a1qax7DTzxJze5FUpBsmbNvy/TXcGxRzyAnwo9U7w+LaOmVCUcNULhjFG2ZsG7L66/a
+MlveaJkX/S1RLtJy//ZnEzdR8aYx4NuPfK0h0q227scMUfEYxg4xrokzG4gqhEjsWyhzpxGcW2O
OOwdXmWSPj9146VSw5Ssh4YV0NI3Xj8oS5hoeVFFIGQeVchSa99KlM/NJPEzVa2Du2X9xoF5CyQC
DVnIy12ARmXrAM9/pTYFwPOy6lZaPUiSn93UBOBTi62D62Y0bM1m18uhNJCHGSTjvJ4Olcvpf1eX
WYNEQ4mOLlJ/E6A1P+OlvdJ2sCp2BhxqCMIFL9i+rYI4fagyaHFnHbmI4cxb5VsabZ//akKMmgwa
pPKDL/AWVsncnym0FJ8/j1YSd/a4URKmFISMPfTCIUjoUwXiP6/ojPUo+Z9ddLR+YzUsae7vk9td
tcYIItUSMieJU3gyj77sJCDsJEjdJKKZZ0BVKjQKltOxNtpJw7042EPPq7PfD1rnoK4O1HUMtUTz
6gvxUzONUB/SssTM1d+nOmxeBA0vzpQhR+ZnjkTmoCs71Zq6kQ1+3oNwT3GeutQbecCTGoAzT+Au
uE0RSFzRZXl8np2rsGiGZtTdkchIfV6eyJ+9BfpYPg492fpds505GhKzID72A1z1Pm9oxNCQwVJ5
xFBNG8IYVIH1ZIPR1kz+rYgtyk1TGyI6KfI2E4ImVHo110dA2NehTO5KeXR/3N5d5dXrkS+w0L/B
uAyzvkL9k/nuu5PdZNXqRZzn27ivpVUlrNn8CJrbx599DM/RYFgKkVzJrnqLr/vssr9pAwu/T9BG
v5EeN406KayHYOmrXLH7sLcvspqXgO29wI3bJJhn/WSLBM2dJU8Md4UV+6Oncu0DZC96ttSbNiUb
ZIlUzWBv9hdpFM1DP33t6ChXYX0wFGTMwzsixwEMS+1v7kJT2PRcQK6AP3Dlzcx5EkVwj6CuTL5d
YisXreArhtiG8l1hK/5lSm8WErUAHy/NmqQ0KWER7PJLMdlANDAQiTPJhfU/5exFGQKUXK3h2goL
8nhle8cR+a8Yy1+axnTnJ24OrpAMpLj50gwYkYOUj8+vaL+oSgZu+3G9bN5Y8TGgmJ+4g7mZp40N
5yVTeh++4oxzNOD0GB14oFdVjKFXxJpYkih7aBJty+jnjcn9eE2+Hc4ePbLrvzxkOxHfFpK3krGU
NFkjGaPMqOOGDhMJLwhlzuVbzRn5BL29f5b6VqXDiC8mc2VIysqVfy03VKuG0I1LsXc8MQz/ayr4
3ZglQHaL5kYq8z7zjMbNoDj68byiikagtWubrS1Bnl9MHs399VIOI+y6Kv2/NkSZC1NA1scfcEWQ
OeB9trrusJjk5audwPzYjg04moHpOF9koUE5nXf+5a6/YQ7DslbhwAQIASiluFg7yTpGjMZVZ3Z9
Ztv3tEiaZd2lg+r+7S7ZKqFhUDdSPp5J4opUf6oPDqL1p7cLKA4d81KXjYPmR7ws5jIGlXR7Vwwh
Li4dF7N50LFL5Zgz9B7T23OgenNgj0bcqna+SzT/Sr9yrb76jhbhjWJxrOm8A+mFShlipMwqGGwt
dzkbMBb3FX17MbcNax2iG8TI4sOVxlVh/sTmU9N1LjKpZQl8/M4UG14XIJVkj3g2uoZPT2BQeiuN
1f2uvrreSmmQnnk1wJQUYarlFd2WaU2Wygw0eRmbe1XP0bohcda3gXOZWXchuDN4ec1U22iV3crU
ZZDSjINgHgaSjOUyuueWeUGhBrIQ2eo33HYehxaD6AW2gNfdSlXxBWza7gVxxpEPhB51RyEovyD0
FAfEAJhiJOnY3l8WCbL5QTnlXqNts36U9onbwO/XUNCt5kyNUSVcPhEZHf4mbkX5uNjtVlD2+/ry
APNoPb0gFeco4nfjV0rcMUPH/yerHzvRVUI6m6tkvWXo5l1EWiz+3WxAjLaTs3iWcqeipqFHfeo6
/btF7NZKRLzkyl0CJZArU+UpVAmUamPbG/eF7mMm1a11U9oxesgul3MaBPr6DsSHK2hhojygfqgP
J484bMwgsIiB4K50Uh+iFn0IRmyuy4BIVdayUmvO7JSoAGInbQ0EDFfIq5iu80xPsMAa6n4/dK1J
o9LaVrHa770ApKLT2yKQ75bwAKAh+prTA1XpqxgtN48oY5Gr1NGN1hOoaqYYed8ThU0EgNQL6ULT
8yIsrKn8FbB2Qv2yOOnsqOSOImGbFvALBkHKIf3XM9h6hVD7JTGm7ExD1V1gGjEJg5W6IVh2Oq5X
Ptb+cex7Bdvj4uvVl/AnHf7TCm5e7Dyj1WHkUJ7gCpwp2AjmHXF9PBKrBqO6vY0u916aszZq+TBL
E5T+RIhnL35iFAZzviW7GQqZggdd0v+av2BIkmA/ieuqAO0hnL+q/xRUc7kKpvYX3BPhobz8XK2j
ffVN2Bw2hANn1c5isOgI/vrSqIVlP3X9WaUhkMextoAbmIGUNm6GtrarbIt7kIhFed+cNhSFe1z8
Xm/tbraW5yqqJk+GBmYSuOWVVqrGgFKgom46SFJEZpz0oH4PtN3Yc+CZQBT5aSikupXBBX7nQWnB
jvHH85PyfbGv3b4jwn611BZ32/3NrC9NdrCumu8hHSdtuivcNigz046gTNeVpVI7UDtC/S4dmT7x
WF7eNXMYQl0UffBAzBw986oIKhFBvo1K4enRH1AkJ+iY1MtluazmaKQ6gfILI3WQbSyXmK0qxNgO
70H7m34gMV0rXiXohtUexYgLsuMrU0YmGe2t8SsAsk0pln+gmcbgx62HYSXZXV4t4CiQVQ3aa0Fa
eMnLNHvQtmIYS3XLSgA4CO00r+IgJZM3a/WoHf9JAY7Y2gnsP9AENbYe9NfiHCve+EgJO6BYd7Hd
mHFbHqYLT1uIF6TYbKqrqOMpskSxIARy9+RwthoTodpMB6jLFDC+KY1zwmHK1UI664TDCiY53msK
ciziiVXWck10XmD1BbeMK6KBHlTnVYQ+7e31EXsUnWjDRMK8vBDeBGee5F+yh7VMpWRqURAcGHCt
KOGpQF3cRF118Kt4K6oZ7bNoRrd3RUJ8/Sl/foWNkQgTnCnTGsp2zzEwRCJ5T0ixOCT0vQ3McDOo
dXntIeywyvLpyDPp/2Bi3CwkptJjzXgRfFmO8hNwAN5ab+8xncGnRUrtg1CFgs3qYeWpi3nIOaey
xZLgfcfauDsYcH4VAt24jKKVLyzGe4PRbbWinnX3nR++8u9Mq4oOrncm+/tWTgmLY6ahCaCaxM2V
CtrBWFzWSodfbRdkZjuhseFj0h7vLYvA52SFEXDOon+BZwSjA5VuO6U1Nhak3ETnemv+dPHu04ie
Rvg5yqL4n55AS7X73XfIrBwFUe8QYhIi4SiY7x94YDLGDG14uSTOVJ7Df6lpWwSlJVLC5A/jfkMX
vs2W0rN/aOimmEIe9yKQE08brTwbdthDQVXS2Zoe8ef6m0KLtk5utBIF5GwiPrzNVNuDJlRvSZPY
3mlR+jijzuUr3qhQsTSGRFkHHn6EyljnUhEmexEtJGYPSkdrZTx+/ZAmdKzbucvfYIA0shXIfiTt
CriHPdVzkx1JyQ3VIPB2GZwjvOeQuQD5hvIcgiSXI9+i4zA2krolzTBpuZGqnn+92RfG7mvH2YSf
ttNrtb6q98aNBqgQ2e/5DwG7LHw7XN1C2Fkv7T8EbTWh54TEliY3grH6r+994mlPPFzQD5Yu5eR5
WgNIoUzdLSj1bboWwDSs4EwCOCeEtwartRjATyVemaWdtaKQ16LMfzVKiOMQmjIl3lACP84kL5gL
x0cRq7dBEEiRU2AtZDJSjA3CBRAk681Z/HDY5Zen2zIxKnojuBOepnVzB75+gtoqZxnJildiOAfR
5JcEdrKNbuMy2b9/mxgnw+4ckTD/jSOYi5sdZJgnTfc2SYyHaHusTx7PTt6JivFana+HkbJaQcJX
m25cG2Ii2jg3zG/bn7g1rbKvQwzFqL5Uo9+RsCbiWf3bF0qHF5tuF5bhZoQNzfDX1/WrKTCVcsct
lcW/NFJctKfeiL6Qo3HYFUuf7phMM7T4MhWD578eqEN0/nV1npYYrCDWwwdMXrOL1FFWrr4Tmypk
et722NSwEVD6P/eCsiOTG3w5EHLkyVGRtW7ZUlkPlCw0V8unX5A8dns7Gb/8r+3PWdXf9OpB4jEz
SD1FPt4lvO9surWSRyiaJVn2Ldv3D+fXWwYQjeyjpvRegLxFtOzL5e03WqQZEGqfbwWhhCblbiPJ
wD+u4USHr0va9yk4QZQ2hx2rflub9aFmMEfVezA+vSoo0DC2G31mU2tkKvhIJ2FkepP156uE2qgD
aYOOyOFNy8IqLIPpXuqEoBz2oEfsLb4b66ChHhy0mMX3yAHQrdMbuPE2kLVxOVf8vPh+e1lgsuk1
6j8G5ahYBVIAotZlVjjN0abWcOS4DtCBkPETVgw9IwSrep6c1Nr0e72sGAploXD6+TvCIwqdc+tM
3TLOdYLoMMbgBHUi2roz2vlOcosMMe2JCOF5ZzAIMNW6d6J5OVD21aE8F8Ch4otqH6+R7eV1YAvQ
AL7gIyTPC+1N/TWnk8esFr41uYH/xFJUXK03Gz3R5YTa8X2atuw179ptq2WxgiPg/7U0vJPXMLE+
NQu1HJNOwhZc56WRxSLrQy89+kTKD+DexTVVadb67O2iR/R+5l4guJ/NITQ+SlupcTxQs31CUhek
H3YRnCfhkSYo37/7oCtiDDJrlLWoCvybAgV+CO+Hlr0vBS3GGXoMH8wBdeAXlBRYGkCiGljFIojb
iHWePXypQQr1vPe86LWzb+tJlolUaFRmD/WraLgxriu8KNZsutW2LKbtteB00ru3owEnsYs5pnKR
cHcyOHEi/reOGc+sQ1b5ciyoyiwTVy0/1I/DkluDmp1jvB8qfXKjVTZ1yMXBMuWL9BBzSL6yRaOO
sQxe4lfhxmbjjq2tWPXX6GGNsV5Mtma5HhUVIXYhdjQbiSA51Zz6D7NOi5498k9K6EhHgGr7byPC
FyYZkTr0Ic8LTMJkylKxr/7sVHr/KOuu/dRuv7eTbJl05+Wewn5zUMQYwMGu06IUvF2AI6UGGXJE
yFSCPEtxDWbqk4L/Iw9eWyAjXHqqaFklaJNCUo5gQdcp5I8+fjLP3KVu/HAdNoALbkyE0cP24snI
4FXP/8FwR2Bi67UkkL4yvOhqrB3vkj9pBWgcjKXYmNBN+3mw2uKOj3QD7biqrtzGAWmDY8lQowZo
0JBf/FWx5l9eb19l6dv656U/lwNOAB6IXComVZ902VfAztEDMS0km9PwFM1kppnWMNuo9tsgFFKo
qtrM9yer8DA8KYzL8kc5ArfcAXA8fVaSakb9pjPsi4/RpcuoVHomazbEVGqEfjHVj01jSwae3CVU
7wPVCAW192s8oYJO791nBG+2HW1CbsP1oz+WpKgRQf1bzcjmtIqlYpRjtkwyDoEIL5pOkke4WbLG
51QFcH8sImzekw8Rbi4Pgz8GRsqY2VZzyAb4N06x7VmWBS1iUfFiKdrEFscUewXPaRQCKyt/yPld
0wxnsJkIfsqOAldddfXxiZ54+R6PjbgpoVUXRvYT6yHCkjvMrBpst3amjxJnyFvR8AJEE2EQ/P0A
NJgkKi8KNjtzQyKl8pJkgY+5Eo6BMN9rJAJounNuCBmGuasCvtmXcg2nVkl6mIN8VYCFHVITJmPx
tvHSpqXI8qf01LqYAnXCWs1KcK5KGFXyJYzE9+bF8BpDwCHWY/PNnKR3ouoXGD/KKtlqGNVwoGVF
QLVqYgUvhiDyENiE10dM+VvTvHHsuXzIeeJktPxE8o5nP49zqr5BUWPa2tkpswvXYXYFfFQIBqlo
eTvopl8q3IuR5F8MVZOfccPFySu+g3uq0hditZtpdaKgyIc0VyCvZFGprCVKhOrgzJg9FiRUktg2
KWSGotdUrp/RtDJjZN4EyA/I6M1oR7Q6cQKZH5a7RpKAb+FLhFf+iIUULyAcYHYISE4tP4RFSZrN
6F7sA8gyxsA+1Q0ahKCvmKyW3e7P0NIC1tM+hdoZfZLLFXdDPBxG4nbUKf0hqSAYox2fN1vJGpcP
dp7M8aMD7hI1/wD99dBf00t6/USoFCZx2T1zy2BPTxLI5QQpsgyl5UyaeVFggw5hx44JNYTFDDqP
9Gg9C0FWhJDMWbBA0AHl0/jGnE1EfuTNFBhsHTRY82U40ObBA/l/DEfAtrby7dRYBUq1UZYOr6CF
1hmF0cNAilCbGfwzLfdnP+Gdjfwp6KNMcpVOBnmj3mOwG5YB2G7ANx6Sx+IgtPyiHfF69AJYWDx/
BzAsDDg2yVN2HLWyXqEPjYIAw2zGbQ9RuhWGVQwRiCZzule5EVdxP+gd2i/4ORJGUnFAF/W5VvdD
EbyeXCKOf5IM/sXQVzXLzSmwJ2T9uP1lNsYPKk9YJRTJwODatmXTIsmc7xORDNmO7rhHlnGLavho
XA8kXyJKdVq0maNqPW1bs5x0t5E7q2L/ir6c/24vpU3Rg4MTnJCzRclirnrhh9WjsiY8s+TurZSe
9/b1EGo8xXwgcQ4x07idPGmnzNPc2QT5Mk5NnuCNzb3/lMH6SFKg/mdZMU3WeqaMAs+inNu5qxxq
4H561DyDdsiEnZRWFlO4jepaElx+LtyQx08Qfl2kCet0i3BTeSub0KUBgKpbNQ3o/F2RYPFMLpVl
DiY+wzMmVbS/eNyfrHgTkAXUYF0nk700/O5dJRFHy8CYkU+muO55CuoIlyLvjNMbR3KLQkpVe8i4
vGE+85nvGwyBezQCxCJKWnu/oMb25/bom/HgtFzp18rD2E2axqoUqvJWNyu7URurg2Yt65H+iZV6
gxbV89QaM8/BfU9xbB8OVJ2apwKFa/50elz2lewd7J+yVwb5kxEZOBgG8TTDJ/pUxP1MHaKfGIoV
HT+BSONBqMlcrnGVziOJP7AK44Ii9EaTPx3eEL2uXjtS/8UyoO9HLwUIzCpaIDBtDdgr55DIK2FQ
Pkv84DOu3DooMgYbLb8LhRzROnWSjoBdbmH8OfFo97bghIRmO8Dt3XEpoKN0nN6nvARIMIrB5fSD
Uvb0KB/AbHS9og48B/wLGZIR6hHndxnCzd6dFV73kwo+nzHPPB3a6Q6aoTSMkTFfTnAC9NF6Epiv
4/ZKpfhVvUgm4l0tdzf2BowDmy1DNHTUiZHvh8cuk5IY5KdUaogHuGvxqfoASHYGf1+T322GsuDM
2fg2EO6TMIuUuWaVUrl5KRfT7+E9xoItilfx3SirwawKIORYKZulObjkXbAuwlcQum19NYryWcxn
amqZAlE5g2aEMWKPF4jIM95572FoLcssFH/AfZJaLbhpT69lmYwXdu66CHrNn5ghbncyU5MAA+Do
rCdedouyeOdOglfYPz0B/lJw/VuIOMxRx0AxISJpeG1aZ0k4z29+ZG4Lwnn11axkDBhPt+2TU67P
xd0Am8pdkaoXuz7rvUsAs4GJW7LG/941Ktc2fvHtFJnclyP4w3KQhfFgzXMMk6fqyN8ZsfFe15iw
giEkB7L34yOrydO6MIYHM84mUuI05AaB37bc7XXIN7rk1geMo017kxs+V8dE0SqQmgGHNzXasCpV
4VAWMnFzMR14uY/FwycC7VGMJN27x5+org+x12N3uzHKd8BoetdDqaSnGgwpUa7sOWlZBNl5+WKn
963VimHG6/sJY0mc/holP30zDUVulXMR3ffVxOOqJLLguM1QaJHcHK3HlqRCM2+Eie04bibq5GKr
/oviqi2xTfgPR6LbZTA/PxNQaw4jVRdf6zXqf/+JyjEw5cH4xQLTfQqshnqYbot1jVlFQxutnSl0
vny0IimTI7s+J2T5lKmrsiq/VDVodDiPFWDjtB7hpg32xFDhQGP9VgA/HD/U/65tuV8ohFieQYdz
d2FUGL7+kmZ3EvsK1NSl9eurwrto8sx0vct6g4lGLtEDoj8t4eVEbdSTzaCQ+D8cGf8IRHmx/G0O
v1oZQTjLx8iXdI4Nmo4dglCrn0hfZzpuj3OTM2yImjzltpXBqCshXVGfLEKfVuFdHI8DQ1sQEvfd
EmmeE96LucWuQLsY7V0GLyTLeW5cJpTtKTIAiyEXICzUwUaxj71IZfXrkJnsX/+XU1hzguDr0Kx1
Kzaa+Dy9klPdAqSw8kNG9OzBIuONxQPMTRW88PDyaK7pGqRCKKPoPZFx41OPD+jftQ29Xju9OoBH
HL5KvXfcwGMKzmRU+mM/SF01ItYPLBjrr5VVZGZWKVkK0Mvw5Egk7cbCbX7AR8dPuYr3zNVxRwoa
tPp7XfHmmIbV+sXYYCgq/4rDFU92d+lvjmCup4Ls4IJM2S7hJL6THK1KPSnzk1hQJKvp2jRMdXFw
WAhzOUfAFCLdjLNd/xh5byop3bimnM/mlAeork5ual9fsEWVfXRxPfbP9o9KZkG6V/M5elPAKGoN
2pE9hgghJOMmjjj+/Nm61Sv0PuaQyWOw8DnuVtFUROqg7NAqa8vifGIU0M7o0qUo9p0tcLrs4Kox
c3/OgUux0o/rPhMb2UFxHR8KtsjbHQ8GINmaeI6xeJxAZOdkJ5O/bHYK1Y6RHI9nz6XB8jtv4ORE
7D568MxQEzd1+5rSZRQsUFxufomSAz1H/vxJueGCJ2DmCY3f4IuaNkf2bz1x8vzyDWMkuEJr8UjV
HblKtYzif/bIElOjFy2KCexp0qvR5TpEnGrjD5hpgaqY4TecNIkplM1B/dXFayb3b6bfayasDQCf
QZI0ixqTjDOTJTY7Rp5c9eGmVPjsg16JpldtslyXtgDbV/5rnx4X69KV/AZGgRgFXAgymaBhYXgL
eyISvTf1D4FVC9Y0TFxgRRKBOIwAHZN3lE2RKukT8Lx23z0IOfqLW0FgJJDNzIhs/DiD+PKagsec
loNT/TaoTedpc81IJBiDTohgpZg3U77OBtO1uhykTr27hZWV3OzUidB652fBjBMuO5iyDIKOUMux
Tjeo92TCGGSi8KGPrK2e1fg3fC5WbDfDW5g2xwXAL+9jczwlxUu6TN9JzcOl644CUECdLVmsTDuK
23UQZJmeOcKRUWMsvQYzmkHkfdBZmDN00vq56UwP7Lu9xnfc9ake+T55P2B38Hn/kBaDhAke/LXs
AQz2je54m5sT4THkOtyE8hUe/nKRCHp1YiYvMyTVvnG8x64j5Fh3/U5M8TJYiq+EMdzumN9Tz/o4
oChZUcIJbyVTsjcbUQjg+XRNbnIcYydKxbNiNstJHmnpcDs25lL1xTy3ZNbnpQQT8Z5VqXgo9YCR
ZxjYoZSrTn9Te7xFzr5tsBo43wspvV7elig+r9trGFsiXTv2HJQBNiUMjbWp3idz5vW1Hghe0rgl
nX4utNcPzB7SDcuyJZQYO2cM5RDpSF93w0FU8YrKQ0iuuFMFsiLFEB5DNUlZZPdvIHNZ3/Bh+WDi
Pgk0e0/a1VVhmoQVLimpfKR7n+BShYnqKM+RXxSAOBGrpYVSaboyyy6CMPsqyX9kTtPA3qQg8d1p
6ujUlp7zbKC6j5GO/3L14zjKg46dGHhvUtmhUjQvw5stX035kGN9NETaRrT0Vjn7Kbt6etRmboxG
6em4rvAs/qQo36hOu+99LnvSRnTnbklSlBRFVrAnIIvnrBTlHoRkScZoQ56eKT8zqYizvTVmXBot
1SNADNxcHF5OHG2f+7A6DRzJJQ6pKJ4AetzsbNXcu+40K73LBUgNsx5rPtdv3fWrrQF5JaDZnG6t
y33u2L/wUuBPmrtzDOPjnKyMUeCGruC1Aigx/3v4OH7py73TsV0QTBnvRnRLRGIrxPsBQnCsKDha
EHxFi3/7+9AcvudzDuonE4myOlKGSs43fvFVcAeb+eDi6HgJLo+Nhf/iDeQ2TCTnUuoK99aGj5X4
4xE31tE7zxzcKtw0w3b9dtGQJxdvqoEDE+U6Hxb68Clg55xjr25C6y0pRxaVLBTQKPlj2gcOK94Y
0K3ZDoBi77uT0Fp6GmSTXS/gCzRaYg3j86z/qgslMPhcgdrDfUWpFeDePTfx+a6ODybiQSaAvz8a
OP8aIrEHbqEIDjqWX5/txS+At5xs3cWc1i8dFu5fjHGMIKQ7XZ6Dq9S7ys1zDL2/hWCkno+dUbpX
67Eo4NH+caPN3X8TWQn87aDa44ba94fhVubm/2DiSfFrKhUTzOa4+Vjx7C1Q7KZDWgN2rPAPYOLK
x8Vwrg2M+iH3ntzo23+/8xB0et9F8OUzT39ej1wND5dVQuFRFWMy7tDYEgL+KLjVZFOBFMAP21Xt
VbApamxoOtxTAiG8yHZijK2rBk05aHtnTla+vhW1coXbswhFiSF2lxqVA3PW02O4797IgOc+7vAG
HTthr2RZq8SNxLAZ8wS9xKN7cZP1EUllKYHU1CDgeQqZOLiqIjQilDF25aWrBH4wUCoIQGOIBFV5
WpwUox6dybioKj+iDQ/KP9NlTlMBkJLSGbYoeik+s01rDzdWXRbK6Ryz7+o8vy1EUEXhHLAdotxE
VLVDs+tDt6D+ak9q1cK2z7R79Li+fQ3Fh6iAsHG3xlVzGJD8VYXKIhkD1c6y8EoW5ToB85dtvjdZ
3X7yDe1DC02RmQ7bxw6NyzaM/ZzR0ZvDV4NSKoIoLoc4DVVxNpimKbWCtg2X3v9SPvsE+DBGk7Hb
hgvEtplVhqwxzQgomT3cK922L8EZTcgzpN6UgDjyAGjXwIpa2/ARFyTQJr3vJsuyQgeI2NaSI44p
Hf6DYVH0YnI7Viq1BxNi0ZX2VryCq3gNN8MKkkXx8HJ5k4c4zvP2zSDWD6Z2ZwOxxvoA41cRYb50
ddy+bLyXBIFd/uHt7KLQmkelM6j3CeON2ywPZ6qjrKR6fqJIeOwhlk/W+PIQ8tPkWIT+BFsMII/6
/XDOzf/bTwRD72RY2ID2Jcz+O7EeLYtcHhgaSnHhvWvPnryn22Dqn68zThHGe35NDXQaapsa3WmL
iw4WAxq0X265CemBH2d+Cs3SD/RHefRqXdFbO+JBfk0PjR3yJ/C2uUC/VSSzhfEMnClj1UVdOt2T
x1UA7sSQqNW+uzAg5nM8tNJ9AviNajO7zIcxYoKlRg1/ZQFG4/aqy1Ji2w3RcLqVVnn5B1Xv0aVm
6or7+9W01Qa640zzGQXJ8hVqzU965EeUaCne0Z70lxd9ScrttfILxaIXuaUdTUoAT8xngwa/E55J
5CVz+7yuSifH4HOr0kG8/GvbFzysUNBU+LB00CZVh+UB014YUiVlxLT6AZfgv7KuGy7eoakIC03M
3trcbdN/7QFYkWVFmOmCLw/QodBb70uWPmIPhstth4eMM1nTw6P4CcbLGQrrG/uxcmM8TLvZh3MB
KTBLiz52UeT4e6TIteFsBYpy/iru+9D45rISHqJ7LC7XjbsZg8Eb4fkhpHSyB46NtXzxiiR3mVId
or7LcnbMiYRqnS5t3/tJukpAD7IFN+46+GkCC6Z88Kzv0qG9uPzKj4DsCzCypWnp/wRzRpJ7ldOB
nzj8nt+l2mHhn4fz8NbWoQP8UC9foMTo/a2pjBDqeSE6luIqJzseHrhTX7b/yOELa2oJQKg0inSF
qoG0YemBqbiRffcErgHqtE80n/nP5DU3X7djsPJOgyR2chjnjQWL7+fB7QqUblsMWW/w3XgMFmDz
MiJpCwCdWaD3X5UFMG5G+w6pIsbgzrAp0Edt7t/9+K5TVES6OTvSr6sD1lffDZig+rG81NYioCkO
z3YNiA8AJ3IOBKb9POY7zXGtgK272E/7yLL8v7zWikgDf3Cu1ADiy6oclfSx6jwOEBg9+8K0ZLu+
jZdwF9cx6N0cZkPUNTZhfFboFhuj7Z/iH4b+KXUU4Tn88vXBiIH24UWxbiraeYYoYPrnTNCo9tbz
knoYm72Jti3nQpeSc2kDifuyef9/4JbMMV2gTTkNBFRh4CEpTumwBuUghQZhnqY+Uqnw/nZotsm7
RJ2jBJ1xLsxfgmUyAHWAetu0sWgbWB72hJxWdbMW5TrvQEXBJ1nkUXd+THXBvH/LeuGF5UJsgNt6
RGBbRlKQEiJE1IQECxRsyN6Kdvhe620Zw7JQloh1PQg0on0jGoZsLNOLzZRQXnYbHpwauUV0Tk0K
1gM0LxDUGgWtomYsf6TIkf1kkoTgIzFynv53prWHFip4oIcYoaAFaa5CVW5MlAobPnB7UuC5mXrY
0Jd5WMGbYcX4no9BG4qjpKYRxSY+LVL4AuBHX0qul9Qu5tEsp9M8TrE4dlT0RBbgbyFN8YbDwlwU
ficQ6i4cRm0KsK1wVcslOXHG7FiA31MrBas6pJjLFVKXreYRxRED6IOhjRBfZ7fPIQ1zX1/+P/OM
j1a9hNvTU+qqS0u3DW9sWGVx2z1wlrynKKac5xqUyFEAYJpK8mQw4ZUqu2VRaRmdvzu7RwofZhsp
MXD5G1mElwptdfx0p+K9kWebvPK042RvZr/NYyRlpbAMGWIs6Q8VhGY/fshv03ORKCppBTuSl2QG
czsdUXuwi5UyMjzlrpxoKuSZbdUV3YqTadte2WXyCPnYPdm7AHCpWyKNyvILpeoYQtRdVmHjqV/o
SUiejZSIazujERUSH1VBY2o3slzeNHhhFmSMFhekO7h0AOBygfM90koGmuRThgxtjl4rJ0hovhTc
VU6eo8/zgeo12DR8N396Cd/lamU2qg0ERg0tQ+qohmMAWrsMQwqCsILwm/Qs5+ch0l9nPZ90n3lx
WHxL4q6Oh3ZU++00FWc/aRcpPqlAzs2f3EKl3uYJaKCNKfRPmCe6sM9zaVDKOSzyD/DPpcJeLtED
yDUEXH4ELRei1cIxxKzYY2N/NFVf93Kn/yPGP96Foqd2ys1zjJ8hXDacYp0XIGt2slisxDlX5EUN
wlJbEfjerO2KTwI64f6rTo3TBt6uiN+iVapjFIg+/GDroU+vflHdHkdkiE3J0tfx29M+ihek2Ous
wX5zwFxRBFxjCepDtgDtMAxvdZlxCHFWbY4hAfINhbWcmz59N3z6oBZq2z6v9O4ApXPqKYE7w6aX
3R1w5nLo52mFtclp1uidiuq3tptg080/njIioqnm0yLe4sPm44ZutRkae2PigToNnrU9IP0pHYCc
GByhrb6FIgLHTbQftpWJGYUMadPQbKijkUfYPDm9Z7vm8rDiu49eMYYoHUvjkFEt8Wek0XXtSUyS
/XzFZV0vHRQW+G7PbDvZi/DnLIKAZAfjg/FPPR2R04P4uRzs6I5mC0T2C4HzP+hRcD3b1Vfa7MPW
GNnKbm3F4q0S407b0EqUuX3jAvV4zXz2yheEnYOTZnfdV/l6kpyVbAdxG/Eup8mvuG/BisjL0tKF
KmEIXj2eQJN6Vt20noz78E8o4oh8dJVknxodHmzL9Zj24Uyjrh36qR53UCFgYTYhrnQhuavLCmJ6
AfKHqqQNbpZv8JPAJ1hcSWV2GDIPjOusKkKo+4+ynJdjJsOT6p29YRWRx/ZolJLP4cLwVrig8VHl
Sefb0ImoOAjBHcRp03UxQ9g7dK610aNut+DpPG9pObMkIrh7G+mpHvnl/viTZRGa+3Rzk+PbNqGq
fIy1ZQi4MAyHZSnFYex5sm2cANtrpAJuQsNGalUitHtCfqm/p6Ff6jSqwpymoXtGAp1Jsbg4p+gn
MssIT5BZSXjRhrsCuiLK8EdorI4jZ9lEVUXwcsBewq/9FScULUFVIL4UHajuVakUFvh5agON+cOr
h4m3W+95YD4gcGrrN8jSKVxTH2LOzd1gVzHs0Hd1qol7xyBtQtp7q5SyAultHQ3174/OlXmN/zzA
zKm+tCvJySeoelChl3bKEOvfANOS0vBFOmmEUt27Ddwpy302mGC8GCTTywhrYo5yM7vPgsSHm8kc
u739rM68fUAy7ci/uff3/xnbBgOzvybIkaLEn6XH7txuRJa2o91ruwFK04QNStcf7ZBJPiuFaUMy
EZClEauzgyjSrzLfFKT/Ujc2wXo25AEdhSRDCZEYyWt12xDuYKBBIPyyJ8iDmXB4jlf6LunmppIX
l3H0xci5QDgQ5LnrsUQiy2jQhwoM03hQXISL3QIEPUozx+VHGZp4lTX54cbQtRYyBHqIU8/CuBoO
Ws69qdq/GMPzdBkwKYVat64IJrgbXZ83+MZacyNN9onWkrW2eYSby3wTyuoQEJfPrD1nDFfwOLhI
e8dSLZECQ5DVDjwgO5/V3WnZb/g4o/+aQGJHBh5PynlRJyZbh5LRemCH03MpGjmQ7/BdUm+FZXiS
bc75NGao2viCa/auAgl2b9VynoA/0sp5Lr6Jm5iu+uI1KirbNsxAsjqtJeyniRT+IDLERlGbSrMC
9nsSVKs3Epsp5zJll/5ftiQkua22Ye4OGI85fOu176mjWcr/J7YCMw3/tdwASBXamfLQlN2nvrm6
Ad1XELNbRa7IZO5UWhEA3iL+YXdqQcLvrkqAoX3cC3/WslLbn4vObL1iK+v32zGXc6zFpF2VRobQ
9Lm3OkhXWLk42F+bfrLBl1FfoRYTbA+vWI5IuGpR6WHScfaLWzbjzecXfvmlp3FFbUGoCDw+ASPf
AO7214dMznlVe98RGRUGAirgsxR8s8YG2bitn9UnoUrjPRFSDborwla5ocVWyxug+2hPoxo4MQ9w
zG66INpS06D41TGR0i507ucCcmIt77DQh4xtswTdiw+d4qsdynov5GgD3riF7w/B9DoGyA0IcSOa
OoThqK+htDPTrwyzZdYXHoRmeDp4Vn0XgyLoWc9hc/ZNZsd+WPWwh7ewsCZGRqQDUjjA0skVI5qi
2SOdMj8LvIhfclIcL71oochpGqj/zFvmOu59aeyXeo72H4L08x3kU0XjM14bE1eqMELZjJ9tC+sU
mNFdIP4a7Jn67KVqwxR9zsr7KzQKlWxLs5XNRSiw/WzfKwDzNFDB2VDWfke+8G0lvvWyfU0oetEl
XUJW8bUqO3JhyafuSeMg0D8qj3Cu8aInzXzmU9xq2QQuT4sgMElbLF3NBXp8WqrXC7ODPC+UuTKh
ISU0vG1zEktV1ISYM770m5U1sXM/YA0R3NjGqa9gN5gtWAfHXPoWRudJmjws4AWmST8RuDyCFkBD
8NaTci0rt9NRkaCKzG2zpTiz6VjF3eI5vWMrjcLXjYn3aaOzhwjJmfugOzgDuSGuK4ac49XsoU7t
yJn3t0CRGup0WQPwHOsEkl8SeSQp1bmRUoEXc5Ei9iyXcw+3lzMBvhU5lkBZIPJ4EVJ40u02sM6z
JGnWvirzPFKXyX3AgxKtRLxnKVzyw/LL5SXnImzyFJx7d8we/JskwRdGzXBB7GmtDw4yEpvk1DQ5
xwnWM2bATRXnG0r953CTySdt7ljI3yzGdkZ5X9BjHO8voy3wdsa3SYksg2eQ2OkRo7B+zU4WLSOM
9Cxyc0ITwfHLHRfUjmJ43clgODJggq9w612Fax/oGrYZACdjvGffXi3nvAOl7BQ81lkHTI1lqoU/
B7ehC0j1WblTUfGBz8jGw3eMVHco4GpYw4Zhv62SvgpH396p74uQK/ey1UY/4CjoqqO7+HcRoylu
joBulE7EC1on2/zdbrtAymidsCmRmWyT0a8bM+iK4o9iEBMeA7wvwRkjTf9BkGDSx9ene05QtOG4
lYwECLOkgoJM5vUiyKdq8AkNjkaO+w2H9od6MGT9m1D/JV/9PAEh9wOGbkHcmcp72u/ygsecJZ7b
YYcTt89bQV6VeHSflTYb0xeo/ZAzYumDxL3PO0xRNSommj0QcvI266cfh2snkUyr7npkcN4zjEys
LpcKOL9Awb+lB39G0dUMtRUhGLwDkhFKC6c8B9beyi9oCjZZm7bJaGAInLL1etzxFgYbWaey/krf
vJZkeoe8mnwwMrsaRd79zUgpFi5HaXgeW4sO/n56BlhSU+z4iMVRVmg5tAa+GnoYk0NkLEVPDf2q
BgN3wCsU++xG2ZkqEmmLCnq92mAgrFKDyNnbIukAl0fQHeSucGSdmpHIGnJ0bPi6GXMHfI3QzMbL
Ru2s2cc73a/wm0Ur400gQ7QsRfzTJaLvRp/OUTBvFa5aZUVGhO5O04bACRZ6oeX8jOj1s4/P9l3j
t5EUpDPU6mJAzfLa59RsN2JOCo8VB1ubziMPLrD3gVCw1reCOIxDtyasJYjM36JktJHHZ2pd2wgr
91tTWgy8X7Pw6LNJzRgr8MeJrB6KziVs3sd/xZxVxgXnFOjVB4QU6b3+YsNJxNfWavYZR4AbGaEi
G80uFnMJQaQ9N+DTXZoINs5+XX76Xf5xpy8iz3lpxCrMrimFdsj9dtPStJO2AreK4owoq2SxQGhp
wKMpfuz+hqvZBKIt/cKdFIFBoonqRYWXWDV6lYKsrSdtAHk6PKnyfNSN9PEoSvv6X67jOxOP9Jqd
Kcc0wDL88tH5AhrL57ILrLK8N7Ksi+LUBKY50dMUrrCvRQzghrdzyJWKUrTcpYNW+XMkpeGyMEHD
Z3sqCsg49Sc5RMLkrO1o4tJKR59vEv88/vY9p3IDvz9EOtfxoXQnLFbJfPiSm7jJZsOfe1/aK3yE
8GE/tnNqj5kTcKfoccTAwJ7/CX2gaQKOBip59KObWdks0j13g7Hv4DiD/DDXj9iW0VQTwOBeIh3J
f6kztaaPiyhThEHHK6ySihUx2kcO8iSQozbMRwuP/DpL96b1k8+R5PSNHbFMoSUKNdlNWFvouXCh
PciHLaUW4DhHQUfiLlShvrvGVKB3Ap+jdROs5o8uClqbcguh2dE3Z7sRXLGnkjJXUHY5asWcObGa
NNMhMxb5BGLvoDMsx9fUv0aIttznS3q5qjDyDHjY0yHUAUR8PyCo1ywM51BL4G/4z22HJNG3VZvI
HXWpJ1xn5hqNimjzveIhUNIfRr05DXLU6rgVwPnsp27wFKwp6F9gJWYX2Du1o+sfXzfopdOJbOjo
4LhGsWx3sibJ3pAP0jfR3Ql3dLPyEKxXTmcjr6VxKQjdJwblzOx6RqUmP3qXJcDUoJkrUnQoFrN2
ILJ7CAFCTsKBeO4EVacFNCF0+vVK11haBikakxWXZT1LJL+pFs4PBRy2L0cneprxW7Uk2/4fFo+C
i5iOeUvQEPxRULI4L9qy34B5YeI09UlMOgoTpHgQoQKZklqsOgAtLblD/VdyI9x8JThs+NDc6Qb+
Gy5csfPwPhO+9uP9EYiYnEDXoFkNGzWlHtzQ+jDX1pC9vRTnLYM1e2yf19Stg3ODVD2eJW9mp7+/
IwcN+iaPGwPBagjBXZq/1ZuoyV5JlHBWWCYll06B5eleBgyQvn8slgGHyFCwF4n0XGtVHlffnbfY
sxq6yLktbta1gHhMkx3cJT3T5pbu9MZTmsp6vTAWKf1HKE7VacKTaCk5RwqBiC22r2QB2AAICO53
JCF19w6RIEuwa50P4jNURjM0ewym/uXJWQBoDg0Ugd1CxoRRZKmF9WXXmOTljgosv54IR/O8YhG8
vsOJP5Z6LYHNckFUMKfRRWHmkZ+TsODMSr8Ii81mTR1pneoe0LANnJanDW+kIgvPot7fZdfZqDRD
N8NUQC6btuGxRN02mRKmxNuLKnGaDEXn0v5L937jef3apJs95q5ELH+D3SxJDYMsrmFKXB9dZ5h1
1Dnsl40j3fnLkAZz91pLyxzGySYZiFc1ia/hda7La1adcn4AXkERTAa1MX/B6RKWmde9TbkBI2Q+
CAT9b9LPy524TCBaYq8+YZxdI3jcYd8MOKoXmRRs/1nfLnBT+65cJeOJonDcbbKNqFwb9zp+8nGp
KOiVgS3EBHkkWeDhFFrt8gSdl/lnBvp/q7dQF7uwzHPGTHTtXgxMTZrWd2K0sd/rpslwboFrpxVc
qdzd5m8aMxjeXVu3QNfaXCTCN957xoO9ngeR1lAE3DAQpsA8NdcDCWmLNYUmaWNLAtZ2RDB8c8bX
M7N8F7fdkeTF//LKjw+9KhiS4QWrplUsmi0lqayh2zgtK6YgashCyc0kUlNgnCvGEsrcgcwIZVbz
qSlCs5LrsMCoOD7a4OajFHAZR0Obqh9BKvA6B2zoKzi068clIMM23t18E7KIIspVQnqni2efbaO7
CJjKtS5AAhD2R9M5sGb2Cc3V9bi9I/FxIz2gBAUgg8oFSXnvjW0crcTNJ7L0Muzv+C60zX9QQr1B
Nh190BwTGTSkiAunrTPMGkKphrbUnHHSbBKCTav565z5zbES+jwFRNBLIWiPTrv9B8HPN8AtHB6r
b55OQeRX2FbzabF+HxrwPgXDPL9XylrC0pRbdsiRa9EHycv+Kx8N9n48we/1CkIP//dd0vS0um0h
k2oyrSwH05zr4fjrkMPg0QKNoF9LsfNzwJXu3X/oOPuhOjzacXzdxl/AZNZjFkZKEeHcUwmGX2m1
beiEx+aPgC1VtiT2HIZFXOV0/tp9x2+bP4KblfEhygzdn6x6npoKAQyIFG53r7bqpkJudy33XogL
jfj7XSw7dV4VDTLLc0qbI+Azg8R/UQSt19z2QudkRBZFcoPYh6pZ9OaJK8L2KpAB3ORtJipunay1
ymmWURO2wvdFhZ4szjoVLKHkvssd1j96DusuxnNVqzAc84mEKpfPouQQpfNo0mBTQAaEyUDBXtEB
ZtqxChDJEwFp8sc/bNoo5Enb8D6NULINnh0ZCdfO8gznBvj7e92IMW2mV9L5/iOTfYOWUnpQqBt+
GaXxR2e/fwRh2NngSTMwCAM1BvhF/cGJK7t0ZdPeE0FrcyrNQdCBIlWnbjEmKpWHJHAdPZP35e9S
rjLUA+jebU3CEm7BVG3P0lnSGtL6bFO5C6Cxhc8TZYQamxA2HY3uyfOQeLdnpRW5d7EpICtDeFre
EvECFDlkWgWnF0KRPmwXytKU57rw8PwX8ZcWRWaqJkQhJthN2KiMVcxmfkayt3reyxobqLzh02qp
1ucOCUtbpjmh4HBxGa2enc9zoimm4VhTw4IRXHaI8z1SO35H6WUh92/hiFc2AkKY3KazigOsf/Si
QRxEwCB5FvIq0UPbNkVVhvPJBVA2wC2Obgh+fLImzY3qLtI/7U5zDfvNn7RRFoa4O7NevT82ZHgh
ZIINHSIi3k3l5r6hSpcKkvnKSiuWqVd6CqvFriCH6FhJ1EKm/pm2XCMrktMQxrG1wdSZioyqxV9j
/TV4f1l1pr2xEOkiGRgFHAadOUtEvfVd5W198hpBwE7GUvKFAZ6rNv0F2jgq8Gko6Wk10S6xPUvQ
zQNBSUt7R16Ti4s9K6buekqJyRB2uL79uAgg0N97I9wnd8rnRzz4Pm+548UTrlgxGehAf2KawrEP
TQSJl8NHjY0UjQ7HfRPyLYIEGs8j0XRkaSbcp/eZsQQ1dV17Ly8O+tN7ZclkG64yGtI0TPlngA7N
HkWhnGVDV5eiZRWs/WcrQn1TxF4ztRfvtGGLgSSJiNdQHbZmFaIvVfOwWfClQcqL12tncszlEY4D
WB3AfeUdwvo48O51pO9T0OzkKnvPegA1CJ+b5ysKqoCeff2G3IGDNd64T4gkJ7Br7ms3Q49HgIGf
5Wb3svnLkZS42GzUovlKcEMzTDxMIvhO8XBmc4LGvwDACHdI+iPFMLHOM4FjCtAC5j2u5juGTOyR
keDXYcPkCZQ8Vrg1Q4IOEHV6B4ydUbK1lhiUWvk7RatSBs1DKFKWI0mIRlgjFlcKWamgvgcaQrsb
o0N5AXdtcNXMroNCvxQaW6C3hMl81BtAt/jUfhUaeWrhzI4lDRYEjG1ej2he2q08KVx4B8dUM2wd
iBV2fMyEhkYGIb4tCIYrvBto3mxu8CzzOS/fGVxaegNiIbe/JzaKIPxMreAgdFbhgPUYEC+F8CLw
UmRctu1Ftu4Q/Q7BQptWFfidNeqBjxPUF9oF1XFN/7GmwjTWjl2oiH+YaGfELhQJ75J3SIuVHCzl
QdtIoT4o46QzIfB/XntcAR1dX4FFCtygwBRPi9KFtdw9pCeyS1b8UQr/yJs53g5GTtbtPo6St6Ao
wCedZocAs41Hn2NH6UUSO4BDAkvxFGLOCLYi7Y1OHgj51VZRJPouMM83ILPG6ueuFQbLEdBizQzT
QUwovlpTgqJyhjgixlgjXTxfeIFH3P8S65bzuIXSytpMYeey+EDiJK+c2p4C/+wlL5fmmL0dwC8F
S+ZtNn8aTfdH1SDG7xB40TEJPB6R72SKgHbraAOMCoZHQ10aAvTmaRJRPgdP8I7KbIdoRrODotcG
7gx0eaS2KIxp8YfmU/msNucE3FScbzq+hedJzsKVtXeUslRfeOXo1gMLzrJx2bWeNYjLw14FLiPP
cUGlnulVsOMm75k6EwaxN5N1NIMSWG0oG1bgohPD1GHFV9xn2lTE3ljxFzfuZYSM8lLcLm33Ld2L
jB6balIgQ1qqc6bfJ5aGlsTsD0qSYJukErWttZ3cLowWHtm9W9arUTHiyj3/qm3aOdywRybxKTY8
MjuBYKS2wf50Xy1a0kZXLN7nVoXUK+wc8zkcJj4qbt4YwVUvA4ECNJCoG1NGZJ2VWZri9TvHRosg
ieLBw9AhhWI7UiEKsAX+mN2sBuxXHJQHD0HCoCpOcaqjbsupNS2ULLITGRI0MGtpBZlhW3X9xViX
hdFbuyk2JDYef7u/zeU0KIXKvZ/1D4lyovfCCXBD13Dis3eegzvOT0KAZZ7sNzpIWG4zgvZvpVn2
CMj9jmOSUUkfn3pg+zoVjSrAUnHc0JLwvZMcZiAv2AOAk7NoOLvBSjv5SXy4IuYiNzwnjb3UIEa9
jkZGcPdyOYjvu90o0VfcMJ51edoUO2wy6f2fwqsusZGKHrMpjhDwUH21q9AlEcxR84w0gY9f+lQS
PXf+IJidFbrDV89A03WRwvIgOWNXm51+X88rwYIjcRxWYsMeGniRXkrL5ZYi+kSojp5qniUd5O4s
GrDeg3JaFocD3abdeFZGue87mCVLm6rSGKgA5h+Qbn8BRXK3qep1dW3GEpmlBNWsQFWQaQsMsuXl
hW351aYRSkKV29bgybRmqDXbZ88VwCweHu2QM/HG31KZhs9MD30W4dIfimOeZ3oJeTgBTJCBMwfN
11MsqldD5TBj287+FMrToJZVZg/39zAW5/ACKIVa2tz97pplgxvAB19O9TOn1bTWOFJQZx/ZGMSk
fqUOcBkQIjZu9NtAuoVrbckL0nVwZ+MZhc5+/V1WITt941GQ+Cj1OUuAAdvvUo+04gZ98074ON6o
PrlmlpPORkbxtsliZcG19gRsJXvZH8Ugt2n6mSbGp9rm5EjyjclUkZNkiqzFibGJa8atTi0jirt1
S6bOuDFQQTE/9XyjPfNQeBDiut8wpdSB+myFpwaYgDUGoKMCzQqdYwG4MSgF14U73+RMhPWt2I6z
/n3BLe0kmy0X07juGgAo1iprSaCaTygJDfZJLoHoLDvSjSSu/aZvJ4AlWnALCXo67SE2p05veWU8
KJuR9gn2f2ibmXRSih2xQCwcLncLFsso/uVFELn84rit7tJWqV+Tt7J0PYUiY9NvAiBcihvXNjdD
xcyNW6dAse5PNxGP35CJ0gHSpgigeqOYjt3w6NqhjbAchmdIdS2aTO3kqpmWgRCG8QVWf/dY4T+m
xYtJE8LXfANdaENT6Od+niHtZDGzlTLRtbrLVaEknr+hffaE+0pL9FRIoq7N13ruPPnmFDxwzEDx
QLrUSWSnqsG7j0WEqcnPdHhcT5UH1a8VSj0qPiG6bgF/ILyuIPq4AKSxdWrlLgrX6s01gdA5m6Ur
x+ZHvK4+8MtHHVR+ACUl0Twg3GzXIa/KZJRhxEn0HY0Hfn5yvU2q+7S9zIIaPVk+r3/+7DDR9EaN
XYwgeWKdTWnmcbjfTAEfg/VHVHDGZZb5LWzbCSOykR8GaTCsdLpb6M2g5kvBev74lUKkkUKWAl7v
XZc+vGltVPZOYNjLb+tswl4AmdD+TMocdDXIpfKLLuUkcDilplkVAPSQ+GZwnkEkDyJDMV8c9QDl
Q8XsDR/U17hU4n+YVylGT2MwkuAN+bUFmPPFsZyuLiy3BCy2ln6DoZueiZI8YYy+kq1Gp+4QW0pz
QNBRh5/h1s+Fjo5//gSemvUv18xQas0KUaDdZ6nYet0X3eijtMotS1oM3ZunlY5CdXGifKIG012D
X8t6xv5yXlljhhNp1ZyqWlgKgMy1/hBiijqVhBHf8Aet1C+2fml1g7/CC2VSYrFRy9dsHNqwaiUc
Qk7u7+RFtyjSPMLl/C3/23iTrACaLxoNdMqsbooQgL2fVOHy9fYxl0Yvs0oSC+m2YQE9Y426k2gr
wjtX+u6tbkaSnMszPlvsrznV/hk2wGXvton7Pirh2dgyExkc84/Jye4opJQnI/KZ3Ulc/bvcUAHl
fvMMgFH3EAcOIRAZQrnkFBJM4/wytnA0ur9BXZYBrsyoqeFoka2mD6/MAcFRBffBl75wASC85Hfb
KXx19JKIy0sLrORrguVUVm3lq8eDXuBBBR1tq5lYc6H1lSlzAdTtuZsIKpfdWb/pwtad0KxiqQg6
YcpiDPy7zaY8r19/rhxUgOeWz4JtOuHzv0xkLIPUnovJgcaAcvcmSpIytX7Lq335cX64MRG3xkv3
pbcufGnawvCPbXJbhQ2Nz+vO65y/nBN8+yMQ4I47zXnRjBXHpvRnX4IIF0xzYZIrOTziVIi21yYM
y4x8Xkl/B1HJxXsvQBW0hReJT8BIJT3br23r1vwtnWFAOXyDhsIABYDBT9yO71KXilMoAyytHIdU
ncGkfn1+8IDQfXVwa91cckaIVUn1vyDOLVsgi8K7UNJyr/XLuvbPhY2A6krlC3qKJQtfHLZfwPyb
jcsT80WLBDWKrTm5LaO/NU+4trqB5AWBrbFP4KfJd7317wC7cO7g5RcBj9sH7bo1ChZ3yFjXXn8q
aSzWsZ529K+VnB7sgQoHF6wRihV5LXSTPSQTBVcZBj4ye3gurGSYoTCzH87uyg+IGebAGLm4Dtnu
DRzxUKXFV/EqREOW3Q62fDfMmE+8Fag6plHR5VGtPeuNULnn+tp48sT4sb/Z1XA/kVYa3TKgiGE3
D7NR7oLPnDuEzKVwAggl8BD6ObI3PwCxJ4hkHrpgJTEsW6j7dOBNeWHUs552twhio/otehpOQ7vT
UkPRpYuxGgYPUIMEExaLDI1Ssl4E+BOCzrgWJD7TUArD8DwuVESU24Bn9ZQb6o3k0RJrKC659cLS
/O/i7PsuNZ1mNqAcPaQRJ9Itvz4OhQkTkmFe3XeMBkQGL+xuwWfhRWqASI/4z6m/5m2R6MeDxMXo
90uqWQncNOUWXWSOGWnAs1l1SiPQy10QxKUc2RzCUwLuCXJsCjoXSXu9FNVbiaa+mY8x3RbV28bo
SGpo01xb2hJFyhTrvo8GXAqaV0KGX6HMDrxmIWZ+RX7mjQMYnstXHNnJnU/zoQFlHx0mSUf2i9sy
Q0TVI0RhvAYCagbF9RxK32011X1NCBoY6GFaHWn2FujwgwLMHH++Q8QhsEG7h8S1yurXMwNlhrOB
UE+oPyvxCfK+/t8Ra6kxLhrtjO1vxUz26QbIWNqX0r2whDvVFm11CFGCaBgSfmFZLlRUv/KvoFyM
ez3WFQuNlAtsKkz+N2ePCE5GrgjQ9KBlDvFo46Qj+HoPAvBWNpbfR+o/B9lSymsEdxT7UByfsWPI
uJGX37GKoWhfij7mEW5PAAFdxthprtGcNvKSIAsjwl7To+UsK391ziYup0yHGaJd2KQIhlZASbrd
8MvHx7OD2MSMw5qQBlnhGAQ/303ndtU7yBBJ/oBC3XH2uJseYDXiWeiNapTZEhY+5vgUahMp4ofi
dm8Af1mCjzKK8PGJEivspuFHjuaUvKrwsfwo39CLj/SfJtLaQYt4afkxYRFMeL+9BXfsKYzVAoIU
HCtmQnHWruu5J3FE5dqSfQedRed7/W//rL8pp+kM9WnkUiUY/fcDyVl01xmiPUEL2ow7WorgcBBi
Ua+NxubVnnB9LI6AwPYBh+EqyO8prObhr/KAoMn4vTYKbDq1iawGDext62m4Qs73+wx+rzv/icoK
e7R1JrE297DxJmoonPw+zfW/3xQF1kcVkurGKdXK/upRVLQaLVutcvnaTfoGVlbXKHOuVpWiXKMo
GqhQJ50HTRTauA+0QGThy68IGa1kZhIiDiPPtimBiWjeiqjC05adtQIzC2q9aAisLfX1gxOZJvDn
DZQ+d3rWjqqScyOVszD5+HTo9fHuEH1hcZjEu10IPqa6mAslyXrGGQyGy0tgoDyHZmLY0VKBuPGr
di+vo0z8CNk+jbPQNn3zxOMycIFuEjySu2l3liLT2ScqEPsD9pZMkatxzK2ZaUX5Oj7nguKXF3Fv
1chOHz+BHNZAcxi8I0+QU7yuR2RLGt1D5ObuV0a3MwOsjGSLhyp/3iEcSVNWTRJLkbWre1nmXxFJ
2vRpkMyggyVCV8KmOvz/rXMbDW0kZJFhvIEBLkz+w1aJvkm/WdscJA6iBztvALtvD/k5dXFDhKFn
YWicGcDZffI7/UaPydcW2lkOqVxq4R9DD3OlNbMr8nLMKN9TnwiBOmN7rUyAfrsRypPdguW2Hc0J
eFsCYMKLgTLhVqS1aewgu5CQgxwS73ji6YFMh+SAiDo0SIY4ChtTJ94H4OQloV3kQWKTv+XrWo+a
KOFih7VqmSMEpuv0w+uuAnfye0bMAXHBaWcOcYXxcjJoHJtpabLhASOFvwXufBWKDzuq2AJ1LrW+
RlTwODZ1rMjwYMXplCTRyLZha8bIQhqJ3PGY+/Px8dE5xuTMnXZWxNETR9wGx445DjQDVo8HDVWq
FoU13w1WOijZrowi9qgK887MrpPIi6tIcdm3peuFKAGfLRmYjryCYAOP2NxFFFYfBByPg+2oxRQU
vAw/g+HLsutjhiLXdJIzEcVq/ePljbVCx+TnoP/1XyKM3eb7p6yCwrNcNVbaV7mcgw//AndhS8wo
Ms8b+r98R/dNYXsg4DDzBvdTkz7WPybIU14FeeDxITYZffcNMug2aNkndvGIMo7NOKy9TulbJ0e7
aeUei0pR9K7HoCda04iDLC4yPQc1ROn01szUyOEB0DqBulmkMjo8uORj3Rz8ONGo26eAKpZilOL7
w8F8KleZRtx+WRredpmjIkjj721iqZCwynWmlxn9gqtWGu3hk2unGXeXbLxgcOVR8JRPv8lmbfxe
iDrDkfnxk/7meZoeAymRCkKPsP7ar7yyKlDmNrSH/Pjd3uHnGD1gTPy5CFoj7t4CiJG/8ZLNxwQP
Xyy2TVdiSvZ71Hg3KFavRapLphVjOpzvwMZxtq4Rc/2JNUuHEndR2RolX4lRJ2mQOhI+2+CUs2S3
vfw8QYJA8HGEy+cp+a1z2K6LEDmLqyEe5L591oKiKVh6mJA2X+QOVVVJ6s7clb05cpMbzMOS6Vs/
2Tup1HtNXJ6BbNXahqALfhEB8aS7byh4wzhbOoemfu4lMWLVLW2SdHdN9Y0UUYJt0EdafWm7KcuB
JjXuW4Ap2/gIqHwJ5+y04UCJxLNxKH1JGvWbds1sHqFoVkaG3rWHiuTrJJZjVzYCeRyUt43589am
apXokMhaB0mwc6yvrZxLleMCJglYEUrtCDurOR5e2mcRBjSxCrqLyhG/1GJndSTWYopMVBgDv/g7
1CAYcdOChBnGMG25u4s2YSaLzY4S6xGz26XPX2i9hhLTc3GLDvp8+REuoyK98t8OWh6PV9WW1y+b
No3C9aF+PePlACONfaLlCNbLl4PpRLZAPtFe3mRQGweZqqt/vhjFf/awMy1RGclH2SLy1FGl3rDc
TAF72Hc+Lmzs0fi5X1YHc7aImLkCUC+k/ZYhIPjkDznIiuZinkOCeuSYAY87GbK/9bFNbzcYYJmz
RMNY94RGNicRadH0LnGtRZkgFyCaaymbQC+g0GiXKDlFI9vrJ4uyfp5cOEAtF38130XH5Sx51m/f
5bkfuwgkjigQyqnlqV3JSKL0S1jF4WRIFehO0fwnYRFFOojkwLM8hC7kOktSehHnFVapnVoFn8IB
nq4aIlpu5ZGogZcmwIJtGnIx1XvZ/tfDAlSnQ89RUnFMK1LeU/yYLiv4B4kJEOnOZh+JL6Gqf0oD
afmnU+OmCuCiJJQnf/y5DvtLa6NDVlY2pLJtFAuOH9KlZHBEvJcegypwWznTTly4p4QRK4cDMl7S
LeYnmHgPjFOxXYnW9fZg8n1gDVYhZ2/UrKdg8v2gee0LbP3Aomx9TGLNRrru0LLIcG128yADck+e
6qZXt4tUVaZ1XBrYOEUYI74ujZHXVBB+eM3R0QmnCuaZNYkddHiWHX9bLWqGVZH8S2DfKkxsk92w
zYBJZN1YQ/8o0tr9AbdEuBdkhAbQ5opsB0Ns/dLp8OJVfsXttM5S7Ug11nPLGRYvv3V1t505uipy
PHXRhQIvi8vaF9Xl84gOR6uoVhEq10fNlWh4W4Rfb7ilPfDrLVay9ryPYp9Wh51kyEDFBgpa4pqN
FFEt1M8NgLUxqSAO8v2JMJp0gfTRPfggiq5scj0qtmAvGHhdGJz/d/55U/yzlf7mVCahnotiYN16
aK4wmCtej0XnNjXqGjttlTowFaMT6uBy5ldRHcHyPcPMHE2uCcPDKi9vQIrThWEv8SNdehJk9n/O
sLb/8lweJ8lqx7O3TrKqpGt5SGwkCN5e7K7QAbo0JN/9Nmd2oltlRvr7EmYAkaCJaxZy160DSUPb
WqjhfNyQ35E6cOmjtBNez6r+mSYo1oKCqMdnSWPPVwtTt9nrH53FQPDgcAEz/XMUsWf5eTcbBI+f
NyZPYF0/t9aHjGDpkx/msFYBZIS7mAlOKvpSv4bgQzdwMnXkLUJOvHD6bFfHfZXLM2eq1MH5d4SV
XudNIj2hKa9Ieh0PoV6ZCFY8YKXksUtW+6IophLUlBPnquT0Zm5+YMyxWLkUy0DB0ibGLpdHyLsJ
lJavyHFccSFinuzZD/kIUWZ2Ytv+j9Run34BIj3AWSGT5QvbRoM8T7ZtBI3PCkwdJrBjNfu1X9vs
qQq2O3Zz4lbr2OW2jJN8zdfi5dXqzG++2M8SBR+0v2zn8KA2G8rgvFo3OSUqtOIhYT0qMTvjjb/m
scRb20hiowGUHxr9oFPsfnkLO2iUe7xL1YElS5E0mB0ZQaIsEUNX+BxoKtV4907A57pUcVkRR7/a
QwNK5+1jZte1ZZEi06QILqdhWwJgcajLE02glno3ALs6aosSVHsExvkyTmGbIV1dgVCZXEld0rxp
6QbdragY1s4ZyPPJHmkmKYWvLgLn7f9lF2/yT5R7vurN9frBTqQ4LGBNFNXXpWAS96KoJ7o43Wb5
dqyxAwaLlNzHOxxd+wm69GfbVYXQVsx5RLYNd0TQ6d4jAWUmq9UiFTtM/2wzscMFwPBmxBIhywJY
qd4VccP5E8FVp70cUUTjTuRQPOJbW/x2G8zzXkzSCAiNHVv/dvzOP6gqP7yGK0QgnJvTuM1tzF+W
Agg7gxTSaMxA2x9AX5SS38/IlSABLmSZjNmvFkl8ACu7qe01JEufU88/XyBf/vAzYm9Y7ZyTGCF0
9OusibPBzQBG1xaNdUVXrrsWCkprTYcIER7I5tIqN589YWn7FC67LZGAlNzaR5CKoOyiFIkAbTTw
U32tKRx2EhHuxdVltkRGKzV4bOzXgZ4FXH8mKxG4GiRqo5ZeWohCgsZFzJFVEwnau6NAwkgz4vX4
TcpoeSCK5YrYpiQp+Mais2hjbcxP29r7IKvRaAsJo19f/rj1Ed1lW9sWDpk03B3VuGwN2HT0z1HG
BDsbtqpnTbKobmyjBPqz06OjI5D51+EQr81QtdBnTcwC/afNp2W9MNGPEcZrVdgP6vQl9pkKOtDs
xWhguLjFwz2xqJEW/b5W2YBqimneuHp2OHxeurISSIUP0JUNCtLbkL0ik46vrvk6d77riOEVrCYE
Q7zAbrcvbQZDD0k1S0+dgo2o0qRajSryGs2ZAYt7k6PJwra9eS0q1YW4RVI3RUv4z6Sm99DlFEvO
cdHZU//D3efmZgYLlwpVDDe8wy9dI3+p9ChvY/UvSm9S+Ad1H5eW3vb8aqACjLB99gv0SWx4DfFb
3ZofIdxds6N53AF8xRBr2OLUI/R4XAA+wLwlDhY3paBabkaW/jg0OFuMWU9OXD4wyyM2M6ZAP496
STjBCUdyhtK9/qpUADbaHaaWXMT2wOAektRf6lb2Qs2lnmnUY++J/d0H+HwvXeGZ4FXuLUxkkFmI
QXrQEgt21MLv1YHawjI7XHgkQeDRy2X3BJ4FTTo2iN9Qk4AnUDVuB7iKcW0+Kr3kTtcGwaMtFwMe
fbKlDMDELruLwZ+C6DNI8kutb5G+1igNQ9pRnOrnCsaMSfRh07xtCr0XDHO+eUfsrpJiZGWo7UFx
jfe75QdrqyI/YXr497G7afL+IRDzxP265hgSnnOmWgk3vjUGrgfe19lJYbHkrzpHcodKZhBOVS2t
j4+hj8XpfelqNgkbeFKGfdy6JP/ifVq0F7MVopyqpyDP9fgRLmJ3kKThGkoWVkLUjSwz87OK/WKs
t09+A8sAiGtxdrNVUmL2K47n+b51ig6kC0hFQ+slGQ+2nnMKulhz27acOkP5Ulfvvsc4C3i6M5YS
kHwNCWTqcBV2Y+luad3E/1WK1d/JWf9vKgTtU5cv22QJd+5e1VUqKrlJdyqI9L8zp+JqamN1qKtR
y68pI3Gjlb0/JAPcwTaq4Z/E+w586bfGNQ9BSx0edf2wpYMxmKXB++1TOX/3ZyE+uJ7R4uhZLjua
HuvEbB3HQJJ2Qo5HNTRFhh3ZGlNymGQ1IZ9PS61q/rF5yHRU/JmMATwQqjx3CKcLII2zwUulsdRy
gQjU/dFpwyUv8xz6nvno9UgBdXib27GxvbwsP+eXHDk6NfY/zcB9arMbkaBcmkKm6q2n61fNdnZq
YXjIIFYMEDnPSX/CaRBz68oddpxn52QvwK+VlFKxlWBK1iZQ4lwK+rjg8pjFwB1lxOJVZ92BixQW
lWc16iFmbZ01Gk8zwhusUNyhXY3nf/iulIne5yYTl7Q6WJCs68TTHIwD3Gbx/li4tjB1qUr/dXfE
bkYapVk18TZaRtWYg100SbNiEMhFnAeWQzWsQtVHfvNrpdsw7TBMZsx/K03+4sYdz7lWSkwf9KLB
5adIX0fPBpOR5NNtfeoYAwMHIgg591cRCusBGbEkt6QmJTLXty2hUijZ1wZtvO+uOjPWFLdR0VJs
fVmf4I4AUgS7Qyi8PCUutqZRDcOqNRTRae3VwneyvKsf9VYWm9PJllsQ0T1hmdERzbs2/erYw4Zt
enwcjP7Ae7HZe3u9fSRNCNPOdXY9k6t12V/Fmt7DUScmfT7iWhyBDby8Dwf/t7fFNra15U08Limk
gBh18+Vfk/aFV0z31JttvebZbarKqpxstDR8wZI5K0YBGcatVMV6tKYheSzs9Zb/woChhQEIcYd/
lU+neDMuOez6QrSulz+oE0XoA56MeB7RSHakbcqF8kRIBbPS/tP7MMyG6vJz5+LWvbYK7RB436gE
3g8uN2Bski4ZgM34K7V+/Ivpraoy7q59j//af8IpN73Vc3m9qW1PvpKSsJ15kALkSaLEy4iquZEu
n9DYWNQHNBLeYTDv3CqWHC2wcSKPJZ0Qpo1H8P21pSgVR0M5mmY45t5wqyGdYCSca4S/tLlt+I3C
Mcc5qNLFs1NdBsG0ITcwg7LEKE8edKNxEJPXjOZeVpq3MOIbr2m2o1o4ZqnXcY4i8Iv5pa4Xn2XA
2OQEjBSmn0feFLbD/7GwHSry8yYoIkRAv/zPe4ot477gyzYKZ8Dpu/w+kPf/AlTjICC7PbtwwTFw
fbNSreRFlT0d8X7lRypIeSMzE8hTe72aYuppAr3R0BUx87PRuleG1WUe2M72bxeNdlDDREOqxqaw
vZvEZ1blt7N7Zg38pGCtkaK59bhaq6YHIBK5uqL4TXjXq9+q4RnZsjTdSPeIaTrMjc56qraWlScE
mW/uatZYBkD3JrnwzO4BhxhcP+6CiEtznckJ2KqaPW/OWf88kISLMTusmV7qTTH+ZT6nyBnDdklj
GdEE7wdW5mAw9qKTE5EsdB6efJsicsNDSpkGmqgmyA7TzWAlzMvMJBcRCuxi2qiMcjsuRqR/eXfn
Hs+KkvvZGcd2vXjRxGEkNDH0NG6+GFsUIIuIqn/MYyXPolkQKP116AdImz5qDqtmVqxD/RdIIwya
sC90uw3HpLSIjoAe07XTLBhuJNb+AGyhsJQOV8ntx5TZY5zjitf0YbXVSrmPuSYQNg1s0MUgUVaR
pNf5JDrJqmRg+tCthTswrKymK98tJF8lzfX0FeylvCsm1nOyPEphG3edjZf0RO9o2uyu6sMQhu8y
zOTI1PJLYzyJAjZ36mPuxr0DIPFhvAK/TZr64Ln8uV5qi31ltU9MZKd06dtrslh98RT5K/FKdJ/+
T8YWn4xPJye9v+sYpjpKfxr90TgqAufV5LOuwROjMuQ7NRwn8oVtqPT+BnnbijF/neZhD/8HbICC
iNJGMw6sTikYdTEdJ4OsY+wCU2+IIOuxeJBc3gY7xLzaGH1qpsARxw2qNg/zDtXPxO/7SF9Y48TP
XLTK9Y7yjjCLTqBQxkvHyzCkBujlgMZ+UEf2Zy8rrnukjQmiLk+NucuhsmC93S9J/eoAjtIR64Th
DUWiXCFfDwKDy3ER95Ee4NNdDAYZNQSE/DnHjgEAEfvj+8p5opV/ATEsDMYRxwTNx1bwv6wg4v31
2uB263yBnel+CK9yb/4/dO29IGdUATR/rgZI3I60dFM+H4IGdp3LmNH6JQ32gp8KCcbrUuML2Tye
lbIfCWkwtXujs+ORx2ttQZBK0e5W31uWJ0mXGrQ+53Beb4uBZucaGlo5C2ctp6ZsOCDSnKNQ2ubP
0HBh18Lx/ni/RTkJuvth/MhJnvnnJPamD+NWLXXXj0rG9tud3FXXoQNdixlNb5HHpXDZQ0jKUrQ3
uRZMRAEbOZ/pR+/muonhud4l72+bTeEV8YSIZmTx892VuafjBlSh3qp1HbnHU+LIEO9Uiq0X5mlv
qmzugAe53S/sLU98mkCyPc5nUdaqirx1xJVFtyat1iayONJZG5P0nYOKvV+2RRrYPf4PZen1Zn9V
0+JYuo4cDSTXxV2BTFtG4UOWlIEtDtGNAeNbMg7DrZ4u+qNc830B0RUQnkNVLEr7UMMQZLG8qPDc
wfcYcBr5BlDkMCo3ClQmohfddqo6UHdJS3XNrfUZWDesMuZaYfDahVwAL4XyiZu+JqxV/XAZ1w5Z
jVEbI+mPcTNdtXSdzTNI+q4I0P+NZS67LQmh8/2MkwTvumQzUQlt/uBSFXrX/qKeCAphcQHOfY5m
JYakqxd6Y8dTsPjqYPOVLFHCesmm7Mj/JfSw4m10u0E0Qk9MFie2TLEO3kmO5EQG7FsPyNfikvgP
DpSBwsGbA12K5VPljKAyNz3KudS9ZrQraag3LG7Y5RusVY+yuBizAkeqOK353PXLwXZ0IWpgVU2n
7hbUMw7Z5lwjAKMCGO8gxJefxz+SkkPUdUnWyeXquBdMu2Mqll7v2ekPirxYhFWJFPGKFl/1RJCT
ANQukNYtNcKm0iwhDOL1fjqpEnaCGheIumbA96+oUkljggnb9Z9TcgMx3TETuWWFBKbGHdyPL2hQ
lMdkcniHQ++lgxFXhdjt7GrtDc9AvqzYcVLMCC1+bFJSp8NuronmkXvvtrlCVenqXewnJE+D1YnV
pOD7WDFEzC2gLpwLdM3jN5qgWLdRgsnZyjw1i+/BfWjEW5GRpUd8aIEPMLHudtLuxgmUesqWcQEZ
S8a3Op7r/OG3CLeD2GjdWX/Z/cz+ltrXYFXrFhCfHXMA4GQLShChMJfhTbpYqHZEWi16/JxOJ2RN
WGVgJ7EKM0td3MCyD/LmY0AbcmHMxfdirMWOJPCGQFvtm0A9YDgfyOqZHSrCSyYHXzeEQJlBVDG8
x5vuOo57rHry8TYzGXpzg0D0G9roRFIGQWQrXi7NReoF/EVvwEYCXfv79coyMySDWKdJ7DiLhrwS
VKGgzLk+9LA+3RDscaILp5RkMWyap6gIF46pBPrzbwDgs2NAXl/jnHeLm18NG7jarAHOCdo+uXYq
O3h5dhlLwJH+AdG3TSuqDukTXDOQu0xgtN8W75xIfz2QL0kiqznC+pG3JNDfcbunff4cqfSI7UUH
jaxxqGeb4eANG+MyXYBUmSVxIjX0ogvu+dD8mMuCwMAHROLu9D5Irdp6hZKcIgATxKLm0hFWvGwv
F+L1nnfE+2mNjLsUY8G16vxjrG3CLPPuQYMqIvEYJKqFssQE/J1BmDoMfS3+SkqPp7yCDSrvC3l8
H+WoW+JL2BdQ3yqHOLa8ZZNgDhd68px+QvaBMj6B8Ox6JS+MkEDDI401kM3rPj/RqxEuFvgkcp3W
NBXcpofGA3zmnXytrxrLwbq/8qkZy1LP7wP5OtnPYp3rusoISqeHfvUl40/elKMKCOWywEMFzjqL
qNdwUSOCmJ5+wanZlZgWRJAqKO12HgV38QV4qJtlS8T/bFNumbNaw/LHqnK0eaypPSs/VCo5LmJP
CgymsnBw1F+yOozfFx6thC2YDQlFegG67MLdrQqMag7vlwqY9fMaNCdqfbD+CBv3bFDYnbLApbRP
FsAtMYp26PYHt6IbMyU3ROC9iyRZMdFwgCYFoc7/0MSC5ylIJdjumJf55aBv5DL8MwHtfzggxYcM
VfK7Vzf8ojbrWjrNuXh7cGNKeayvDuN2GRxZ5dQ6l2C5QvinfOzg6AzJUqtyBJjXI+zvcnOioQhx
ScGF+AV6so31iLpwB95Td6X+55ECV86j4Zbtz0DIZrF0LCpKMMpsLhFTqv7d3QHff/HwE1JQonTy
Ps4ycTLp2JD1VH3Akn6AxS44eruolfuvqBvGD1JylG8QaWaejme7GgeV30LNTxH6oqFq6eR32nrR
CzCfSc1vz3w3z660qT48gWeTq3Tm3pXZdmufgb7F6KFZgEcF99fxiYppaOjua05UfKy+uP5xWxjn
QtnzORBsV2FWyQLxvh48T596WiTLq7k1uk7HWlm+99jmoyu5EV3hiPfXS3tbaRUZy6ekJjdfcR4k
FgybCTdOd5CMsjDeL1hztyIc1tcDSJVWznPJY4hQK6UJF6+QTCRUNEBRx+TFMD4U1VbNonbqtigQ
qYqYFcfMbluvpMjenTjokoI9fzgqaDR/8xGyvUPBzZSuGeMDvkTI+9u4Qire3Q0ibu5QxmNrU9sb
Tnd2Dpg82gjoXmgKqEh7ccYFHv09O1+ydZcPJOcTjBvHlwMQKoIlKBZYo6vMrcFcfOPyWmERmdhm
1STU8cL0D9eaabSmVY+VTSfnEIXp6pLp8RKASAlMlkRNYroCQ0cPFecg4Yygg+XVJ5qQBc7gLXtX
ATnHRiZGRIcwnmB1CO3sqgxMhiTFtsjsctvhbGy9WMMAimqCyK55jjN2/loD85B9roT590js9e01
UQGfiNzrxv4YH4/uXGqKhNQ3WgOP1P5ynQTDWeIzoSjOOEyTBNEbE0z8s8pTkmjao7JtsqNDXzoY
HJnpHg9Itt0oRxPP5rBdd0tWg76+2ZKs8uTeTHZ/PqwnjRVapP/ERSMUvd/RNxFTubepYWg0dr8t
D9AuQ4BOha47konW27LUT+0ZJEbLokSsERoJyGwCJUE4DQgT5quLVReZb8x9c2hGBgmrVCpAIBTt
I7XdNxbry6Tudbbr4yyFjFQfQlWUVNPJ3H0r//m1vQmRYl5fJvzKX0OaXeHyNBc585+j5CSwFOV/
Tw2xqVx6T7VBA8BjP4Y2h2XpkGWJSIB664OfBdAXGArutOXgcelFpBA1bn5zuADfXHyjKjZFlErg
fUHxe99sQyaYKcyJ64eiNeggP8b9MDPnLenZX2n8TFv3937iwUQcUwCg068sOARAOTYzTrxaQoZn
311o7RmWxJ+EKMX33Nj1N58zy3fJqq0zlqLHlb74dGtIHo1/Ij0H0Rf6tVLdWrWydNmIbNbUZmMX
BocWT7EwRWALWq6jBVLtAv6MHDwjEJ1YJ5GhhslNKlrCwvVwdJhqnWOHUeiPSYk3bZripQxcThg3
fu79/FUwyzzMhVNAtZqAdRJ16syrPvUv4Q/WundLc7HV4zhlWujeDbAy60XaummODXMLvFj4lkJ4
yEwy0yS9Zo3ssptDg94YZOAUfo1QNPVYGJT5xSbRZWCh2gSk9jtav8431IXfposZLzkQMCFJ5jeO
fYpquDZ9SQPVpbV1vcOx9lcJn02rA2Y+s2jClmmUdBUT9mU7sxW1BEraYpu5A8dDMGdExrb44/eZ
iPYSR21YjQMl7Z1l2cT66g+YNinncSeinNdH8xxJffcGHnn/JeJMHoMtFG+XrcjL12hbjGWKur3i
juv3HPOb7JXhctHN09f0+1h+QjW4nN99qxQ/mQ7QH/00FPiBXeOjW7tr64+vwMu9guB5Vp1tYg09
+Lcn8TMYDAeI7/GgSojtwLRKSfV6uATvZ89WjU76nmdwf13SRZLR+BhdDkP9kbgkd0D12qizAl+w
ChmufATOUjknEAICvU7SQR4KPhYHNFHjwlixmLq3tiVt4ya72dGBnJrqr9uVRGts4UspSHobFJOm
91a+zdjYNDTvW8W/g302X4XKMaliX8zHZtmf20EygCsrcx+LWs9qPKxYD+q4yyBtbMpJPz66VEBI
FMfK14dfSgo3aGI2TQM64/GfNl/s0S4jEJY+by62G/q/TSJsa4AkErr2qPhD0twIImYJUY2o44pM
ao55rJOAGVl68RrVkOcOc99DeDI8aVDk1FCirqARjCwUJ45xpbcqtgxDMRgKpAdzmptzh60X5geO
S7cJBfTtZnO+pS0VHMlJQRRApLItMY5mIxns9hPGmNeKAtJHcIm2WcvxCKRcgMWxQ5BZs5rWyFih
c4OFUN9O1rxqWIbV2M+G+LVJ4in0C355vgzjY07lhuZdmWFqaXbZn9MXwgn+3rkOcHsZ4QEea/nO
4yyOLb0LxKgdmEuH1dQgPIJiUOLSMO9a4nLNtOpc5r580VE0J6RvhvK42WwgJJYDKZgJ0VTEd7Uy
Q7wijuVy5XyOJd8e7Oekbc8hOwXCF5ffEjjzi0Accx3iSc28agiPiGlF2OczsslrFsdddIuO3Eoe
FBYHwSsqV6ndPpPdlfs0mgjQfEac80YvTjijj4sDaeVQXgwcvjm0kml5mxyuOdIchudjVA9BFqs7
b3FUsPYIUY13+igxnLCIQWJvEo8usLwoeaootixm/1yUQMGeHZOzju3f1Y2BofSp9ZKrmxRAiGKF
jaz8RSFcbbOaxC/DHi2Gvq6W8UQojq1Qjh9r4wiV3EMvDgNStUPbu4gdQRxFaOVoVX8+70vFEBMe
2hGUsVVffiNwv53W6Q0XJocp9rWMc9Rb90XXBT/HVe5+dHhpCreDbAB00tm1buD/73PYq09965Yp
dAxr6+ISKiNLl7PtUVMc/LOvjjj4xcisZ7H8GSH0roSAzjHbwYqwL6dNBLsN/9vfqpbxsMTcOCwU
4bA/FEUZFNRd80zYfjjx8qrh4dugthVqKUkFXUhhgLdCjd/gyojo4A5diPOyiNNymxIylNnfvFV8
OvMF3dJnSvPQ6ifoEuPW9S3wGt36vHIFk+N8mOvl1pxK+40d/KbrYyg3PG8Bg8K0bYWQr0jgqRZS
KaIpBjFw4QQchmEKhzpOwn7sroT171GZ06IIUyoRbVxbTcQ3K4m8ncCJXcoargtlMlQPW3Q8LydE
PaoOWPhT7DDePze3gIEsGI1p8NX4NNOLjGE5KLtLQI3kE3U7d5i3nLN2TWHTZn84g0INp/kp9wve
cV6x6GmjmEG7Odwju3hKe281GGYHxSorWstt34DXfUwLRVW+4uCr7R0HKbAMDVVe8i2q0UBqE0Bu
L3EXV+xSfnNuS+j9n7bPByID4qvI7Ueh36D3N9C9BuBmUFBfHADwr3vO2GDsf7/1NDnUt0FjKGCc
gZrj/dhkPEIIWMVaLpy/I8pPtRUkCvHY9wwWfKDfwfVsA5QKTvpIj9gvYbX9uBa/a28uFvU1pUCB
7TzsnJMaLis7hZ98tUQHo0otc4VpxIIwqxRcuV5YbxJn9KVNn6veL4z7pFuJkHersiblip1+2TvB
3KQ5EAUsXFaSWgGo5gIvf0UCmUAJrvgpE44twzA30nhCUPo/d+Hfsay8WeFBzxzoZ9Q/jpERAwvh
ro355FroNv72oA5C5fRQfpCPVi2CHQ/xVg6EyhVI39L66a6Puo3ERgipwAns/r7Hps+qMCXJWNDv
9mrMZG/pJYuRcx2Ab16jbo8nQMJV6xq2351OjA6JXWfAGqDNrQrBG1S+0esK994MZWdKU4fvqFNJ
f9+tXjUKDm2nT0cc72zvsr0ttGnyi6+tugU7RTcEtwEWIUDXiQ6kNLFyoPo4Y9aYOc34YYLufJtu
m1BMCIHORZU7UH5uKnRmmzynLcq95oMseXCvrf/+SuB4MpUGAuPtfkv9hDPVTcOCQNWF0IrniRyn
grZSj8NNQDz8U59sv49JlUE4n20vJdJ9Ez7BpIgThH+kRZdkF1ZGJ89bFZgl+p869spJl2rUa81h
DTMkMdKGOayZmOSV3Czx5xukoRbJMuhcSkI4WK/RlPWt5V4lcgMJxRw7sPvP3sNDxyheVDMrvSYv
2dFx0OH4kHXFGvsQ+lLK6uvYX3xGq4U1VhvDi8yIQBqO4PuMNsl2YwMMSwQ+s8QM2o49vPhNnPvO
JI1iKJLCByX8r5dM5QodiJ6/7seOXFL+TQ1CMaXj2Gd6kDMpwv+QY3mtfR9HXy7d08filpR7/Gw3
b6O23jibvyGcL/N+ZSk8arjqRcVnz+xjRJ5zDLVkAVI9twvcRKoS+Kng1uIiaobeaHyxlB0kXBzA
/VG8M1t4Y65MteaJQTCZzj1jGRCiFVsOJDPD2zVWYqBXih6gwemMcw/Z6si6TDKJ65UA3VuD/iAP
JJz1OD14HbKbPrpg90hoh8XSb5MegnSRkd7PiqrN5Pl/ifHNsPRMC5QR6F2i5yUnn0xMXe3rU5Ad
WPjg5bE3xpjCc5EiLWGJag09hLrcKrb9aMFUrN6VMVXUFYUerYF7B2uMhGq6iu0bZVLrVBXh8mdq
InwYCuaKZtTHDKTT0rAsru/agGIsXHvsLvT6KmAUivJhu2WGapsxKFVh4IE5ZDuc9oALT8duhgww
CuKVQTlvu4uVUFSt2BqK8LOKM1UU+oOwebsgsVTtZpEZp4xfRZv0duz++S6zpQ85dzpc5DxyDf0+
c1IWxLL1UBEz+pxmI+xjNmeBQsw+KbAoWYxcAhvuPJ45PEuY05Lgbk4cDpUVNOT8wJmkwi/tyCOi
AHej/67SFaST/z+w+0JyPhB/H1lIPBFaBhIVmSCxRGhcPCYXcCVUwR8Gol8utfwOvV32tF4uZ/6B
vArEbKCWoHnd45o1Z4zqMMVIpWCbyPoJ0AGGg3Wx3CIu3ZJw7d1b5GxwbVw64Rw+ZdeGjox0ZpRr
sw6lSv3MoCEx0ifngyVWfA9SNgU23iC8kYhX88JcW2QlltZA3AXWO68uPvdPhBCd1sjmESZoDAeh
9pAYIsItYjCrKlACDh4tXDfgM52oAUdMZ8aiVPniSqcQbcWVxfm15PEmDhHOYblMk13FOYIGgO88
MGm7s5sFU6N43n0kvPOqYx1R7zLd6OrXgJ36sN1rxkzud5b6l40891uNYV4/sAvijMwQGq8stco9
Imt0+S7ZMgpg4OiFrI4wamxdSE+VmHnUihRVbB6YgjYJjFdEEwqUb+ZRFj9L1wNP02K6mXe62V2g
MviJK0XXXYxeeWUiwwrUIXOovQEp2T+tPYmYvmKD9LHfuMJ2bLrBHPt06P2xqs3P0pI+zy6hTzBt
WeRdZbQ/nt1klWNoF0mV+K7pf+jnhS0NWUwTCsBPVn3SDrQfX4h35KJdzAmAggIvUOSmZQQLhEJK
fYrnY9LaVZucpyBSidPCogxx5PtTAtmI8vYkF2nKkZK6nEXFCvRLbt0haJAtHVchZSAifHwl/HhR
lcJvRR8YidDlRYuDlA6wNH1+G8SH162qsLg7+HB8kGPoyzKTjSA5wPG4Ppx+gqX7YEhnRq4IJn8s
f8uTkZkGttle5MLFBnwwx9xvCWJTSbmPUheDXXKrl2rQBT12I00nO1hT3TQKWN2BgjTGPTvdJ6Kt
2qQtb9qE09hHHlpEKFydqxwuyY+o8DPZuGDKNrHq19QXzAaSf+bw25szajYDR8U2izjrd0+cfexR
h6ASXEKc0pyzgF3xGFieTUL3ocXKZBn5QmijFsXJ9XTAg3w3H/i8tku2u8NlJJ4JSpWXMOxcyI9X
DaJwhrZsExD82GQ0X4Urtf+VorEYpVdeV2da4ebOW9e9+K8ZBDyx/JKW7JpnLLiuEtWU/QtjtQFO
SwMs26uEnBXZzT+mP3Z24fz8Gel9AV9WGNvd/l1tEchI3wJKq4NIvlTjbVfaoI0IoNFXwzyyDKkv
ZEft1hNE4Wwqr/LZZiZ2VaPFNOn0yXFp3eB9K5a6EMioeBU0ZHEO7v0bbcG34sobXpq6Df9WI4Kq
oNuZx2TvZPBtT1FNxXAESDzySEDOwVbCiUHRoMW53QcNsGOjNV+aPgu2hnTSPAhOAs8xtikRdUky
XotKuYIPpDyLDhNlEL+IUVsNdBf36Yzyw8Hq9HdNU/RmR8JE0z4XYTo2R5g3BzYHSRHlXFQ88lDY
2TwAPAnKPwNu8ulHqzwPAdU4Sos3rkUBP2t9mxoriOtfTwKF+kkYn/6LXGEsNshbXgWFGvyUNcbK
q2o5GAWNrV8I4h0Vp6egEAqCd6M7Fi6mYVjjWs9F4THyqUYs/enQkftAa8S9SEhP+V12vaxHBzS+
LZIn+n403ql5fwX27JmCkSoE6FRvNvqPOY59+pl4S2cXa3KrN0us97IVZqdoplZCKBDJYimtVSb7
TDxHOr9Yv6ofi2Un+eEWSdrbGG+IB4dH3Vh2cuUzC2sbER64MhtxvraHHI37TFemxFs5KGOknT0v
lJGllGQ4wkAgYTpJvUBBAxRhG+5aWlx+C5kAXzBN00OA1nwCEXasxWya4YpcfDkz2QGPcULyktD7
5ygXUfO7Jq7i2Zu6Sjx2X9gikqz89j8hPz0NX/NpwMcXKwD/cwo69SgAmGUwmELGWjQLGRdfDFyG
pg+6S9oFZaS6w1HyaUUHHWRn8G0j2Yl4/F8htTzM2JV8gdKHhIzxCitwbPbP12xat4CM9X4aefnR
bV3j96qwZbPa8K31HTcgEuQ2YmkReBMbGqYSfpPbUOsBzfodgDlwifpvDf0qKXairlJcHdOG0jWW
S3q1CHK0wGPLLOCxmwKlYfuhfZDxA+lBhtIb0qDetfsSzT8PqiNoYsGVoxw/leFKHg7Q1buKzzLh
XMMZdPJobI7AVeLR4yhlrYdFl3Ly9sz8iW0ltOZWLSNwNqQjvAyqy0Qkn3LCkkeiYeXFxMS/mi9w
Du1GpiPooJdJ63NQUkDD22EIKMbvgIdcioZ/+djlclNRGV9oiaosF4/gSEu7vIQ/ThvblYQvy/Xv
kfRAmmXhhHRnOJa81+v51Qh3/knST1u3ddhknTVpWMq9rFyDNWZuTAB5bELiVzIEdnOJUa37Y/Kz
+QmPkMsIuqz61oTPSzDxE+vSPhwTbnrgpOQoQEvFDiACo4eqiXr69LB1k2WHjAIJEJw4WhMEEm1b
vZIYMJzKVJtl34/qQWknNjNZGjEv9+aNRnQNU91zpmJpM2cE9nFtmSL2WA7zi1k0lTE0FFnBBLAy
mu4XmM1+JWAmkMstefdO0l1KKB+UrIXu5XATy6pEU66iT9FlKcxSL5tKX8tLt61ps4ZP23MVxJ1t
/6Gwe4tsEL+eYGkqhfej+ETEiTwI5ydvUdyeJOdpwv+vg2zfMmvDMAdzcIBz6RrzXvwifGBeQgfY
hu40drxWb48fo90tjvgsjduwJc3V82BydHegJkE3B3Zzgc6HwcG+cb9jWmx7I6hW6XkthDiOHhZn
EIZYj+d9E69fgURJ/19IaeJtntF6Hp91qm4CpYxcI9gIfGXlgzsMXD3MybCkPnQ6+BMkzQh6vpvp
75HGsLonAd+7ObXRnwAXUF6eNhEyzoWa5gP+brXPKACLHMHkUE02Vdw62jdRQ7Z/9L2WNJTYXDPv
3JGYGiCjpqc99hf3vwkZ8j9HnkflwNWiRo4gsT+bafi1yXqVYX49/JRchQR1/QXBVITH/qMugjGE
DvXBOpgbbRzcliNmTlomwNO6Fh+dUSpDsZorG+nivS2+kUeLFDcLPtRJd/sdwfrtfVCzmayTmMQ0
vaMLHYHkSt/yLYh2SVD+z2hdR5lzNdGd8o2C1meYLnNl9JRxKkhiEz6b/ydjjzMayx9OmAq/03ZG
5ca8+P6/d0Hm+dHYNBfEKlppQRVz+CIACCUU9sSBG8RxkJVi5jzH7/ynXtjxvsrMDFElV7LG5S/b
MZ14eHe0FxdSsXbrNjoaTGoRiFoUcP1LpR+15GM0GWwNOyNslgQBDauBOx4gtVOOg/XPbhKmRmC8
qN0ZZ4s0z362K6FJkCW028ldxCm2Ko0UClaMmAMxu17yYajbYRAxG1tmRdTuy4DAOW1nPfoJPFY6
6BolLms2poINoFJT02dBslepCV8hku6EQ2eg3OSQsfz9rvC7u9z++gjPsh57Rq/OtK3EJiCv0qJh
stDsH4Do3qjV6UTRD5GbzJSDMP/4th42p0WUxdhUulkKFQ60FZ0V+PFM3GnU2wouzQ4mQ9Jvl8u1
suit/+i0IFj9Q0IHTs78szQ4xuzTAST62akVxLmSvwL9I3Ixr6DQ4GM3ZcW/RnPdsI6DopH19TTN
8GHtSOioftaqt9ZQuL3EH7zyHw7qOwOHTaGtFaXWbgWZl4ITwuqn2KqHVzinHOXjATRXwphVQOlj
tFUstyNQz4OyzVdCnRDUITIhm2C/iY9WJdwAP+PeTSok9DRh+2V+CPS1ylSZcp9Cdcf5SmZhNIM5
vKZT9c723hWDlShpd++6FweejmldnV9iJUAqvZyLIA4cIJybDZ04dcFE9hJHwTnDGIMCIivzrzUr
XwdHcR45kauSeRdBcEylaj4P0gCO/zKnD1szFSfDcrV4A3F34R6A0irgUBKNu2VexEDdV2opb3Zt
k1E2wcoM41yHALYMoxx6ki8xiLyGBGJFA1DLpN/4LqVKgi8nIAXcfwzuEAK4rtYTmU3PYyXOZz6W
DbgzE5/p0Xx8nvN6oyIeeZIFseFL6tdgE66WLC5rtejBYrxCzOWl43WecpOwLNBuyORn49i8DCdA
thPqWSdGfSHVMUnY7cer9fUIkg11BBoc2OrCijtPpiHG43ozWnQqVrLNm32Vjcl28t0jHUoZUoA4
WmQICzB5vq64jJNJG4NXDBMY82lxeJp+SKhBL0rAetyK1gln+eOmlquJ3DCG22dFymNYwIYAHt21
dRcAFDm4eROkao9pzAobchMETJDH9OAdZqAu61jY9wIcCvKVabwM0ks14JYWOfmaEDURO9PSU39l
cUDJh6nO6vvEzAlQmcy6oCPRUx2RbZie1VS4uvkh8565lg0reqEekkcszVPlOOb5zUlAGXNSugGN
1lwwvrn3e3j0rGata5xdcWj6k3Fsa+GxNUNVNkUTrUpanv+PA28e4w/Vm7SWVgevVQee/IDz2B1o
QiHl81gZXppI0h2WvdewV41V3bMrQfBcSD4TV9Pge9ivcaweMnmdu69ikH2adI9RreaUKB8q+Y8s
N/j+C3OFI28b0kTbLPoBFOgXnGB8dKRJmLzaMrZ9E5Vq5/iEs2zrJr3mPfgAbkqMpl/pRmfbavj7
A/cvVemjUnQbTmQB7yNfWt7S6SWLHrbKP1YfkfFZM4DPvYLV+oFSPWIDrn1PDwrSwWbnesUyuMFb
iKPVSVHXWa3G5msvhShl3fY9w54bVCgjrhfSP7LN94BzvMG20+9FHRWBdcrQBZ97wFCKLFMam3Zt
EQjJoBkm5itzdz2nfPXSYU3EbHk++/c3vZG5S2ShFxMzGbAhuJYk+F3x/t2znmGzvVUVOeWCwT6J
9dU/VGyk28fvNZNin5Yw8Ot4tExUoELy9gFRC0IiD1cEVTE8aOO+OVu4eWH4Qy4g5pqSyiobZJeg
BjvKnv26KJV8BJsvsJDTmn8ppZlFBeofFoHoXHU6YU2Xz0z7yz0Y5tpOUYvdrXKWkD1IaE1uuSNI
WY1EhkICQA23blXoJIOHVO3smIV8gLyF5Lr+ppt873WwvtjOZEO+AYLCxVseQZuaIdb2G4rE8Ny+
NazVAb/Q9HnPA8OJqxr+hVOHIpJCVx9vA5OUis/g3ZaFKDGVrPRrUpujKf+7GFYZppnLYsyk5TvC
pcrnSNfHIlYB1RTWVvAjI/nA3CgfeEJeCzLv65H8uWrYt0s0Lj+Rk6jRXefBwzYIML71Vvg8So2U
6ZASTAyjKI38M2p2024expENTJnHrgtNYhe1zPjs+PAGV2Bq0blu8pHYKIfG/DFEEIKPnAgrc8SM
stY+id7GDynE94myz0IaZREFOlvvLWbxbwqupNfCnfKu7pGIg3nz19v7KdfHVj2rysW7ZpYTbqVn
SQFpG81yH7ZZaIej2KciCT7+o/NSv7Kzha+7WWiVA+bAP3MaECYsruxRBYVpOLX6+u690KL2reP9
+MPPWIdgEstvtKkCMuHkYJCJg0I6Ws3swRC+Cfn1VVWTW2WsCVi4Ud6uzTo8QnzP6MAgyKEb6QR3
Hfuv0GfXwTkt3f01EjVvujQYsxfB/CHZZoz1EN9+WUBtjHzbe91xPyMjVHrxgUnSB3Nd7my2RTUQ
zS5b6ghwUbR8BcRMtOn1MRndf117xAT43JqjkJVPqIVNiQRpLmK8tcJXBH41XtU6PPCAICLldYON
CyC1ptV6ydciFbw9SCQ4DTav+VWFsuWOUsg3UrzjhFc1dSSw5HA8+3X8k9bA7gM4pNeKs20ZkQHd
BUJOKmjo7ffhf1bOedAvNJdDOLRwNBAjpeeVKPm5Gf4c/4raGu8rUcSN0l3Zlxysey63jcm7qSDN
04EUn5E/LVmsct+1Nbs5DCYv6Vc8OvSPw6k5DTK9ESF1KLc0UZZ5inr/FGX/NLqgm8cidL3a6LWP
lNTooD3uK5hgqwEOM6CUBWVVc9iNukjrjIOkyyD4N/beTSxfywPkiaGVUFkfRbQWnVU2z4F6MpbU
3LA+NdLm3nbQj0Kn8jJV78hvwxuC7aF+kHj7TYZCC5o1g21HWSEKRHEUVhP6NvPzjuD8hfdy4OZZ
W75oRHW7txIV5g9DkLLgMok1T3F0dG2xuZX8y7SY/3E+xBSLL2faGaJNwByB7srGkC1ezSkwV+rQ
glvZ0t11TmS/N/JiiQSUkdjxLZDN4VMULoHHHhnqMGy/RZPrVJIP8h7PZonZU4Qa2FkF3f6dJfRm
TuRU3ExYKYaAbUSPmKiN3LaeBJbh5IYWKUO/HPxQ1P5Y6fSG0UDQwGSj47dus6ghP7eZpMcKjT5r
fqe23T9QKHhBuCxGl7M2xeUqLtnpE++J418/CK1iLv7p2p1+x/WFtdwq5tdJj8faxXZnIPGq2W0f
eths+AjSFv0sLr1qRIEuRIDIpWy0NGJC3HNSC1/a3zZgrcTx2Wz5u1nOZOt0JIefaOQrKS1nM5XZ
XivJLfsLK0PgTVvdnyVycXMWVpVcMZD/kvNS/m5jv6Tc7K9O3PVAkrl9EbP+RcsR+Ez6GmLcs58b
dvOl1p1pzoF4sMrRvRTQ/6D7ONTI/4HLjxEn6aaMtN/ripPjEUc3ex/IkbDTyn9mnPLa9wRv+m4I
WrJnxcnm9pJdtsDegK/oGxBXCtymgC3yXnYYCD6imDvAieEpMjvp0uQczmmww4xhyMjWEm1/0ZmD
RhsWJVpKKrL0EZbSvSNT6gCd4FU4nAm+2Od1EiNFilddobN3tfc3VW3LnhsWJTVhEj1sI7iMyM8u
gcJMXjBpLLHU6ADZzlsUiYKhaqa6MXvcXABBbs84JoBmvZlB3ZJ9Yaa01Bi0Z+5fqdw1H64gqAJE
1DcUw/fTdG3IjDXyZZ7pdHBZIXGIoZLBv0O7ZiB5hqAKlVGZkdGOCDHllE1Nlcql6/YaFFUFxxH/
E/b04Sqs7wCmfB0sziJPilaRtfE2REwAop3fstBkaoAjkHSbvNhhr73kDUIXPavXuT7paLOPs6ba
ueT+F1MY59aAwP5ByUuzJKgAEO61vCmF/cNaj1/Mnm4m3kWhMB6pb13/dBgXvYt4JJu8wS1DdXEa
6wJKDK5vCSrO61O2HzqdXCEUKSDEFagSyHH9e+5tljgVAzzueElEzIi6immhD6vA5JyR6BmLa+IJ
MR+SbvbZxZRkBD3o8xhQ3tmtE1sk/+kBuA+RwTgLzs1u2LHmBxzQL7em8mtU96JCuXJ3Shk9GNWj
nzoWlx2jq/oVGUX3SAHXkcu019wdr5NuFEMVk3/oy6h8hVCSO8Zcp+yMhqI997HK4CEVOk4m5C7o
zt+MswZL9wDGUsx3YRyAwRqxvyt5UWO95UdZ9UZr2gol2MS7rD6rUA9lAv6AO8l70mI5IIoNR7HW
thu3iCuQ+XWEo+zQa73aWDGeiJVBqgHHAFXREHRdJ8QNHCM+CcW5EviPt+ahkwgbR2E342XeWLvZ
on872ZnVSvYq9YXSgzKG8y6vwABA7sUy+4VDCh6Djs7tlU1DmvSeovIwbXDe7YmKOLdJuLA4SsCY
vUO6HfH7eSqdLfumYETa7fcL5OqzyYvinim2D+iBWrlKOuWBWWCPA+is1vrj+5uGR0abQAc7S/vU
MXVt0+ABACa05blRkbKG0y/JLKWQridSD9UH1MislA8oFnSOjJGpAcWzmigV1bP+Drl0+iRSFaVp
jwAQ92TJV7E+WEt9uhQmPG/chxa1g7Kdxl1QF7wxpup1r7qRHg8Azx45eq9RlAEoXzylwRAiX5DP
wMTLGEROp0CgmryAUTnqJFbHGogC86WHxYAdxfGqjKwWaWELsBlTdpkQmcxmhdSunss2XSru3Jg6
FnB/mX3qPOQGtKadshkIRFu9EFeklAmLqGRvgdIefmhrdhtC0tfh7KyxWClyIbDACgLPmlVy3MF2
p1W4duf2LY2hqxvE+p8BpdfQPRHfAkMLN0bhmfK3KsQe8oOxtQaKMXL72I1qkOC/RrkKF4gSBK+Q
/8HzfcK8gSEiEf9wPUG0dxAG2teIOo7gdT9ISaJQ/okGwLs55uv2BPux10ZuEj1TFUBxKoSG5UNy
XTpqZIQU5Zdt5LCkpR0W71jpMn+33IQrs6jOVOJz4m5z0UW9uTcqrSNithrNfbwAkQYQEm7YpRWM
ZrWy/6kDh6ZOFv/pev8g2w339SXAW5uITvKKKF3+rjwS4n2BrrOstvBW3PmcQZWhQhnbjwu1nCH6
hLII5zYS0TGE68WOg+85z2sM3jzJQmwQefA7GGshz0Dbwlva/r68sgBsIoZQ+LlawHVX6OPoOcAU
VNKbMkldi1O9GFJkoYqcCJngt1Pw9dh9vgtCgC6vgo3NQ94amaGKVmFTIzYn6gtCcAHJY1fNveJr
nms1BiRV9ODBf0i4XLTN9UX6pL0e0omFG7WfKCR1Aix7N53s4Q7kx/h1CqswFyCGxBq/NY7L3GLB
cWwa7S1hQE3kVBpfAvZHzC47iypvn5PfSobgWfNJ21zbGRUiHpjj/Q30sJXZSBo/vFkj3Dgrl1d5
SbOSqysUmuZtWuxaH6tbMlCxCLYxzj26Jlb4JSwdtDL7E3DLreKy8gH8NW8k3/Evns5RBUDbHN/t
Ixi2AZ7CbokvzV3+PJQCNBzrd3X4F/ZRvrpq9wPoHrAtj2Uyox7v8vqK/Z1V5motZeeok4H6byF5
hwcesZPPelOvYmuBrNS1ox4GuhncfDSE4PWh+NIfNJTyh8qiur9abnbHzyTkYJX5j9coMFU+ZnEY
/FYv4N+F+6TjwZRVM3S9z0JcMfDXy+edV+4OW5ygwIzVkZP3jqGnFGRKdcOboQiag8szQX/FCXyP
INpT4Q4pCn1/8spEAkc36GL1ffLRF1otD1B2KIpFEXPA1bn5IluYH+256PbclTpM2rPMi2j+s6ck
Yj3Uj9JptSnDRM0MkrKKr6gkXb+or5YZnkK1e7VoDpoZ3Tc/LY0DNu7Mtl5adEeo/TGgac3ZjBsU
/SKP/ExBd0GwEyiM0fYL3SBzSKwAuMa5IdnQkAUkrvOp1Q+HMzy/ArA3Yx1bNjssRdWkQgQT/opN
WYa8eQIYxLE3uGNQxdpSJGJER2Mk0kFyUCZcO+AGCz2SGqqk1LrTiXuKNxLE6vGmFq0HJbV2MK6T
a12SrJqaPnuzBWtjLlbLjhBgN+MO8DWNDVKWKUWxay2YQC2WmM7Y9OS+O+rpIlLq5vE1xzjW2omt
V9XOCKh/b0J4SW1kGoJs/jW8bcL190VEEweSKjB7Foq8ASsK4VY1EHhIoa2ocyl/Sxe8EDSjcOaK
FS6YE6ABdd+opQjP3VbwSVgJ75NLYGdMJbQDLtdLJdFnAIQOTclABiqvoh2nrkGy1NWU81U2yNaN
9DvNuJpdvT4HoXTi9VQPr6CPVOqd5ovOgU6YOFqMVvw6lmM4GN6bTegPPbt5eyyk/obTnrEZ3hNf
1sd0fHZTPJX+JBCSCozM9Tdy40nsT6A0qxyc9FI0qYXpHeSDoRpiB+sA0tQ4R+t2bOWBSd1T9ZiD
99c5CxvFHQBoD0sAXTCa3LZnwMFq2WX3sLdFq3iZ1vq5tr3g/DuSBIHvC2UxeqWUwBXN8XYYOpER
5fE0t8HgJHhNvImIIp8vzz9IQi6tR2MpQol2hiuhqigd4y0YFWzOGjLXfrppy9EgO9fCeSyPh+S3
7Sarcq3AQVtATFr2JFpH/RAtzmy7OKVGrSGU+1Qs3TbvzEpKA197NhM70JJnFUryhGoIhfPv+Eym
OuPhh46kACggqGKsLsEd7y46P+yoTIM/5uogONJDNfmd2r+yjIg8hg3wKhKX43JjaknfNFMRn4gJ
gINctpNpI0n9ctPwkBdiy1gf4UA0i8bR1b6p6x+JsujqkSB+cO2LknW7TLvomrPBMFUtrveBzH0J
HgUl0BBHAZ0BsRHLhDbIoqwv9c7qJjE8QuQsGaZeEne2Riq3hTRPVKPkbWiiJTvnU68qn5Qhk1B7
e0znMTOrUkVM1+hRwq/04enWtHwOVdAmVywRkMoOyTM+6/5m2OrOGYUd/TNZzlnSH/82b6Jy9aL/
fxyRnpcXZvbMyHjkZms/XuVTHxNrOMb1eQStj8Xto1UOwQu0xo1+aEWfXc03HQccVEJ2i64vpNNq
VFBUSY1yR9gKfl6EvZ46lXvhmLpKPth8rJdDkeMkcF0iGbY1zcU7wBPZ30eWVM9qi1Z5dTp+NLKR
KtPwSgJNtPZBdQHlKJewM0KYDizSmNodSAQSgNs9DoKi8jlceT6qg3/wP4TuLtm3myk7BSm25m1g
Ui4aQmdJ4shf6ygqZnLYENpQ4vksKdWNoarQTzVtjhjF8NZmdIRTJVrkrMXRlobq5ghDeEq35efY
tDSzcUxts/KsT3k6ztr10g3t7Ydv8TqywHuHRLyCuHOeHY5F/FjBdVRYuII27JJz2cCWVTxjFOv7
9/SrOFK962PxTjQ5uWrm9CtW0HU14poOxYNigG1Gj3asi/92mFV1cvixTD30hX0spBKd0LduHwRH
OC0q/cRUW+7pfLDfr95CvA2csmE6IFztB3OcqgggSd8K1r6lPYp53zUTzVO/8mXloNTaYvdg8Bff
uaRn1pARn3AExWQllS5+XEinCKErkma4q/FkGZnrnctXT17DzCRt5NMQp1l3/uzg8gBYIaEKV+N1
0PUnLXE5U0vyeexwCSbk2wFtlVXXlDyaRoK0tWL5w77QYGJhxNlqcaFXBDdchxDxREomjXX5bnup
AKu07rRht15AQlPHUMl5RGNu+CbBpPkRLWtDkYT+hRurs4CCacHNWItGMkwFTejAbNBZKORCWiXv
3kfPuuvLqFIUzBnCnKb/d2CSXX88V2J/L02oS8bp3fKSvVykhoA6RZ+qpety4bXc3rLNQFUfHEbK
Q76LYCMBMGMDuCr0AlHjMon5v+iHAL/OdY41GP7rIPSsCH5SW28cs6fcyx8PXGl1NJKCO6ETbjwB
OIbwqnziRGlqZBVzQWs5cgEDTKgDXFQjv3GxMDn8EDpO/5pO6eiyuZVqzszcClmcg0qwHRDP0pGB
ezbYwYVjBuui8uKWvglERok9caD/RTl1hPmves1ow29avJqjO1Z/5xNwWDFeDinRsVIh3+Niv4kS
foMRcAsvyq5sNx4dQgboUA9OsBhNKE8BO0OGogy98DRAcdvidM6F8gjrpwZs1oZg3hPsHGZo9K/l
HjNFzciLiH8rOH9PGTNhZL8YomRXn2vQZ7uYCpVhk1gGCZsZOXoGOudL+sUrPapUhBq5DkfRFPio
oQpWqlFZJWpLp0RibFRcw29/+bswbBpOJHS7EzDoiK55wb9q2beHTdAk5Y/WQ3IlefMEkjVpifot
gct6MeJGQaQdFyLTEL2jIOcoV6qfWNYiaRtSdjwdniEvlRWjSXlpqr+5S/lOUPdSjWR/LIHjNWyd
MQcFfktUE8kU6eRce+tGyGozCpGKLLD1D6tFK0tGF9xE9MoCrIEOfpVbQAq3uZtXNVuj04jGNJCr
iGVg8NWxTbljwgnGmPALlNZYQbsHZjHYEiE01eG4llvifVmdm7wRhwK7OaTCAzRfnB2rcmlwFqSU
KBwhnMWlI36lfsC6DNKJzoOXKd+Jilen7CTgOj2jEVbaV+PoKuAXqi0epWoabwC437Hpz8Muaj6x
e/s2S+a8YM7Hud8VaXvUxpzSYM6DegMITgdK2+buoDGulbCRaqjC1Og+nISxyx/1655kiTW+XVuE
xB0xUDU9cVqYXYBLxumQ6GZ9fGHGSYzM59oO4Z1XCiar792We/fQMMxSp82+AEN0s0FdMqQ29ZIg
HzkROY1unNHTAfABu5lHQm7FyobQbxef0vk4fraT3vp0BvKeM9OPTTgv7fZzQBgQSHHNuJtLN/L/
hLDfPYCLEmdPynglX5abQxemMhudmNddUh+wWouWQbMIGOzwggSxI0JdPJcIJ8eeGI/jJAIIb1ru
Ip6pl7VLMaxRyKMN5sGyOhO3WjNDUJl8TO3kk2R1pn8opWQBpmvXl/2cmIjqboVj1GBB+GgkTg8Y
Hp52U2rRTG0tBa92wUcq4vEp8JrSuQ3kXNhQgCNj3MJaxIZm3vmeSwMj8/X029pn9o+6m1AqcR38
fyxbc2q/LCmxut/5ReGhb4Yt2a6fqnG27hK3LSoMpYasO0ovQemOb+pOihdheanSiAAid9qLdoyu
8439mBbVL1wf7q5gYZRGXrORseN/BM6NXsTPo99vcC26by/fVa04fbdjGC8MjWNGQQenuqLIk2dh
LCepkIdbUWp1Bz49Xef7z2mmvEbTRxmYh1xWQdoyyQsVSO77XJt/3p9HyKadEoIT+xVkpbTZKOTy
s14jdGm9LEZxD8f5ngvZZ0GeOTecdEJT+mN7p3vbd4iFSjmbhZJua5oMVggWHqqgQsfkmBtWGWWF
WA1jb5p6A4q+5FRjDHLzGM5dIsG+GBR5rYMIdZ0VOrbnsJGFjb5jcMW2zKhFCHac3vzuhRub0UN5
252U0TKs6Z9qKGJ+VUOGV7RUdRjgz2Pi9SHeet37evBVM1t4kwUhEBz9kdNwPQegj0KS8eXTuKdi
rbtv8Rc/N41OrpM3zDt5J6xroniAiVMR1M1khjV75eVPIOyKwYSoCEDGfKdmqmjeh7HBQWgqz0He
WKozPWbyJaBc3ILQKHTakLZgbI8MVDkMN66neo1iZlMTPWBiEuVbhsqYu5hvjh+XksSEfnueb5FA
Z9rAQe3RQk5hDe2jcWQU5BwUdJxiILuaLC08WsxS/d5gQiiZOa4CPxQlGqyJ2oxCkXKvTSLsAIny
yz6FQn1xdtUeARym/TFJ4zK25sV0Xb0NdFI+N18+R7H6+hdv4q1H2whRKyhxSW3G2/H+1QI2oYnQ
KcVLus/Z9uBCpCaY5U+eEj6oUuNngKpHI4mkoMxEJOyUIHpS8HcgNqGdzMoNk3PKfhDC0tjq4ut0
oOJNb6n/1Op1JYY8nX4JjIvcq2RyiGJYBfYgzglKKsarDo7czjf6alXJ99DyYJlMpPmIb16KJMJq
aAJKcWBJqmjE4fNIl05kUhT/XEO8nS1Bbzevhlkvvvk1lv+X7Rt37Fvvljxc59BsvMFyh/XwgJq0
XJheWKb4MLNdTY9CNiFOOsodHv1w6Rlg6/GAuAAMNYeuZLaKFjHR2jOk9CxkaSMpUKRoj8CEirQx
9dqQ3WA82EXTUYRIiNYk+2QFvRJcKJEs1N7hHzTUpWMEd2zc+dwhY/u9GzI57okvXi4BXIrCqpzx
9SBeYbB9jhDCdaQvxh0cunYuYRIiMxykxYL2Up21INOaCHj1Q7GUeu64/cQuKrfecW4YeUD19a8t
GZJi6qXKv2yzm6lkpkoybsQbwco+qTCkSHIp1txRI2AUFBnnK+Wm6WcTMM/M14OP1aYtlQ1iwMY9
PM8l3OjdDlXFBOQw766Y+wFOEhylNGe1qrQTJm6wyu/NF8smOG+rfGKiXi0q8YK1xZsVa5FdiOuV
4sifSbdrqHsScQDJLF2b/YA+owFrd8G2d3UFajMJCIpBHavLQ4czjswHXZt/bbO2CW43G16185mZ
48Lo6CruTvlEzIcJr4bwRZG23kXP00UoKjUWJKF742jQQ0Nse6Bv13ZS+RZX8jGGhoo7C+m3h7FX
B+XipC4vUW+9V0GGiYTSglLKrBFtfpn7cPmfmi+pVjEv8vORiTt6t6ATL926p0m71H2NkBQ4Hujk
dfNRVjXNhESgZrcbpLBr1bHNj4aYYYpQZmJU7OD9mFe3luPBsDoq8xAES3wdLLBGcwA9nMK7HGDA
0oSxmpXBZgcwjtUEnwjQsdxINhgVfHGTcAbwoQ8AEMBY09/WsjETffjbq35QJDkKCA0XSMxYt/Jh
OTbkFAVX+jRAiOgrCuROH7II5gidkRcYwtdcc8rSdKCaPzpQtEXvtwfVvf1uL4hi6s0EsWe5hdxO
cRxG3Nmx7iX4T9td/HAG7mIk8B2ywluu0Isu1mLyEwswkjGw1YCNBRxAy6akQgbxf2i1IZX4Aprs
zZeK7+vLCJ4OTpTS1K4vAGI4qw9uj6umcLOF4x0AUrXh146MyySG29DmRkApdbxentpteTNyiX/z
Umj/ZOAXVW8dux1ocV7W6jX6L7n7nyXGedIWmIHvvj5itKFUtdppmIH89BOGraXe451a590gZ91w
1fF51vm0m8ZmuxYQzOlNYbMrXcRxRqUpdO+CEYUm9psHB4dY0yw50wPKjD31QcroFfirO63d1P7l
hNqX7ftKuZ2As8Kbc/fZbwnhz5rAY+tBJ0CI5ys/a7SZJxGh84AdH3L6OOwjf7XDoodNV0Hbn6YC
XcZVGsYGV5dAiAGGvkrvvHI8PkABBiRia6In14iYW/fcXtusbmBhukSQ0FjBo+rg01vuVtnNpTUJ
F7IZFCZUPBd29XYOWGaCXLAeVGjfSWvPLevBTChmceN65Myk1o5AI+RB9B8ea5WrzbzAOUHhOc6J
hw5SWLMVHEFlOxFGOpZbVl6ZLlfKCOmYfvCjjRXi13l8edT6XVdCQ1m+LayQy3gfmp70UHNNiPmv
XsfHZxeMZ6kEgfE4/81jbmIZeAAPq118CsbzXT3enJ/xX8h+879DxkkVT9Ka4WvTqrLIFJfRiI8I
kYo5ux1IdXATcRLe3qGfDjJQr6zG9E20hinptA8O6LbqIxRzPJSqgXLuMzgtgThHNK+n3ieLfPig
zlYhEOzsMsX3RpUVDrXP5HseAeoEyoedSgOFgN8lSbVYLnS49WkScmAekgw5KrXH6JwwlYrpCzvn
8gaNSf9AyMe8Vq78GRsjj1XYTHJqg34uVwvUgmiAoULC6lqEp9fg4aCW/KsIPzBnUgr519LXQenA
dqCcAGCBUyp0//z1NGm1ZO8qVFDpP56dVc/YjR7Lgb5BUFlmjyP20cou/4yp7d1y3xJbNmFEWvI7
GsYHeRgVjCEzBHjje6wYfJVgwgSzztOvVImP5RWd/AUuRgB0jhNL57DIYycVZqmKcnIeVbS2I6FT
kDrWmQhoM7/B5B3naLhkJTKc0OZwowXsMji2FOJQmFV/X8ug2CUFehMSFWqDD0eVu2K2FjCrg3wQ
decXCk0nooyEoVk9nNg/yjGQGvzJcWc2KnzgJQOVhKZkIz+q1QQ0wVdL24Y5ZY8QKfB8nq9HOshB
+CohOcsXkKBDMTlREhZMHLo36OpJRCbaVzjDUvtzM6QxJh+PK/rCXtMRoVM/GGsezgKwAVwZMrw5
2lTWWkdwRXFnv71Q2vCNv35SE/SM3KuldI7u+sroevHaimVLjOqgFkKZKEhJlp0gJSb2xtU5mFBg
YvYMFZDgf8ITVEjSwd1YJAgDEF4k0EeFMDpg2qsVC+ADsE8P5Ns6rf/V7ZXTJP1DUeoaXLt9MXB2
qGrB+CE17zk8LI8HNyPDs0vIg2+EbVjRuxIzY17qVpMOZTId7/QfNSV/MrKpkgkDO+t0gst6A3WF
Yo9LjAcT/a+GupjnSveIeGJxNywqbgKZecunVhCTgNQkcS1AqRNDWpztpAB6KpwdwWwLtLQ1R6wM
RU+MWuBOxrDcL6BubGg7U8Yk9psVnjd5AGX9Yfmshn1RiJWfQLM2uT/tdlU++5UsMRXKRdvdcc8v
FEwnl2SOlnEK5M/imj2CjrA4oxVe9RJ4QkRTro6hR/oarf8lZirqPRArio2S0+iquemEQ5qvi+xe
OVffPOeezK5zyr+bYDGPu56mlDPB8U0hEONZ5Q2ZyPfEWN5EtPhcYuyZ2nvmROxKsIeAtGk28nac
IPLzde28OdC5LnAAmWaoIbgFFtU/B7l6S/eGTaBCflC33KnwbUfnKN+zZ4GHC9jbtWSgo6dB45e2
5HSW0claxihP22I2f5wpRo5hF0693MGxJSr0wrdJ3cGZQ6K+gRrmK6Gns+7DnHHasHJNFKnNigme
AxAlV9aS2a4Ik//P4FZABMj7gJg45U99lnG+MPfWzjmPgbK/V2C/U0TelJBJqVxxPl09n9IO+OAn
kAUhvi/yVKHK7C4a53YMAUWV+XCpcQ2OuFo4dHewUN70Rwan0A0lnL+i/cIQ+/mspD7peYBUf5lz
QzcuN2aTwYLPId2Be4ZQqY2+KKe4iH4V14HELdp+sUG6QlU4JPbGI4XLKtEKFTZBuRkJSfxRtBar
Rwg91oHp0UPKL0CG9mdC1E1CoXfQwI9QLPgRESZF1ceeG0j0XN0pni9p10vhBe5IfGZaIlJR3RyG
Ep/hDT6yToeUlqa1Kix8fxcUxhq88Sa9lMSf1qeJSh4SDJL7OoJa4TBk6/jans99xgIOyz5i3xDj
Im+6V4WkoW3VoaWWmL59dP1m15RN8iMmM73Ihdo1Jy7zKExAbUnN0DbDx+4zi2r6RfuIMHJPSATE
FiKJecbU+jX035ChN228TJZzW1x5BiRXwRXSHm8+NbmcYbxMvvQmBz9TXyB2+W3fCxGA31g2QkWC
5KLY3FX9nV1p4fFDi4xG/YlYJMP5YfXZ1B/CbmkhgSRezbk7jUA+weWycboQbHGTi/tN5JwuNrRF
0wkT38F9+5AW484YdBWBxmhGsOhJIHpj11WO3xC4xTbDvsxf1VIIoTrvyWsBGV4LM+AER0v5C2TI
ElrO45Zbp1l+C1ZylM6GTt3f6TLmpwFwaGAz2Ih6IpH8c1KX12ntqm5tAb2+DWCKz7+dGcOKMzpf
YUct5Z75BhU50XVgRLK3KVpTHP37HQQ6OJKAb5KZRQq/tgaOSuqvfeEWYSfBSPzBOXrUdJOAEhz6
U83PAizmkiRuTabx0sRkht5ZDjRyuq02Tt90PEerL/oqiwvCeKMagm4uyKHrZQ4mqoNi1Jo8BvEH
2Vpw5yOoMUkk4/R2BjJ05P+1ISN1/1Kgf4TEjY4t9zkIvsx3h3Vd3T8nnZJBmCc8QASKyhplsXj0
zuYXrHYts/wMbdSD6LFFDqlPtUnS9AgIa8kM5hfo+UasmkMG5M1hQykwRpg6udZYXJlcos8eKme/
XiHsU+JXW9fGIC5rXmZwOC0ctwzAAuLiI83ZmRdT7Hpdjc+hqF+sGsB4UYYxN/aiSOHwKrhxOgDS
NsLdaPVG9cWat3GoauZCYWLl8QoU1tTjUeQrSCYf+1CorfDGH5YMKXzCkIhVtzP/E9RpbenL0cRJ
tlshA/RYGBclMZUrjYfdD0HnXzeRFvX/wpRzcTlLuQ4JB9n5mHdcaRv7iBVdPAD7DIC/+F6uDB7s
29G7bKLg2nojFp+Rs2yiI0GiNEBkpgGrjlnAT5+CGiMnwSob3UPXGI0RhY9c5vqfKAhAk5lwaxnc
WjWf6MCSR0SaF/AIhKohAokbzfixOy9u2Cf4Z6bwe8BwJIi9HOTWo2CjI5BDvvNUJQyDWJKDlyUz
NcqESC/h4thUYVaMCBCxBfZWIUGQ515i6OsAfS0V1AVo5hOHkv8jPGlYSwlwgKdk+mfsfumWKJFm
6PcrEke18iz5SCr+t5BWxwooI3RgHqrrcKIXGL0UXZK54eUo3gTyhcEaH+b9/ZDQQsCp0fylb6ow
Lu/m18JW7UqrI+/lrJuBPQ1bL36UavKqYgLcHq11EqnFE+1V6M0bETHrZWcK9/FSJwLQgSz1JL44
aks03HawMQVSQ6ll41z1WClfthY4hCgDJSQ8Po6H4R2BaavLnBFPvSUtiONdBYLiQz5GHIydQtxn
xM6cxNT4xP5CKFoNgcfOjz+M/0z/I8LTC4txWKMOsxVUqzB5/Qw0NkQNoT1M5k5huBK8i2+8uHKl
15xu1c6vssiaVA/xUDwkd81SJ7/2rFAFNWxIKTgSSFeUg66n7XPYNQH7+OG2/h/23QhJ3GgmzvBX
8FN2hCCbc7VKoSETSd1iZyWvsgjsE42rm5R4CV8bJc2YWBnGQjQ2AGJpRt+ryGmdnRP7JeHCb3n7
/k+8lpA6MeUda21ob8YtSR59ZScSHcI74BNTF8xPPCKH148NwhWG8pD78fOwe67Y7Xj75i51zsoi
mKhJWjZRZvQMd9H1lMzuzfJAOBNCTYANVAROGESIUIqs5dhj1vkLKDgw6E/YQKzbCziY8LhOInkv
4poQQqDz9vGiVJ6Xfvmy2Od86+U/K6xrHaI4IWukOeNHWC+jDyvss0qZwVQ1FNW4eJuopw9K0Tjq
8kngWfMF/yCY1eshUvd2guR+v7PiDilRzprK1qMRLYm9y9d2pGoo5+RvawiBT+FXi2/yNSM+2Vsc
n//WVhKjL6n+TrL3RAE80xRDT1D98CZ6mgP7MOLO/cKCqi52VTsdbhxSr09/p6ytEIKwM8wbOlMY
q7bz5K5rO+d1BORpX1iZ2MV9K+yBE9aLreNGw8OOMKIjEGUhrR3ElOnrIFrTGX7rh1DNTtHlayU8
esYQDhRnQgRx+GHPxeuT/oFR60ZD+gpTv+8CiV+ATP6UFnWqz8qZyQiv2TcAe+s+lDsG5PSaU8Cn
v3XXFcBo8n/CFyPARCs4EPlzGEzls3iOvx2dcHaBsT9dPZklf+4HeKHeWNVTZbOgeSlDS1VqVt2X
BEVZ4Cgc9N0pQGCykmKmnU1/PKrPIWAOOg63Wzfcy4Scbxm3NyFyB9H4M3f8Zf4Sj/zhyraGyuYV
VH73VF1GEL67XjPaLHwYN23USDwiAFrsMCsR/t+rxMfl5Ld4wekXBbzuPF61X1T7JqBuataDIM7E
pAUBVfDLCyQ1md3L5g1vzQLz0DOsNCDE8jqpqa2PmfWo4SDmQo76Z1uaiiBrKuBcT5tdT8XCqODV
HJ+ecEq0EKBoLI8zseY2IPOgGZQ1EV79stfGkQ/LZ7gR7NkYHHEu+Y9cwTtEZnTYSEQqRbBUkHCL
fZsXI3Fw/2Xevd6ZvgBeABb7KdhNDViZZAOtkbQPp8YFiwp5Xczz0U7w6iBNVTmYZe89CW7Pu4aW
L5WueGlBtPsPBOOl5Rn13Da8+taUjBtD5mSb05q98gfCkHJCduWWaok43zDWPvLyFECfS2PLvMdP
Z7OOv+GAoHW9PD94U883MuliwunN0ZefR57A6HBLuMOFcBtFa7DojksOUC0NzgxQo9DF3KPsJ2Ct
2J/XYzBcpxKFkDjX4FosOzrqeGyfWlfPUUlZLBY4Hy0bUq4Yz96VWmHrP5QZC8iMuARCGChd7YBg
3Oml9+pN/fER7JgKudfg3+zzfoJZkULrVqRiVp4uqdWtf9O2xhrZqRe2jSSIvxwOC3VIaUiiXBg2
SUDAVmAJFAG6KqUmmJlKeXG4JNTK7fI2P6B/NeJLCJ2ZuxkBQZ+wgns1Lex04VXYFv2n4ZP7x+HR
PcJucDjrvC1vxnr2wcrt7/1+7kD/hxCxXjRrrJE3sY7FChPcztXvgpGs2+8axwYMmNaTKmnasGM2
45001Yho2HkCWpPJCnTFzAd4yNNilKZ6pPW9W0HxFp2Gm6lcYf24VGrYJ6tHsdUjcLSM/LdTxuHp
KYmBTVJJ7zqK62iDozVDcoiRJelm0GWKOu2YTDexkl2zPHotOvqFD05I7kKg2zqJ1WvkTiw40Z1n
i/zbSL49rHe8Bj3fWerm7HuODS0o6MVvzLsAfRJuV3WNEzE3mS+dIBQ3TfBwyApl0iGR1XGipeEN
urg6Dagv1afBAveBSSFDzBusm7Z7lGorY31wSB7PuU1jlX55pZ61dWuiqaPCF+I13MNhcpvRKtFt
IdeYCtWwhRDVvIiNJKXrSsVNIalwknJrdjZlBgmsJSuXsY5Q2q2sMrE+hZLT00UIXpHN6gEExFVB
vcJogh+i7dDZUxNkbzx5X1n69E/FMAtxBcvf+F+lUjB6E4QQhe5DFt9i7wqzfpEogMGDBGdd5+MY
PMMGf4bgFRAa0tiXCJYNDpluNHEJQ3tkkx1pojg+V/DZCl2ii4MLLowrSvNphJnya5n48yi2F3th
mD4riHH6bK8PB+mtS6QhdhN1FMNiXneT8B57IWJLSFgfsigF324LAyhI1VqKou20YSljLJ6E04Wi
dwsOUSqrC7zPQal+7jvpSZNB2Yw6P4Wqe4A1/eP4DYCqIQ+sA1T3nyEfUwwgnYgST53ulVqTplWy
XI/goU/g1kWhgWjnLshLHmIPVhx7X+vXPc+4L69ZUGuFQV27rMiVW84FiHjFgGu1ht+rj+esgILu
ctpapFqZ+kD2epRsh712FJbbDzabdOGtuzoSkJz57mOxt3WP3SsIXxAjmwPfdJ8/fiX8olTPu88l
KigclEcB7MtEEgiquWbtYY7ExtuH+SkkneePSjiFfp0TSrr1A03r2IRVBT3aKipccZPJkjErvE2G
sJvro6svNMrRxPeTM6qr8mj6USyGHPqPBTtFsTRY6tThzg91ERu2YTKE75Egj9vAI5syY8x80WGj
6fsgmIlirVez/B/dVnrfYcf60vmNt0i4atMmtJTdvVvriwwX9gH8QbuXS08ICVe5kJi/fAVYlppU
mJYwSmhGYqdB5VR3leEsoveVUiVRshul3VYPXkRd8G6fvyOJLptzxPn0KXL750lyfZn7sK/K2klD
LDh6ewkM2Q0f8Ri1OU2uI9dH3ahWg8Z/NPncibmzROsVCzl/jgXThY00HxoyPQ0hXjilbiFwhVHW
RiwClE4wxBVSSux/Wp0zMpvjNcnV2oUXLDDvvCngNtO9qBCgW9uayRTwdcBq5iseMDemSCQ6CwI+
AtV1RfBYAJEYlaaql/4qkFChvNyG4arv/xwcm7KxntrfLuAY6YUpiQ+vunDtPeIhJj1kZW+3O4vC
di2iYHQASr4y5GcmpQFnQQvI/CqvSL9Nj1Me6XvuUhFnXCqInCXWG2lCgA3VqY4x3zW/ROb8fPvX
1m0gGokeZA2c8aNydYm5ftibRx+M/M2GWmqLP8hvhgGaEanYs5vcxAk6FaIH8arCSqQ7Ir/g9KJe
OsRyIG/OD9103UU+Kb6tmSQoHEFiKZNW+CinTv+3FWibwbqTjWHUBDL+LVfvoJg6ofVUi9RImTHu
a/Zpp41VscOJo6/33wcyONKdooK2S/L3p/0PE0Fvmh1S8w49Cl3orQDRH/ntIVElS98LUpf5cQ0I
C/lctecngciM2mAy+Kv5kojiUU2rP/DDZviiyXsHg36c1ICkC/bZ2lXZ5Aw5EJoUmxXTMJq0JDAt
5puvBOoW55xP0gMags6tXAaoSek+redxEp5nW4YfYV8cTZbQre7SxuhEKcy1ReoxJJ4jhH5ZU8f5
5XOP87gL2+SBi+fb8+bboXdrSFwF7gTz9SmJqFKvMHpZD1hIThjT5lMxN61l/bTT7JJOl7XvynkQ
mFZfgPlJqU4/uDOb6wnKSEBga1KRIde0DD0sE5U5zRIg+fn8ZOSOIQRGcO2U80fBGlQLq1eXnFJj
sgg5+ZAmbYgE/nfr6aK0owO/ljWJL8g9EgNeOztYBzwDsgHga6VyxhWT+ZqkFos9YfUS+t/uWSGY
KfK/J6zZVXVNXWQKPba4l4UezkOGrEUzatT+dKZAjeVgzRM+cY7HQoxLDX7cg773He6jl7ZwQI7l
GWPxLt+ifhgo4rS/mKO2tckKaldXcYBd/n0/FDp1m6MxlSgd169QxXxEW0EXkTNpWqz3HWK/Np7v
stW+3NRtQTEMlvChmXqjfVnBW7n1QmppkwEJBQZLrXIPlH6+z/KtB2Hk8whkzIb/ryTduiEgcUdy
3k3BkB8nlWwnhnvTQ+cOG2mkTB2KcBm0hanT+qm9rTHAGC/vLM1klX7mdIiksiGhEtcUptDuGPjG
LmKmCNKiAAMa/M7WF8r9s5tjYx40eUvUvrr0V0+aUFHyRX1vLzRvT3ca1XETMtXzTgOPrKgym+IY
OM7zdQQYXkGdZSrWxWXKqRv5GwWPVeU4tYbh6eI1Pj1eUkxWe4DlFLpyxPCEp9FIOppsyZLp9336
9tVM7FIxGGy07m9aOuwUzigbD+RdaIad0vP+JcfYZ5Kc0saeCKN4TJaoe3ZMsPQ4LzyVFsNyoccV
GDN+il/xVac6IOm9ohdxPFa+56QRu/h2ZocidxQ2wKxpPRokyC9x5h5kxzwYze55zlbvfpj+CjjU
BWv1hnEApRNgiPRltBhM09kre+feGViuteO+Pu7DV89Z1bgH8nH3o0A21se7jWlPhpCmZaBVeQQA
es6FX6z1Mt0fB++Xk8BheQygfBR39y4UnPftQFN7vTlLSTCSY2/pbC/SdNWQooSzLYI5eWt6XGmm
KfZ/9dbRF4T9WI9RVSJYRCE4gff46RgByv0pG/OVx50m0QpCv1HMveIELQEKrBSTa6JkizvtCe0I
xGdxG6VE8DAmhqAEaBFrQX4D6Ng4lAzFw2rGDHV146rXHVa9Tn4T5wE4Pt3oLIvGglOEENvegFSg
kcbplFBSMEyVI+SPppJX9oY2X8jgJi1w3i34RU4GLT2JKlFlsD7Bmg88dxM1d2ACsGQ98RxIcI7d
9pqQMVtzCQ31/gMv9FzIxJ9q/y2d9ynnhkrmnEolt3caTyI927il1tvrSYLogtFqSZsTZScpB71N
c+qm2RZqkxmYD0uMmB0C1Uyowu7LW0FpIvFRGS5mXoAdeV2/WgMldUkmdPdM265QZ4GwdqFR5UW9
2mZK5rwfkAgOqfzBqlGXl19SrwfWvYxmTl2LKfVBhhDMoZI73lrcypMAKE9BBHriZ84/d8OXbR4w
UCOmFNMOijDGDjYocmZ3dJ1iccOs1I66y51tMA+ru50tTQzoBlcw/Nn+vBHWQSToSXksrp3iRmfZ
egGG043uLjoi0uE3z8Vxo/D/yP7QNI45WkFGs/IVj7l1c+N42LJ+ogmm7GfNEXXpboo+ar7pOwFp
1UK4EO8zoVVryeiMRZVgB6I4ZnkOdwT7vezBxHT5JwjuyPVP3zyLtekJ9tLgq9mjEZaCaHORv9II
4PbVtzPhk5tZK/rgsxCo+DtboI2eXDjl0JYx8d7bcJN/elQNYAT/dyRtLIp59aL0lvVTEQqI93sQ
6+VilmldXhGH1mVJrjSQcZA292n0ips49wuYCYi1hIs/CsUsx1uSzvitXpvVwY+T+eWA+b4sEj54
oCkHEC+eLueWdjySSfEmrhVnNhPB0b8Vxt8/AGyhz0TDbBlY6txfrbEhHAC1D4oQsHMqh4h2Qkrp
0AdhKDU43XlSkn/f/614DztT/WjRuEIv7zF190BqYx9xmTobCu3UvXl0BO8E0pVKZPU5QPngqMxg
sI1Dj2zgM/x5vsx2R4K7nFKFMlrX2aBxeLnV63IyNAhkgyi1FUbJUgBiHbQF2zhoATAzRD6STyQJ
8Jg01qUin+5EA/iFn5DVHJczBkZX6VpQBFN8MuF99/tWlSCNXEXHopLiAiKljp1Z7/Pw/7WtqgOH
YBT69oFfrJAywUVHKAMQr5bxwXsKgQvUEW2j7nZp6QLhSyd9xamC+G/DiXlM0+CV4sHqd+EysjI8
34LvMpeuZd7wXO0cjk9w9Jowd5oU+JFIO/hbpWPCsRk5DaqtAObfdTnW85gW/a2WwStCC1eRu4wl
3ZnEB3YWO8pPju+g3x2JfWQX/wV8Mhuu4mU6ZVQZnVkpvybWqmFBLiI9psUHkldl3k7gH4nHxJXt
CkzNw93/TQe1NdvC7JPiX0VQJbRXMSFX0HukHgnUGpE2x+XRMdYoRIu41zY1sdTViOkb1RDha+4l
4/b4fY9+vqDaIeIo6WFXaxGEvKMQ09g4qrX/qXqrkBgrifApLbG1tJ9umRBxKqY1fzYoOPaISdpR
/F6EnpkxyaJvAs5z6MS0mx6T8WJwkvqzr9Gs671saph4Tn3QfYwTc20WOIzyf6ajnWpSgV0YhzXF
wWj4qMUrv1HLR6YQRLKBJgo/z+txbePiHoZ8vbxELxA2AU9REfZB7AE+uSv6dBsKNpKIzpbcJBwa
scA8dPvyq7UUO9pPRVYtWehs2TzLx26oaQfSR+68h0eqttOwnYcaH8tkw7iuRH3+KgBrAi/jBxRt
ql0H5rzLuqlCz0u4oVp9qrsGbkQzT7kS4FEsb6VOGv4sWWV90XeTF6edexDRUf3b4+j5dCp94ML1
8MOdZAcJ2ZsFZspDy3zTFvAH8aQ3flJAjMb12tjRJ51ZjtT/CdPIzSfpkdgAiXxQPSmd3kdgKEXY
3sudEWde8xKQVNqftiVH2YQSiv5fjnTXBsGD/cqep0beiYcvGQ563taUhOGl9Bz/FFDxeFfFWMC4
J6AbHWHIbdW93fTZPZpsdO7j1E8vG2DVX5GQErcqVSUJoUG8HYQIhpi4NcU9zDYTmEi/JZCcuEeN
fLR1g8ycw/LWZhplCP2gLq+EeamH0Loei37NzcdzkF4AthF5ThoVM1LEF2h+5OlhSsylPfEIvk9r
bmyt7POS5hyX1MSghNShxnQ0bhBNND/vQ2VMMy9fy/RccZinWdcIWYKjztuSO3fD5jgehG0VR5T1
0ndckk8RqDzaGq4GDeeUrJrNqW6y17owjDMi1war9dl+lrm2jXySaK5Rv1B8ofU9TTlMQ8Jac421
lPbYZVFX0NzgVRks8YbZWON83SBiCB/vE7Ejbf5frtCFDQ+DEaHn2kNTqxpwrGOjz6Br3UxOxtoY
8jFChdZrSusmRWHswmDn1iCW4ctoaajCU6WQ76rGr4cZdnWTPJ7ns99xDd5mPHS49cy7jD26iL5R
tf3OiZ63pX93Khf0Rc5rLJA44KDNVcJcyXbxW+0yZ9gxqgFRk64yojKqANa7nigei2EHvtwBuGbs
1pu1JWARmnI97Q6+dqbDvPIk2bIBMFBOj8M0yt7b87u+Bo+st7r1ZEYqM5B/nEREArYnfmOjAzek
x5uEEtAAhTNY8eLqKr31RwjErVH+QLqKFY7xU48o7y5A5THoCg0+5dd/UUjH3Fa9CFl1y7/x1x8h
OnGkIDfkPYREpHC9aJ7RfRi1mxSX5PPpPfog/r8P6DtjFp2yYJ385wZiO8w+HyaNhSoH006WkqrS
S7q0VpP89br8DUdBVMVhiSpTEcQ9nt95UPHlajQ59ErB3n1RGQ+hmuVs+teKFscr8Ijez07GFBIB
KQzaqq4en+DgWnJj6IUd/YYQQP+sn9spw+E6eQ7g48/+IO5RfZcFFQT7BXC+CSPlM9qNcmMtwrWb
nHYN2zogpwc0f1YdUTuwuiSPN+tmPMP1t+4PLa3SOP3H12u1hepMTGcjiAzwGROjBwMcHgmG4W4l
WPuRrGyEJvQqvxKGETN3B5M5wTPcHsgD7viGtIaA/DvOCYWedew1ku0x3O5E7b1Rs0RqQM2AqCfv
rW2Yr8Wzb3g817JqXbVz9Fq72Tyb4LicBgi5ixZevQnbMzfUk2xObiUcr6a7okYCOR/Qkluk0qsP
ZCeXCFpDObJsIhaMRA74oNWc3nXuDomCvZaS6HACXWvEv4N/QoI9rGacbHXSr+gGPqC92PmURD41
arii8HTociy0gdOgEfqcFf3jaDrO4Vgc1+5zGzmwnlfeWjQeLw22/xBvPpOFmI47hKLd6x3UGd/E
DASfto/e/n+rQ+OS3shNOYki8NROL1Nv16AlX/lyUOrhS0TUXR6UzeSyRYMxM7fs8STmvHIzGzKD
lBy6ilPyQAbXmZAQWG7fhVS17bxA96zumRJ22sdTCFe6M7WRjucsOi0YuyL30FtsJuXT7PAffXg5
qKFDVwM/Pcaccy/o1fNgDhXtZKtkCjGhu9AOKfPxeq3j0YWUu3QomGdyrpeGQomRtAnXRmAZcVPZ
L147xv/tIJu2Zu5ABQJCf0Nhc91KelkB6254TzRA3cPMyuEvs5Ftl4Y9/sne8AUySzdwUxZg6QKa
rDakTh1NQUHmNfHpQSBHVLccuoHTcvDO4hreAU1MrAezushNDEiH3W9R6GjLYgD2MOUimQbVP2MU
4ZXmrXY0v5qFcooiFhOwxBEpVAHDkVT5Wo8IXYoqfDy24TXGPihbyaGG5EDGtVfzP0raZzJakydN
HvqsmR64lguoeZNYtRe9t99/QIef2SbQbvCuyeffHIuEys+Im8PYcPlmkEbU/n84c0KC1RpnMw6G
6K0vGQw+WAi8o4bEXrQEo2c+Mz+zc16DQ1hS5EXWj+1aJfym6oS45ijDZy40C3GTyovtbYhfGGnj
Ig04c8eGWazP3mFumS+HmWueA7CsSdPnkF33kseoYZinySmV9t15O2IR64Zvd5/JaXm5epnIgxPV
lapQJpcof8Ebooz4llNpuPUV0ghfSDN63Oo09FphbPktahrP0IyT9IF9VQ5muLrDcloxJr/ttgAD
PzeAai8sBjVv2BJdd3wPLjtsBZh2LEthOafMAvLpvVToHX4Eaqiu7lt5IEpS0ShGhWEV98HxwdSh
Uo4kZzSKgzKMz6uEGstlM+yVutHBqy0OtC5jAy1YYfdSewgkKNGcegvLGTnkYQXgyGcpkDTviUQQ
p5V3C/yZ26ehg6eKXdyEa/vwZS9yq81oTRkESoOCdqqxnqyJsBxtxxaxkDxGq+NLOMaWe7ijKe68
yB+HGqKb7vMaFkO83JG+NlyfHc/g1I/bg6LlTMnwFJu5RdTFAT2+l2OC6etCMPonaNZkIREH4ipl
TuLKSNn0x8VrwlLdaQMcRdiHpPLKmcMszMWRBYgHdtiR9d38meTjzfqaTt5GZ/pH6cPB7+6Svx0K
RRa30cLFZrdyb7e9LqB7qVffUAInxOJywLhj0QlRYhCLFAjZSG9eS+4ZVV/RlGZCqe7e1cL50V+J
4VrPFmFA9QR5A+FqQE0aU3rGMUiE3ifBenma9aLVVtE5VL2OhWl46gQfA4oKv4U4hQaZmpQBFlDE
IvqgEP+GS05x83cAGQiTSeO25MXJEZsRupesh9p2x7nkhzn2w8u86B0QqBuI7Y4i8CVyFSIiWU14
uINI2HUvc0rplaE+zyH8gfoYwvdW4umryQQA7TYK9n+YMZJ4dcodijPEoNo4v29GNUKxZZ+PO8+F
4OSYiBa5FQxmK9TS5qV4lKAtBxB2NRtfuAHPA64xw6hewag9gcORGGn5W3qdq+P+ofBIWpOyTWO8
Co86iwUtuF+Yu2rrWEQCxZGyw9SfAufbbX03R73ipVtUSJUAxYHSiB2Vg+o+ObwlRQFse6oJTpNN
RD2wh4AtjMjPbDAak5Qlx454jM2c44MFPVi6jvT68d2UO1lyaJLSmxlsqMvSMwMOgqzu10Zf4gGm
UxEUXT2qIQxTnfUZ6yrq29gLZVIpFnRkAkCmojYZ7dL6dB2wS39DDkIdF8awF/wE4MFXbRnEon+c
uND2l4ScMcxCJTEPvbb8VCr04FR6FqRSsssxBipcYTH/yjIPu3vOvgholDa/IM1b16Cn2FxLeCuN
sqOKBOyJf2hTOPUDdsLSOSnp/7au4Mg5p+dtzHskTvpgDVnDvkcqgr16OqCY0EXHkOgSSejdBta+
qMmXchZRYIhswcyjVfsd7Qwho+x2ec1SJsp4e32vgJasoAnB1z8Kf3IHfuuWtQszlmjzJ/Bbk4Xi
U7zByE+jXCsP4Fwz2jaNnel23YyJ3xlYttIQ3UkXNPv9agUHihi/Fjfnb7Eb+WhGQGdWRjRglRHp
KyeXRPd6x/swislfYsOGlyIfbhlV0jxv9YzmfkgEAlHO++mTn9XBrODOVKOyEoMT8ETafl/Akl6w
TS8yoz13OWDMHEsmsAoxAQPZ/TpcuZY7INbKOBp1tXercasjkNU6+RDAe2y8HZfp3CaBSxtxFEBZ
xEGUwQ8u38/8RUuMSfdBJlAD9z+yunecEEDmRXFZKDbCkeSddGMAmqm5Cmqj1qa6euLtkAVXm2wL
M06+Ftx9JnOYZO5G35NEYu1pcPHm26YWazdwnfBxH3FNBIR7Hurvw875tPT9dgfyQ3wZ3JWg6FS4
kycK20fmptwx7PL7UjkAhZY+fx6zrbdd66/dSqi1EjfvpySlrxqYk8QVPCMEWGkYGaGPl2XPqNyq
SxnMWtbEm2RlUs57olbrCBG7NobZU/6qnR5aLOec7SDcyl1sKj58P5UJj+sofB+DxoIC1d2ySXAU
kMBjjKUNLwZJCFEIcLH9arLf4COG9hnupdA3EpVE1sOnbo2zeIcM/xgCM3LTzwRgYm9OAfHhcKQS
9s8QDR9ilprsZTIXYVatoiLhJI436Gr97QVP9pUOKWhRjd3t/tQM6D7FpGRyVgIPgmfgKsrfwwyX
UXVwSUmjnGTN3WFf6OEHCK9iCZ04SXrgO/igPypwFygx0qvaTQcda7y2zCSXcu6CiDl3X74+45kJ
+36syPWNjY1J15J2gdSD/fJqqUkcVvdzIl04refYuiAQAt/gEusxzGdBwCCwmK0I4jA2FPeVINxA
zahRkhvlbEMcIOZgHUxFkytoVmF9SI4HvvFzSbuR/CnIW/aFvvn8fTRhqvARebk3dGz+Zu50U0LB
4KuJszPBQCXBzgLGpZq4gk8bbqvRnmbZ72R4ZoyvDWb5nEXONk1cpWSNxrwHjeJ6iVSpq9AmoibG
keKaR1mmOJwoynVXMaiACIwSDwKZNRzS677wMA+fNW0QXAo72oa66VBW8nOK8ScmEqPRnDjaxptM
RdCvaSiUY5M1oaNfgWG9CxsZI2lQNi9B/+Ol2iHPlj2S6VMdbUgS18i8fz9Ad1Tr6yeYlBI74x6B
jECwXkaQ9Ohp2LONBHmWWKihNX2hWFYyv1cfJ9LQbJFG/75bVgCCAnYZocfr63hooPqPzU0WzyJ9
kykUT+8lKGYptKjvsOeNtxoNQwb1QcGsE1NlmThp6TB+7lIUjf9Z0+Y59M9aFbyfoEIvs2k/nir3
X7FOxmv4IZtF+GUJe4kSkgAmc99Di2Fyw8Nj1OC3CjUP+6SByS0lp5pfr5Po9hvHefhbhfPRCqzb
HK6jLogqDaBkKjdWPMNfeXJ7ihRCGYLdFWW+YJaeO24dpL/jmQ2IzpIFK/KkhkD1dm0TiAZ1UJXd
ZtQOzMAGiMjTqxNz1YN7zzIJfJiL0wnk3KvbV0IUdw6UKE/EmayVIcNGipSs4zKfIVuIUggcw7Xx
zjc75uBjzh38kZ8Jry51dkhhwRvwQQAEDojouyI4YftP2vED9KMrN0vtFxL5hDhPjMM9WvqoOrDg
J9IiuY6Tmc4nietmTjXVcvJWbUTUZp9f9YmLcmOUZbu3w6K2C/Jt6VFfICmVti9YyMEZw7ULahwz
k4P/4wrpBGE9loAaNeXcxWf0g/ZTwGbZzVJDnDkLX9HjutNpk45oDJ71gTBgX+MOSOsho+vuB5an
GvOXgGUGPEpZ9FFIzXmFkYOVv4I7QC/7LXGJwoMzlDmehowwWgpRsUVG/ohOgHzsShayODdDXHp4
TxfdKNZj+pTNSYFEh5Znn4BBEdJnr4H1lcz+KmovCp/R6qqqRWhUKS5ki+4LrYRPXZ6AZ2vkquGS
snleGk4ZvHkMsfvU2D0AewHpBRiHfcaE/qk/I2KoGKqauqdXd2bWfklTdhSXBjgsYOvBiJnZPhj8
2TuLBJwm57WulIWDmYFiketT3EQsTYRMI4l2JlUBV4xu5xKqTStNgSPcfIE2rcraVJomqq6Sy6n5
tOuKox88dxS/xrkwkVMR1ikQ4LqimygDJEKj2y4wV3izS23aYnaaA5tMM9WDCN0rOqD3O7KZau9e
5ia+UNBmISwACQPj25zfAQUhQ4h8dVzMS08CAEcbkg9UIcjU481N3IAra/Fjn+Atk2FSBWvYiNqH
f9WD9mP/21XNsyEAYaPikL9BntPKdG+JduF2MZOlqys2Q6vUEZ9hV97VlI1Ekqt6qiZXgI/W3uPA
ieqNG8/0Xd2Kx4uXNrg1bnGjVl2B/oL2I6M6C/pzzV7WXn9cMAW3Ma2qCqvAH1+lSjlF77A7vQZ9
XNgvPfI6/SsL0r9ZZoM7KFAJGX7COp09SGpu7WMShJGBumYm/oR5rAe1bVUPWRjOi4oPEwm0l7qX
G/phXA7GcD9KKvUFUYC7MWP5C2Fn/KUggC91bYazz/aCNeVGVaidbK2Bax3bjaiIUf5v1XgolOCT
qYgVYU8zlN/jbomR17kt6nw4JFnhZdY7QKTQrfS3UhPrlU6IOXuNjNTMwJSJ/1TVknFh2KC+o0CO
8SDrUhq3TrU4+nPYffAPGHPoUXkv3x/4PD7V3VAUIPU6AxjBqRpIbVmQ+ZrDuEL4zwXJsd0r8/4R
ot9ImLqEgQBfBUQZ27azZUYNDT2A943JkQFUd1lerJSK9+YeuhwZNsa39sSGWRW4dk3iXsYptapJ
xNCBFuG85ilbmh9Qu5o5H7CwnnV22UQ2pC0++7rWwV+GAkq8+nvjCxQTVsiG+QW3fmLm2T/cX0rr
yqXiSrq8yRWrWoXuP8kquLWC7EiFuQKLbP+h2/nALx3W9QdnDcyoc4HFN8uC8bWA00D3oqCMdXia
TnfWwmA47k5IEgKe1/zbkR8aXDVWnPnjLJnjNeJ/t4+wrisf4eA6DXnqejIthYw6OSblvMhSMMlm
BLfOkWNyNKNDDbWbDPd1Ov4Mb/dCYU/mBWQywpulscg0EeUN5GEJPQFE6+whfprbkt7flNvA5wsm
mu7PsRQV2JzXBiW1I/C0Unv1NheQyFSFb8YUTsroQ9+ScHaSVqQukvGi/tmMUq9RDa6e4fa9H5gP
wwDM8kK2mAy+iWEoEVTtXRVObo644KAWz8olB4BaTpm5apRKajpl/xvfTZahjgC9UPeDN8XwFiX7
BPHkbtp+GbobJNuf0BmuUk5gHn+d5mKhp2R7k6imh63U9q01tUyolg8+mWjGvhITWPaBn0JVn2Kq
JLfruro+r9dO82gN7u+slkYphze/aPaLujV/fY2ukcrEnFCbW2oxdaI+qcnsTwyagWp1fhYeQkwX
S5AL6HfbY/Z4Xp89t1qVso8ozawhaBB6488DT2wGVzJ76lBSKnPEDREe9ORIEd6mMbybh8GE3tKY
L8YTFmQBZ4acWtYLilQ5RvNAhyh9JlpHaWk3TDN/mpCZVGcnSCKQy/VJc0CTr1XldCUychZ6WUSG
0AL6svyae1sltg1Vx3c0fUE2YBN2sv3zqdA5Rx80lc5c90TnaZdysMJ14KWZLBuI/E5HDHxtDnPe
kGl3z+hDG0UOvpYZYg4tGj7ghZO7WwiwkDcR2PlCX/sQ7lYjp1S9CCXbQCWSuEgKCDERKJW1PRtM
qbQe7S4CJSzRY62iD3H54Kxpxz+RMoiR/ph9t3gLLmGZA5vP69e2wwm4CFNtCRpa4kwykNjJ6ry4
DUorx8JsuumoouQR4KYS9IxNLWyqXl1SJ0cXQQKhEhJQak8T5JIuf3FDePdRCe3jJ4MwaArykpVk
d8R5cY9mbxMZsxga+pCUOq3pwgFd+7nX3jcL5Lm3JJPwhvUdbp4/bMpCGkENJUMyWZflI2IBNUlP
7lBZgCsetb5sGwl4h9kMh0u9A7GIhyGfQ4ApYyiRl4w45AnL8z0hxm53v0WMlm0Xxc4cLecc3R94
/I/Dxx6iDji8OW7A0GsVDtD/bf8JHBHKPPLqPjZGPJoHZc1fMwhbO5OhcXcTh0AOFlCqXQS8mynX
7FxWb5QFffQWbDxNQ9cOQEgJ6BB9Y+tchx0BAopUFXOwO2paob3X1OaongnAD4pJv/vl6ldKQIlF
t3/m26HrYoTlq7osMYz4K7tBc43naopvFgfX73nTFOZOi5cc6fWUWQJzpDQIskRf6TrF7eWqjzl8
3gtYVuNJWLDut8eJHa498w9Ehl30IZVviDYkqtQ/eONXzw4s3ZC5N/P1U1eodZgoAneH0nwX+rRq
BopfOdIXdqgBh4eZ5nWx0DFZ8Cdxvpt8qrWNiBIV0TZ8/T3B5nfQ5XH8WrJkjw8KjAb4yVRE6h5d
crCIfsqxXVo7TRSA04Nn609l6BCFeqrnZ/wj9G5X1zKxNVEFOo8lAkz+UsZscP/g7oUY/5AFkBgo
TrcD40cCgZGQe6zC/dVdZ+XmkUgpGXj2Heo0nRwO392YqvR18Jp4YD4FPu2abTdRlyFPMr+cB4kf
DhFPAvD4kNVlJbzZCzq7hHwFv+uNozwrsgM2SOBo0C8gJSLSvJt5Py1zNnuA9e9dEgTlGrWlHXQv
jS7EfAUZdDLIBgpAUR1QYVvJrp/CHpSiPW1cW64ew/9q7myf6iHU3HzOURrYNj6MrOp9r4KQ9/s/
6/JEvI2NNGYkVA0cxMPSAJYRqPjbMztXeyrqAP50N7TtXGGSeQ+00S4rIjJfz3a5D5O2Iu9Pdrt6
Aa2Q/Os+LsqihpFgmff15Yla65Y64gcNy4yoV0wf6TLNvT+eqJGw2y2flJLx2UF8ldI2YC+IW49M
Mnx689VNSADd4knzCyYsEogdNE7MqfIVBvT87kEPhnpTqeVZQeLhZjozSbcYQV6inStVVt4c3bCF
jOgjkg/2vhgRieQJyqNzUCMyJx2+zwR/sg9PS/Oxka4sQY6mMKBJCm0U3XhgtU/w1FTbfORbDczm
60Lhot/RcChiL4qxvQpEna6G7vc6RkoVBgLemaL+Jy3GZtC2r4UCz8bXg0UWeszSLy6SUe1rDc7q
XRlXA1UxlD4D7da2qNxf0OTlLE2OljSdEjOro2xZrsi5YsVHtFRDPTGaJmmOo0svWk4QngkEaE3b
aBsoKVhz14veRDEZnDVN/wD6pbrsmFkw9i+H2QFJpYDLJqBsKsy+124NnUomq43T6U+7qlqD+88n
OyQ31thqqVL5dKNJSPo0oIuQ/7/LMZOJsahbaQSwYTqaEcSeRm609H89pvdKAMvMx8/1qC5ljrRy
uIS1dcLD/6p8rHDKqP9gNWH6h9K4MU3Gjrnba5zJzgKnGc1rmR3gqL2a1gE/N08FfT627LURpL/S
kE3jSKCEe6lsdkOqtpPgSpoBR3itk3rbzDDrSBHNMYgI02Jf9I535vJXMaGdiMdYlbdSeOYDVORU
mXzwT+hcTWLfUSk/KQlCTPbJEDNBPosKdRZIdN4mRdnLwKPYird1hue1djbfWl4PkZZ2SyIXZZDf
uBm77MGcWEnPxQYyWCkcjqJVm6Px7rVX2dU42vezYcF7hlFzjtJB4/bKw6ucYajtuXFPwYqMy6J9
Y2r6e+OHpdcvpcSe2sW1v2PFxDF2SpObw3234vP1Ul/grUOjEZn9Z44UJk1vqky2EWQhurjOHVKd
39SBT+By3RTq69fRQBqKZy8rUYkuC68i3EItcEyqAfvyRWbGVz0tngBxVqvG3UpgeaLqd/j+HsQg
s0+Ogvzd4RpNYpDVIlFeZ/125lHK3ZxnczwqhkI1mKTtp7l4FgTPkkbMgmmBltvjG2bJzpk52en9
JbHej5nvtiId7I++0QRmEYVlV6ov3WNpav4iPk+UcP2FVIdmQ/3WTn+I4UwrpYlQkq8CnZgLRx8u
/il5Afm8hVjIHiaJGUxzmpkwuEmiQvspq5a+kYuv8VSaUmXpm6WvqWsQbZLGvzrQM6NJgSxvWOLr
m5Xhku1Onu95DhNReCiBFtWqm0Z8Nz2glp6ANjklhg6DhDlOaPmsh9ntGQW7v5vu5T5jBlRwuqNa
e74MPdK4Z81KN/X/kinvSNLkVcmtWqyRgYkLdzZ8+EI2c+9cj4YyN8/ss4gTEoiMIiGDmjqIrYon
2QV6lY7IiD1f+zuFm4EcMtX4O7nNGMyhArrFakmyWqx5uOcj1K9pMWfPQZe4NZlCUrvAk12H3TaB
ZzAjkwJcnh1AHP3UYY2QP5THoiGO4SSW0la8rJrgh92Hq3dlM7/JS4Z6r3bdqfkfTxv5ij6+OKo1
y8xOULJKTo8lYZ7di4L4sC8qOv8BLleUO7TkmDGrb+9b8q3DZmwyO10w+CdFPyejeQbosD4eg4Ri
8k7XjYSShghf9Vi3suThbN3fJWW5TTcPb0G9rsOmUQdtx8N02/0XzrQF7EQF3z+OKy5anSZWeXRW
xtbJna2AIyObH2IXMbe1dIdaNuzdp/7eC4Dl6B6+fSQkAsvDxytdfKKeOHodWUTSPINzj3AcVGIM
5nc9ijE98WXZ2PAuLtv8kQUjLabuTd0Bm9RkwyYnjGyAtSXZrfWWrQ761//iS/cD1vs7WrfyHSY0
GyDAgkL8hdV6H+QQSLUIHN5qKclSa1Mmn1xJ9MNMVD/fmOg6r7i+sfdGWh3GRz8GVmoE4A4e3SPt
WL1trGshjMeTnqqWftomSZhAyLx0/EMwkQkJ6mK0lUiNUl9iM9IFrKxJ4mvZbkVPeVj1hYqBXQJo
KSLFM68WKODQOLnPAtDkuoiQdANKX1Rp4ZCuqc+zPkOZaa4BUJRlCq2rajuw8FIDH50g9v1/Kue/
/klsCQhHOWy+jpGCiarDrTQj6MbVv572+rx9qzSBvoH2NaYkHo8JQVUNjm2nCmXUe8gFmTm8uKW4
+54T/U8ORBnKtS5W0U/eyExe3jaYqSF+NuQSyUhiC5RCEIaZnZFFLqDaO6EazA0+53HM0H3WQ4iK
Jr5T7dDzy54gVBfIAaveym5M23pgYk/tMuloUy3QCrEu7RdwpkT7u30943TUrYzW4Iqb75arIHsM
WaiNHUYLxt+9u500HERx6z44coEMiNcdHJZ24FFBdXb1lk06EofYv/XYqJ6QCDf5hmxogNZqepHM
FxBO9AySEqxSlE42hEWiz44tSYoAIbwDlcLDtAz0jxSn6RK7QL3WcuQmOAnJaxmARQHZNuSJJkol
1Ojwa810UDwXt8/bdJ3F4SWr+JZq73/iueNqvwZEYdH2rJ2RXjqUzVxe/28jYlw7nPRBz/jcDkRU
++l5TBcACG1R2GGyTE1iq/pot+ev1aDzJ8zuU77RjqIxn475wCRshKUI2k3W1JyJilgHPKG9S9Aa
CKivmprC0DZKibrFgYyES5hNiMQRqfk8HOKrY/V5ZIYVUW3sLeJ+HyPUxmo4cn6sjqDZXEz8wAr3
thS7glXe/u/DwoPjTLI44yGTJMbnHEsW7/PSHZoCakPZWoLE3W92brGLiXH2LGmKX9Q/R5UFeqZ7
sha132sg5j2E+3E6j+C6X1A9DCQ+A8BWj8SSGR/W2w1qrqDF7XLdpd3uOeVC8ecHiWWBMD72YcFd
sotMg54cVXKLLJ2lqNcdkuJRF3YHOS94gc1HsLtD/Yxc3yhZ78gMZVtUABe+cj6xO6W8hJwi7Cqg
6G5RqrDVQhJL7lGGSyg7ZBel/OFM2suq1p68cs6ndzfmke2kxj8dHD9DyUISsrU5QMQ5wjDeSTo/
s+B5+sZq7DVS4jj+M5d2WHBE6wFvlHmDSzdWWdO+G2TLi9GT1aqnp+Dc4BST9a9ybW1pzEzk+nNQ
4XdDP09Oh3hl7GxoPalIqdxxMocZgN2cdWW9fHI5KZ3RWvURyMugbIrOooCh99XRyx8AcfZbQpoj
sGuzAiw23qlwWKfxvZ3JBwdPWd8v22QGqyclBgB2Q7ppqpIH2pHAeYCj/OpTRI2sxIxWi/ZhErHg
qGBr8hrHXq1/6mkeBOW2L1nUlZDEpsyXRjW/T2atKXwTsSLiDR6mf9i/HmRdw27R+/pJOlo/3UMC
4Bq+xfG0Hljd2e7i3B/JkjVk81l9DjGZ9Yo2+5IunHZyH88ke3wPTNvqJezz/M65waw6XDxRIUnl
Wgcmvr3Y2KDqMJYiKtawTTRs//5p33q6QQaKDZ2oqBXfeG8ZwVMkMpGG0J6QyWXBx3FnAky/WG60
n2Kj/FOxLcArmyQ3h4IT1NYIkmkILz8FFInbU5V7QCiKVaOtfQntttDnM30TVBFwsVoco63flgGR
oVxLuzOIFTwxq7Viypud4K2c9tbM66komM2AJx9TQeREqvQkPw0WDwIVXhjrwTtwjxkjxpkLhvwQ
eGNexDzSP+SCJwa/WsPmwY5Sc/rzrfIpZro1HlcqZ0P4b2NlJtGA7g5xojFYu3O8Tr+bXpnhPCWt
iuXqVlUUwgFIyII5KGzOjJGcLAreHGLDr/qCesUab2ClPYKZybh3iSpUMgTS3d5wER2EAi5gXG7u
Lf6U1YLfrSS3AH3V8sc849CSUaI7/19U+hbaUMufedAzhhj+Uq3BvTL77kQFyU+yLLBTpBkVOGLE
/XK8Bd/Lx29xna4TwIIIG1DZ+efQm51gy0uGZJ9SsrCBhneLMwxaEsBtdfTZq3897SnrsJsXEc3Z
kzdElslwL5e03wNZbPewgDCPP1QyjrZwbrLt+8YQwi6/rbECWO8mzv+u5TUzKa8owe78xDnwUfZp
0jLhd7PBisPFivjsoekg6QwK2QUVDfnNeqEtW+JAHcZM02aR1JCtGw0iBLvuGSuJZgJeYAmsarPw
DTTRgjGziFttQ6Yl5KGVECunW9qMXb7jS9TZVVuvrLIVEuew3tk5Y57cw5e+dEqAr1/YIsWPDVQV
jZjNn/XMiHMT3FdCnMWoFXxu/X8ImiYhUdBoUeHx4RSIxY3wJtWBu2OQW+qvyrPlsALtktG1C0EX
CWMs0EV+FGGZcDej+G8J6u8aAerQfDEKiTBs9l0MNCu1KZZyKl+vw1igD/NEJjAFzuIS6S7I1Rba
aKjHUQ+0s1DyV6OucJQFvHcB9txWxOo3D4GS1FnrVy8WBR/dtiAylAL8yZe1d0SZS22dG35icdqf
EC6rLlxLrq3V3PY7Z8BzhfxPNbWrTv2qYgZAmu9utpq9zowK2YOPTiKCT6jwF2qnlxySxFab0AEs
TC9gRoJmAW3Zqe+Ec2q1i84YSvRXgqQ5OZnrUCOyUbWB8ykUbfsxEycm9d8W0LPJnruvuoODCS66
eA/2K10Rh4AnseVafr3NrvHuLX0HrSMtPviiADeojntEtsFf/kLHeKEOAYE0XJXO/tzWq3Hz7pzp
VtEpMs5kI4K9Hkap7COTwqoXXkp6hoi3NHrtbY7EaZ8cXDmkN3x7tm3AVXSPZ5P2gJPeSxzt7CZE
UrQOssG8KvuUfjEZLRshQZ6zPVksKuUn+/v02jenskHMliEmP8nUrglCl0L/IXAtyJjwGEfT83AT
fpFEmwMLAC4bGz41PWjN28a3mViY/WV84vJTYKs7efYi3KfSYD2ylrKQgLgGALhA1Illm5oc9wb8
O31FTB6IryQPTwWcPghbGIE4JPZzgndlCyq38ffTGlIF2bCAf7e4ylKYxf0JNruKprr+7kQrxn4D
2lygb6pefn1d8s8mpS0wES2fUixyqKbTdr4BK0MRtIm9haMr8lsTjKcIKFgiAZw23a/VbT3okKZS
aay07rQTBAdNp1VWxXAruVtTHVR5wrH47fCCL9k3inHI+aqRukZeWwEImiArmiyIGdH3XE4sPSRk
Ws5gHR3Vadji8dG96K7jmKu9gyEIr4rffw4qNkA7kMvRUEv7MESzjxX7eB7NTrA1hyXDcPNOeudp
DSpRjuX1AYOrOF3rq6Wl1mV1ISZFds9hm6BaQilDdp6xOuAdyE1yx6MlmxmO49c0V9chyMvRozqW
cOsl5LCMGnnnV6gjfBxI4QyqNewIvtEo1ft57fe6UoM4dFJdOBL9D1rSPfyZjbIW5DyOctztX5aL
hvd0Wxch1GY6eOFs/zunh9fIiglPItM4SAzTa3HGtBkWBJZhJ9G8kTP1N/4Weg7/6neaUHIivsIt
2+COVMriA1BjydFpzkyGd1vrC0vs6h8Nn/0v3Pw+aVnE9Lvkm5JK/g8qrjMwlZkA+5wmj3haPBOe
0FJZiLb2wKgMuY52EuTKWR9jvNtAI8V7c0hnsjv43fj6uJd6RE/6OHiYPyju34cS2RBuTCUkhkXT
FyftlQaJYEkCNbW0CU5awdZ+OOh2eQq12/z4s2IaCJWN3aBaU4VoV9xSGnT8o4tJvN88e9RKsEBq
0684aAPPlkRZBrVbMc9cbeqhXf3Eqvc0NlJV9qK/s8ZBDpjqA7PQpp/ny/eEL1f/xITYHSB3JtYK
17xJEU1Rz1+kGRxHr6xintKgD/uIzF8WqBvCeFsfVTEdMCU6Q/jxPKd9RIVP1D8IGNde3AfcrQqA
nVQnYWBRYlKWVBd049dFCoo7gjb4r/z5Q/Y2wrQD2F48HztSx0VyQeTlXZyAnXOBYAEaIjgdWcsC
tc5TXK3unETU0s7I7j4CWIH8v0GNTDkma2XDSuxNeQJiYJ1Pj4pVDisSzup1KPPfqpQiDpO5mfTd
Hp346md8RTbEwtPSV1qBuYlpQHHON9q6YrqcqPxK1Ld+pQY7XJpuxFhyvNnEZnVm/C2jUjliJg33
yIvmuAkWOLiSfeEF/R8PFAmVpaJKOyFXez/ri59tF89g1WeWge0RVjQyxOwnIy0gGPB5wfa2/AbJ
tjzgdxUcIbqUbWhgjxHA1nlsduxDiq71ocWp+ygf9qcnf8RFExg/lSH0ZhnDzp9Kpjtr0cY8lqb6
bXDbwjl8C2/U76NbRNCMlMPCYaKpd+FFJN8lC1LWndoala2jq5T++PbYgJEV/+BgvVfN8lbMOtu3
JhL0lG+/Y/EvCwCJTg91hFgsNNtBfsvYvhTVq0DZBmgRJZmcoA9HcsnLMhXgnxYtnNZRfC2o+5BJ
4jT6pyweOuHCDJPtzcKMXs6nhAlYAmTsBvIaXexxkGGR/os8H7JhT7IuBWMr1DiPjD32YKqcH9TH
x5WJZw7RC9TYDlJPTddRD4ILHIz89LzFrFfTfgXHJInxnA+9YMTZBL0ZqLVYp6RRYStVow96lmBd
w+Is40wShleF0NQQaewC22pHfvWo7XRrZ17ltmVxKBsaQu96wQ25Q7YUkkZlqiOTCEL0EdN6LN0Z
qYENTAdkpXs3PWX78IcgOvZW45BS7gXeaOUHZ3r1PRtjJrBKKI/MZv33aQHZAXiqOMroI1M9zQv0
jNWfbuBH7Ep2ctX9m/98tHK5O90xVr6kTvzYJlcpYzXLz7Bcok8zbGkljfLguGs57Rdu8vhdeqNh
mZG9OxTs/XkJpETKD1KUpelD8zXLfDz2hl5Qgb+p4EbWSL22Sa9RL5F1abQ43cfYy8/SBSrfUUdH
jPia/yGZ6IWE/IFHveYWk7o2IkDk34ZW9ATc6PUhRWvKNJMSNwofPj9zbnAn+1FQFLgC5LnpuAQs
9ilXMtmNz8ec7Tav0tx4Jiit4k/yEgX6PmDdsjGthYgc88CV3Z8u0KZy1LJwwVL+sasnE2u8RPcZ
c2uQXL/cxcvfuCvOQ67J4QRQLyl0cPEunoC1XWf7sw9rF+TGXOJS7oiFWs8XIlJcJ01YGdTxTl8m
hTiyueV7gukGRWWn/CK4hTV5JGd0EhOL0JeYb7Za7+jJcgO9HtRE3So4PuuAQXx9vKKwZxvmTOky
PaHna1clqz1CQrX6ivitIjf8A0Ahgl5tDlU3boROV42+GlLu9jYJ7LmdyQlxyNfEzwRP07qxja+C
pt8uwHU7IarYpA0i3lkPPfBvLtJD/TgjMpqyZun8b9EWBIUv7SaTUATAduWJ2OwtkJ4h9T0p5jvb
SJxGiPI9JgPz4Mj3oTUUJJVzOoRw0FrP/06Gu3mlDy4gKQ7cZemdR+muB/V8nQ7AS4VbpOaZNnx5
1QNYH83PBcr0d4J0NeILVNUZnutKFmw/jKMwmXeywl0Oc/ONy98Wv24tvF0jTJT7pzgTek7PmuI3
t+G9Dqr5y0jZ1I4xdCzz9sLt3SWCwT23rWGY4++61qEjUrLXn/UCHyn0U7BHvZ6GdEy0CodpXBWD
YrjeAUPkmYS8xeWVorc6NUQHbgGKAWLXkMztAVqRhPCQqDFNQwwj4gdHHT8s+2UK/9/d55xq3abF
8eVmaS8WFWX3Ar/qMr2psM2q5rduxdSV4n2gUksFa07RfVsPZNQkU5gbVbHIWys+H7DUm+Ne1bDS
lHk2WAyM/+2Y9FG4oz2f0o0dpCRDcvXV+t+Cf1FqNpIlvv2Paazby6wQjaYuRXlGTBP/AlOc2j5+
jq+ZuQwrY2FfJTTe19E/EooLaGa7jlI2urUClh0mUWTqe4c8+BsEGPzQ5mwtkXVxsLW5373Oh2M2
6uECfHk0amQwcvoqMMKQeXTbmJU5uwoRMXlp9x//JbHLT1cYBeU/YZ/MwkLbvrKc04Mv0RAoDxhI
jZv3QOC8tgJq34ZfydvgD27vYFGwclQH9R+eYFSb8w5A2sKwL/JpNUFEPBIerhIHHShofiIBzEe4
Uf+AiNn2UJOGlB9ybXMtH3pz0xM3AQ7c5aF5whz94ql66STduZXTtzGNgfWBoY9ZEFKyjELp8l3w
hylRdf2VAmududvXS79jrMpe86l9DR9jYdA4IAzxVw0omSVd2XNBa+11QpcE15tMMM+4Y1NswH6s
eGccQ+zwHajOj2HXjE9co27kHy0JJ0lnhp17lleOdrAj751VI7DG0yRQwjmlXdXhSqhR87bkFozP
D0Bv17hVHmKuKEPnAvVeiDDxRKu4+PJ0i+gtB0ldQcnsXnMPW0Z4cy6KioIJNlookIN5naXZOzTB
MTwgScpbxYhMnTQIUY7u3B47vQ2yNM+i2Fmsgv1PV6CWgu5WIwli0qXnclecv4iudAo/806vTYAf
OYYwKsb++hFp0xAO+NMDdRma4UT7rskYt7BpCtG9equHWIKKVxUlv61jZlktm3dJag+SaWmPA3TO
B6K+l7JwUSqX3CBzGSlnA/8d5+2OJIGtCf55TVM6K9U9RRLYrqTz3cprPCAbBmeADhEBUP6bNxpJ
50oBBbEkI/ufgHjsqUqloA5qBBWY8n2L+1kpuQUaLYtalC8vZ+KCFceRxjOkB4gs473VQ8m0yD19
0eNjgpnow+BGqmHwbHnywvcCXJBOP8dLVnwU/lOpLhS+NyQPkJdzyYayXZojm3rK4QsipgUEuWWK
FkGkGoxqiMSzjybjV1GHVP2x12UUCaIGgrNe4y9lBI8DO60wlZxRoRieI6/1Il3JuYsQgLjKzxUT
F13YxTxtHQZK/Zqh2QOAagEGeBntV3GK2fE0Bu9FoakdpyEBvq0jkrxOJrabuNLd1voDcrHhGZOk
cnQiCyq0+dM/fgBmKUbFaWJKNfv4LwkRKnfK5RBrH/kDBfLBk2fxvBBUco4CZLbPyxCpTdirkUVQ
kNu0TphHpjYzZnSZbiKQHESOTsdeS/NuAatktKimtlTskrzCt44mKZoX8tXrMJTXWAVLnAM4ptIq
1ceJua7B+YjBSDuQYpU/n+aDzooYs3x4PH/Ayug+6fvnIOEeCoTpYalAn91ORQgUhqrMK1FU1wV3
5iZ+lEglbotTsQFtRw04Qi9rK1yWM7KTuf61E5QPFq1/ICiU6EEHkgxmi/AWTlobGGCiz1Pd26rf
zevrwWg0e0RSG600K7Vr0X5FVn10n20f51Yd9H3Ke7jMmZwfK/XSC5DNjhTRHM+g8oVw9+9WSxaz
w3bRFBAf4K/2JhDY+Wqa1sKrS0mgDcZaJHvVZgQyn9xhXS9Vp/emTNqvnT5ivtGu+N7+WAvaGDd4
Zvj6nhH4NO1rs7JbeBpPQvuiTud2m7gyEA2TAMi8BWrSLFbz2iBpFYTG7lIDgg2+7R8OXN66bO0l
RXG786pwDX7UidlmEhjT1Xkln0YVCwM5iYHnR+6l0wCghkwA7wZdnLnpjrXHYtStYMgqbfSn4P3x
BUrNurWAY6cT4fsjb+FLuC7igKL0Jz6+8ULP2zqhhoSBb8urO0aUnDrPLQrSv4+KspHQPmo/c+Z+
NI6QVghZZzUw5mlyUomfFkC7p6yBvQgyadbaoudFCvLcJKzy2V4Z7/BAysVVFw8XU6C9rCRqnxrW
n8JBsWdYaIzGPAtc26lGkY98Gk4Ti46swV6U5qkCByKHP+T8QmVjGAd4Ye9MOTCLlI3Uk9O7T8nb
sNw4l0SFrzx/ge5AbdaZiEkckNs9i5z8rYHLan3mamFugMFI/gKB9MbzJssi4AU/9962jTPpyGeS
mUQ3qJDrPR++q6/9xWzm12nM/d4LxbWohG5H+vd4J64+c34NSAhSJIgi0YoarqnJeoUay9ChzTLu
7XBYxaEIg58DXvusTZZa7V6r4aJ916msvxZsdAkL1fChqUoVghRPBHhcU0iUm7j4jMMiOt6PkKDq
lsj5s1zoIpxUHCicrWFhQMts8+PiD/MGQUhekO9XFmakWgTLV/yi935pzTHh2gsVhKT/NZGB8VU+
CkpdmyNYU/lywMAapNDHZQ8tiVbpH7ZZmbLa1xyNmIDvwyYEO+7TbAVaj0U0ij5joyAAu/6Cvfmx
b3FH68TaTLwtWQ/X5qBXWwSNXWYcHk2DFS4+m4oNk8oF/Y86ugDu7u2dsilb5qCW4VY521qgi+/W
wUxAN63NwsW1BGCKa9z8q9AWyww9aNNbELs+XYwVd54GoAs7duDpCOECRWPQ/3kR851q+HR9a1AX
oJAY774iP6+4zCwtsKtuXuIVd2hTBOmuRUa6qu2OJR/eBK2/fOEtYGHe9ivuZYYOK3DzUvu8qwhs
Ts/dsdc0HPPaGGJWoDlfLkT3UC2DH8rrz6ieEVZf0AM4j7yRzR99ZIqvKaztfgznrLW0XzqZrVpg
ufq+mXFz0I6qShqQXb71aQ0vJk19V9/SGqdmz3l1XUrKagl2jRF0BIuRzkDt9DEjWne9jgXlNzrk
OOB89QRDHUmbH6HWUjJthC1H5l64OSX3FtoT5SRaGMRlfgjMcZmWYI3aOgjGFo4xWVPo/j3jDRvB
M7hVHhVhQ3/R7W+a1NnvHQohP81XIf0kTwRhLxGrQX7BWgcCUqVo2zWANlHQHmdSfgY027jo3hGL
394VOZRS8mRvug2dNJADIqDwmIliL07vi7vvpL3uReXfTquT/TVkqNlsB04Dm5BLqFI5uWDFGXDU
ELn/XvQlu+ZZ2cyuIFxHvHnHdRU5VVdjk58Fz5RsRax68i/moZvYGjjz0k6TABTHu7lkz1fkr3OJ
55feQYisQREQaT6XCTYfFOk7mZL4G/C6JIaKgmsFs3Dls67sS35h0Am6HERteZhrKNPK8KiekzUX
djd7nXCf3X7d1+/JTlCTGnnEeJT3kAbcTM3AgsvA9d+ScGSk/+mxyTKW8OZPtJSSyAIV0L1B93uF
U9huvYEc2B9tcmdoSDHKR9EzhFAiwpW7kVDMaPsPFAXGvCLhmUuSOk36+pDxZ6dWsFJzK7aQ8kGj
wL3I5Dm4XHnqhngEwFfLFwksC3uHYefOxvFeZ96IB1dKmsIGHji47NT0l1Vyvp8ZFEZlZTdhNacJ
iB4WmqDz+JGhcG0ZH3ttS7ykiJ2WMFduDM4wwSnS9VjoqH4Z5iu2ZBYPOexTAp1Fs3zqkIoZ0WHo
4ubK0HKpyMP2jQna7GOuscQhcAa3G7tsSqbrm6nKyWg11ESGK9TSgeNI4zSfM6+Vv34Tv0hPf7qn
xrfNKCryLnWX4tHRgBWAfEDbGfXEAYV/HFDY0p+UEDLX5eK5e3ix2vvvDyyhilFrDkLsTBcfqy2H
u80Kg8ZbPmH8TpK0ybL4zd5ZsGd55+Pw9wY3GRxmvNw6toHv1Kv8kfP2mPL7f0Ebb5NTlCbkAcwH
o//9kag5wbkNq88co+dscu6T92hvJAqjjMfwvx9aqXTepYz3cZ41raD8VaSRUNBTcSbl5Dnz8Hax
g0/5kIldeNdAbsOz+J/nu69mtgyF/ltjaN2dETMj6JmcSYpGi0GCiLn58AbMvdOwi2VUINpA0epD
xwSjuXJBz6FpUO7LPPW/4op7rMSa0e0NDyvWmf4vy6eDKw1Vy7L9Qz+REHyu0eRu0OIf3c26Zfe7
FUwt8vXo82YgJoqccNJwArhUkwtZAhgEunVdQCHBet3/0xWA/ZNvXkFdptGb1Tcp44b1EMPWl5p7
+RM/Z3s3ss0qDaWAid0RViImgRmLNahMaEkHLfZmZqHReEGVATv6nPjL0EqNtUWJ4SdEDfLxcK26
/S2vDKDHVTqAcJJ2MryR4tpfWkea24ltnUHC4xZF8X+tEySCRLhnsMr7zaoDvARbAjl2pg8TcObH
mxCms5Ks9iUBbb/r47HsEmVGW+8bKd3pfkwtwb6Z4rb61SccsDwaxKrqtQvfO3Z5NDOlSAOW6U4a
jvaMm3JwjbOQATlyL5yG8fhSYcC80OO2ZETyGST3/JGje/hadRsbDx9QFCOwf/7NB4gusgNxZdSP
wDj8omsLVvugmH3F8k+Bi6vDso/zOnjRdWQKzUOAycEuEuoIcwAqIuz9imX2+wsznbsSaNEpy7Nl
Ved1QofnQiSca+WI7CU/nFK5C2d/8M9MJmqqKtPf990dU9vyzH+KrvrFxQgEFUgKjqPODWl79DyF
qCLhL3XZp18NWU50gyg/rFq92COkV6wl/KRqO1LwVE6yZBXMmO7Dzhb4C0pBrTMpcBO9qFzN+SIe
zTVmefsAU5HYy8bfRUq06b5TUzuLr5JnoNvtU05XywYtj6+OZ1tACpIQyJRnJIzkAuHalM6pLeGh
GQFT3r5xW0PybRFVcw2ik8X1TbpxQP6DdBXaVVlwUeJ2EePywVmt8f3a6EGjjmXibuUe+zefOHAo
UFFRdeXG5skH/T0btQh+rRWrTW6Kl1A4vhstz5BgHIu2NvLlafvZTOxROU3JNYpcDNNlRyD5mAGE
Dp/8utgKKb4t7L3uiyVLhqEPY2LgnypomaRpyRFzCpWO59NuYKnPAyfzKD2Vm2xTvm9wYJuwyJ0Z
9IP3pr+9l2aaQMUH+0IPAW4VQNCOB+Nvo5qH2+tGi290EpHAxqcA+hfrB0R1VKxr15o0452+zgUm
YbhaBh9r6mFDJ4/92OQTq8yeosKtR/XK9djfcwbjmFATf12pYXrh/JtKuQmFgU+8k+E7hmmLlo5d
VeRULcYv+QhtiORtoEk1HDjcZNrmmTFYXt9c/710/p+rmVKKrCEX2PhcD+61JuKQSXMLcl1evMfT
5nvbD0zQJHikqUDnh58/nwvFvm0BhEOY19RWFY33tWqkyWzdLBwxMn0wbw8dFl7CVk8eMQOpKJ/V
kD6PNfu6bMCDtC9SRItD4ThBqo2WzJarMfzJwpxltD+Yi12iUftXwwsWOSAFnUhsPGo8JpelxYb+
8JjBM5VHdHuZekRG8RMFJxHnLWmFc8tbpM5k8rIKYa8+f5vghA6yYCOAljxXQCrztwCyspsJ/qFx
/Vsjim1IHHyT3DJO8r8qC06uUTWLC4OCdBsUfpLQMa5LlcQDrb4ab1TW067iPq6lTxYHJFVMNeQL
PD/+4OXAMuxTphvxsFYJXfQ+29Wf3An5MfCVCN05v8qwXbtS+la/TfkKneXp3oN0nhm6oTJKOnU1
eUEXeGFt2S5AP2eJTofAHgvdoWCoNgvMUWm+qYg1pYJZBI2Op+OGAwUK0fTjYgmeuuW0pNDOjK7V
f6mwZtizXwHGBMmt8yMJ7uw628VswAHvlgKNDDMQxp6f31vqWTGaUI/FR3TqwLWvWeKbPzJvVVTH
OZwJ6zZ8AG7XMf2OmULjYjdGwYOk8McXMz0w5vQIF8DocbRvpK0F1kEZnF3cpBSHGqjH/mzMiZxC
UPJKvOFCZn2DthO497MnU+4cFnqXSggUOa0fsP2UgYh8cnn+lH3GSzh7JzBYlDfCdW0/123+upPz
cFCX9kAPKDs0CA4Wi9S4RwsN39WjPJyCorg5HikhSTTTO8+7AI9tteqvfKdfp1JHJzLuANQdhmOS
mRwwiDqfJFRuigjRSh37CLsMSsxWwNRm5oqThmu74illlbkJYaUCkeyzWDJAUHmqX3dP+pii51s7
0pAKuEeq8Ri4FgDenvl/yv3Q96lXdLmQC4Wxpsrv06KutvLyC1yV829Kntl3aiGDw3Q/zAgGDsW4
cj1tAcvdH4xo6aSOA3YSHE9ZUvhKOaexp6u3p+dicIQRZ1eaDGqk6W98qtvh/hkHkaLytvi9Nbev
PWI8dJ/GXwnuNkX3ze8Dp/S1YMXtNfZywwjnsIU0cuIYoabOw7OUmwW9JBOZMPKyHGA45/qPtFxL
xmZxwtw5EGrXE2YP/A0vfrfIHdSt8NR5mePuGcWJn7A6O3tBx7OFlVVGj5FuuWdy42aBqbZOz5b9
lON/rEIFVou4cYD3Y658z82CWv4l3gK0H2Iz9ABhcogRORjXq315xzpUspn0Aq+aRjhh3ZM6mXot
IA3NgIM7Msup5gdjhSu7/gl0fO7+7ys2IH1SVPgSJ0aaD/O+qhThv/F7nAKQgW9fl5FehRs3LX7O
CAOXUtAOUhMIPVsYXnSNH/h9Xru8qRPRKnuPSaQdGBrmvTeWO2cVAs2mhSUDo9Rk5/8TUFdcaWW1
d0lADogo4z50GMtUbR1S5/uh09l316SOOIrSgDgq7xy1ibfc7OPJovQxe/2pUYiKFq5Pg1mcXdXB
H1C9y9EzYT933qpTj12jneTb6Du5358Trha6LRqnvag4+yZV0wuH3tXTGoeznqsPCwv3ZY63qW5e
S5tBwwsiJRDA8htmKD0v+0p0m/JAik9zUGdFulsQfkCJ2c5kensuhPLfcE3oeRMhdAzpPJrrUhSz
W2qRnEX98z2qymW0Grqw4hae+/GQZ/XHIuuZJwDtxd01BJ3YSPRdof623pWefVk3GD8BqSmFWv5B
eDJFpDGpkMaGMqwI8ZSBLJwdbZqAmo6N9SjUabK41q6zLowRlogK69OUkhLjpT6DKNtTZ7oaIK0p
7yKlomsu494sC2ikZSTac48r6m+iYQlmie0mlHgR8h+52vf0fdfY5frIi9dr0FSpUFOll+CTYzjw
sZ5k2dhUUajYMDSfOUmhksv+RF5xbN7QZ8Du92j+hRFuvqZ35eD/3KmuOghSfp21bN0p9DLu8inr
WWsqTC9JMjN90eyR54jwvAtQqd07V8WXkYLgHXuofzCBPWSvIHcSPbNvSopLtg5EQ0hlqghksjTG
LZEbfNYAUjKyGbsncO/bJ5RtUJFU21nO2DBgG2GQplihN5JmepWkW9WofqUVCGdg8JW83jayLS9w
CJhPeQwjFeUqym0oiOppIIIebjQGXCmJEqevBREY6S0oFuROz802u5V3jsUoqykPD4Md3NZusPjL
KVne3w0QmSoiBHKFLHVkaOq5Je2BgYMh7Pj67tyf8ZRqFZeidWzZAbWTM9pfN45yx5bjZ5Cr2V9k
NhVQzQe50HmHdnqy8r08skR+loHuFzyUIYUKvv2JfLmZeiLeTU1rCIHCX9jPiOr3jrnQi0BKB6eY
ofIqa0Jqwdg84wCcMGxTw1k2Z1WpPdZMNqWJOcrohSE0oLJtNPLfqgi92bZGyVeNXqZWuspWQvA7
cJZiEC5ChTIpjGeivvH8ZtNOihQIcaQkb3vK14RnK60Tb6HHK3YnL57dWhacsv20c4nna4v01Zqu
CW19FSVAmjFjCz6c4ira6kYgT7fohqM+CYetG8gwLhsPGZEZhnjJKUrcCJrTjmfiL/3E/JEEuTrr
/ciGd/sCKn0AG28ZmnqTzGM3IdcMrykM/QxUE2xjJIJLJaPFlRTmPwC9pogKdXgPXehGS2X2tWcK
QXUYzbL+WWwiBnQLlO1yal4bIB+YTgomm0z6cvhCV2tLgr1mifUu/GgUKbgDVlhxSJrTnZxVqxKr
gCp2tbccVCYUDYZG6Z7WM2bMwRuvmQqi4FatsX8iZB503KOwE8WDH0ldUsW/cV4g/KpDVQlEGuUm
x+fHaDt5cRf1lOxp04ySP1WCGKqwdf1Mu2XjT0Dk/xBpKSjxADxdnfH8dQIjTuoNRX3qtVzfKwNq
Wwm5X4TGuNXgVEXJZ9rHlcYvJT/sF8QRd+1n9LukaRXec3khYbK9hz2+4v/n40RqlWJXfUUHz1wS
Q0FoNFy2C397GcElZ8TRYR0pI4dDMwv3Kv76Mo3e+oWHb8dL5/MuEN6aJMIbMx5/6qa7soDl1UBE
Z8lW/Ind/izdT9A38dnlWMo69w3GWK4LQClAvx9W+EMlOOdhJmZaQDp/WXKOUSJ/K49cXOoM1rFr
FeHwnixdclR8eyy4rNyrG8eOf0RybGqjuS11Lg6O0N2Q8uV1WGC9EM7nzdFTyt1XA9LrjT+UJH2Z
M0zT7ZbBwvVgNyTks6OqNu6nMx5xas+BFk4ggNA2GV/D57NO+bLc0bwszqzCFFX1vKEnux7+jGdG
GJxBrFD6HlFlx7q6Z6ztEF9C31ImkG6p8LrjHALp3oXr16WsIIbAtyF6/q31NnzPumam7utrogJ/
aRlRpWPsKQRja8fuvUZG0fc14e9JXS+SUj2p7jFVMa5plJlOQYuf6HuJDKtAjbQSS4cjoku/DU4R
XbxiikqRr9X5T1zytol7ScKedeEApwMfF3jL+ilg8pA5YYu+2tX5lZZgbF2liO3BAVovOfQj5uj8
V1exCatIEceTsppuNrI50Yt/a2whr1k0I7POrrfuR8Ac3n0vKVahmGmB+n2URy/EiDbqxg1hWl/9
DqtK3cstDxv1tw+TV1+wGXcJq+lss/eUFtW1bt0SWHZSOxFogFo7jKYFSnbcmAysO+HWiL9NwE0Y
NdNB4qF5TXz7oryvRpe84BocFvtaSnoKpe/MgExWW4powMm2AJt/UNgc9ngjjMBs/Ch31H21ZX68
n4jr2D0Ydi2Dggt9+Xd6NirybyHezIza53sL/AKJNx2PK+Nxjr1FmKEC5YSk6KJR6QYGE3xKvcIg
WBapK+A39TJXV+EuzJuRzCkjoszH2SNj8E+eVyDAMXe2BJ/nIjEAGRISPxSGsM8a3jvmrSKuEvct
KWF1dfGxrEu/2KrBTBD4SLjx6jKpPZUTGuT1XNa/qSM0Qm0U8SF+17u7NvIROKMKHDO2tBWxHQrQ
RQveOHVLAMf1aqLKTRtclamriNnwpXDR6myJgeIjVSpJP3zuVrIxeaMSXk/kLWgYmFyJ42At+uK3
CoK/RBNBDAsweGRyCbRjoBjd+q5dBK0WUADq228AW9+lzK7at6EKT/a6++N4Hz/9NfZj3XNUsSPR
yTUIZJu/2rk10b+he18EMZzICeK5Djph4mwN/L7z0HIr8idAJrGoEdTtGr4H3MnfyRfJnASrT17f
fqGjcYdrtMYRP+OfY0q9ZMsvqrY/y3GAFwKWt61RDgUfuBR84WF3ysnp4IB1OB0FAcJxs0Nb8nG7
rlRYcXmz9+laTqiBnaSBvHd13P+auWuClMmmKvACBf5GCUQfaRbO0COhUlNkM+cZ7NoyoIVhMIQ5
FWGzCScLHt80ns9ftxTeNP0dkCyjtkP0HABN/vRrPhUkzFTv18BmMrJKCtPsgZ2wrKk44R2QozUx
0hRmiz4qHfkMVzG5SxmlEatv5Zx1d4rpr01mcEJs7SKYu6Yc75SSTR48DuSCvk7iuzSVlXArWzNs
VxdbM9koltdEASbTqRFiir/AOMPE3q0NgfUzayP8BwLi8vdA+q4zqpI/9Rcaorjhrxnf8NMScEFV
otZx+1wJhFJu6cNGlPD9M8YV2vJWTbzonOBdGiZy8DEMd5dRrkt72XieG3/T0j0fk6siSq1dhzPO
hNwkeluPvTcZ/b4ZPH2ZgQyN02bRFRtaNYb/e6zklpmiLm0G7QXvQrImXIvf0ziJeykdpz/273m/
PW1/72MeuN0uGi6ksCa5lc+waPg0Ab8dNPLzUjIHcduBrpg6ogMlxJFABOCy0O5upDnJs7MDnMwN
adnI/UKqXVp0V4XH5fOX5fgVRp/26YXnLh9artcKVXaef83TtzKODr5NpVpZR1Gnr1Gx8MXjbGUQ
SmOJlKg8wMB1ixAsjefj3vLNwFG+ZnGfXxRjws4LgUiHWDwr17GnYByD0xqjaxtj6TqxttdvwX6Z
No5zOSRRpS9FJh1gxcP2YVyeTPXmJM5O70wxWg4qgSohdtiSNeHPtHxLiLa0GNP7JQFExSE/xtLV
7UgALblqz8lwOSiwy1k51fGXuYFtoESpawRxKGJ/D+bFzWyzedoiuXTn8BK2gRYUXzOGd4PQ2B8C
wlGEB/ABVJskYwjYn1EmkzHZIMUysYAg8TOkcUC7BQgrJRWP9Xm1xpVbctQIR7VU/7WQ4ZD10Apx
w+LVhNPjLcwWMopx3COri5aN7pKcWqHCKZnodqMwaVvETHoNX32VaPn5s1RU0ey4FJOxM6doa9jE
pB4haRmvcH2k9jRfg+ZmxHAmPx6C6qqyHhPRKe1hvvfFKoHvsvsQyRDlzBencJZ98RyY0c2kCVLI
qB9Dfpq7CunulFZzFw+6MvTBrTxKng5/mWKVDIa9Hh/0fe+4z1AIu/K3IobqXWnZdQphzdyNSWyf
I6yD5bMElYmUflQ2GGIZMG+On1AUY/3F4pZb2hJ7ALUCyPrFap+aR+xCUpkb96svmZGAlg/HakPe
qTc8uvREb3GyDQz4pUIdwDWwLoEuqVviUfqrFJoC9CmTWRtRosJopKSuzZgW3+IA3VLLJVpnIdj3
9DDtZDZuaytZ2EACoJuXFTBUBzeZVfa0m7963g95ZGkZwn1kUCNE1LwxJHNiJMQUyTovXpO1rvA8
UvC5YT2WY6Wzp6f46Tw1qJM4ivmUHnRyMGjszwrYyKQSX08GBdcvUyXCJ0R/5lH1+6kwg3XC0tjw
Wu9gMjzHUGA1JUsOGR2u5+XbqioSNXCJoY8JvIP285dtkn9YSPn5kO1BbKqVc4oh/0gjneqoORUf
vw3wtwajOHkQaHHtovcNRkC+p234M3e4ndAiDhckGV8stNkYuMdAeh24B8CHuy1djdJXPi6eDU9T
Qp42Jb2o6uY/sgHaByq6D2xB6OZDmcFWppmi4KOonLZ8+kkFDzZnsnAB0H4z4z635LSpFwHjUqnD
EerDyVcpBwiwy2611dPjGE5Bdjo8EthquEU1cVlpgsp4vf/6pbMu5n3gHRUQP4YF0JRWbDJ0l6M6
kIwBuH4WAwkLLIDSUl3Op7/Gv7zJ4uA/BejQZEqcPvTPiVCq/cCYyguFmeoGBGjokT0QcXlOC4Rl
KJhRH506QOtaaM6rT/NmiQ3zFHJMJnjJzzGZkCh1OF6NJyEeUSNS8vPUdbYWZBcfPbHqLtJFxWWO
SrG0/UOC9vKydV6aurSkCrJmQLaEaxZvDD00k4c6tloB1hTOgIzkWpPrTVWYSTaxdS/Ztn4CtaCs
zlRss2Cj5gnJU48pE2ouQYp8vQZwbDgp77WcMPksqHSM+FB7qgivLju6vuONUP7EBFGsV5nmEDXt
8ql8uMlqzbqKVxM19C5lirsmym1qyoYKy7dvw+PJUWiilQYyR2cSTUY3u4qOTQIW2BztpKgZWZww
U0duDjl+78XaXG1ccLVB04CBldNsthjqdxOEf67Z0WNud/u0+aSaLEHDb35N3AbJVPTNjJlWoWo4
Pty9Xo6B0Sfta6WI54FgvnPHQ0D8ehC0Yzr0msImL4j06T7uAv+7t0xhilRpVo3OhNbWthte9G/J
8B8VWH2Yp9D5hlnAm6oZ6sZ1qegoDnB8uy7+5miokyejFe35CXocf9mhjJxc5deyoWj4yn/ESD4Q
O0t9tz5yYVCZ45xaXY+CDCpmQyA1fGHeH3lmeyx85h/VDCFKySEhuCP7qRb35+Z5IjsT4vgyWGL0
9MS5vOy7k08Ywi0F+tPpkWcHngWCrhzFWAJ4XzVsUCESd+X47TBwuqdz3/a9huPkxoTDKmr8mJ3D
kETX3lb1dlXCL5v+0mAmqLskjk1Ob90RgoAxPPFVgCdB7Wiv+o98R6uS6lVpiGViWbCQIpanxNct
laJWaaLvEFKtv1ExFuvdA2tJURQ/x+GOiw2kfw/cYPQnMdJqlGBzBpaz8TgmEfkKo0m2XQBH974g
q23S2oy4ZCC+rqQHatkSLL7RakCFLeLMrAewkJqKLeV8g31dJKPboEc3//aBUfwgEYsGTmnLfsVt
EWiRWT6D9ZLGtc7owYvAUIto7+YxD0mCg9pFu+vaG5UIu3tpnWixwMuispq0TKFXVCrMLVF1wkMK
xxoy3B9B/2gu6CrgegN91YClqf3buwuxKyV3iormxtp6uwyDNMPdPHS1Bg/1TE8bJ3rMDU8zWpeD
0Aq8BpYpPSlP2+1+PWpfKyhnW7Gm1ARjULygbTRZkKLI47OV7QdBVajvkgAnu3OmauWgSL/ZyXB4
fb6BsFzrZTS3hIo/ocCan40oUngu15fSIZ9nW/IgBnKObDhXpVKeZGbyhhsjdCO+Iy6j8QW43um7
24dVQyu9oC77gAVj03iBIKyNZR6qSPoFB6Cp9jkNJv1Qi/BSk5cYz3FCgYISnMRFjBS02WrbxSnq
tAxpMDRAFSKccG5Fzknti8D0L/dnQYQ/skzZz4roHGJ31yC9cGjQgPCu8T1lqLXywm7aI1PLOaON
NTGcLcXW5/zBV71Eu++CDukwsl2cHIxgU/5/ycGIP9UxwtoGF+8VHtZ/U6KWbFCI0ONwmH4d2Kt+
KuWgc+FL4X5qH0+052TpaJP5GAQOkupkYnF79qySGYdjixhJ5X8ekcb9h0Z9xZQg5S7YeJ41t0wb
+nmMAZ5MFLJyXPNFeqqMsWsvrtQVXmnFmI76mr3Zsav3ryEweGBTYBHR+6++6w6I7ohQKe4xjMKx
ReFmO9sK0oGKSYvCkyRnlF93WqjjJXye8qyFKXibWybHjEh9YILwPfyLylv2B3mRGUrXVoI4UrU/
qaR8UsFSsEHMVAe1W4u4TclEqbtxPOWrGXThE7r+aVMt/lHKTZXZ/kI6jI01oqboCxzYxuJdOgac
521rmDe2xTG2+6+ad1py0WG0eDxRLGNKmgxww1kmKLjO0v0gPyWOvQSxNtDBJZD19FLcDuqJGzDk
6DGpv3ax6pM7EE1p43Fs/8clS6M1lum5eTB2Yx5AXLlQ448kjMtVb20aze0Y07hBmciwR8SyjleU
uxSRH18mIag63872wh0+qowpRyy5zjiATBJumjWXlh5ln0Dv7ZRWTiWppyq27MS7lBznSdskta+r
QyHnl7N8PuNAMAj7S1x5Fy6sLieA0MJI8e3O4b57HUPir3i22tt+VuwdFjkN8DTSkAb+gjJFJrvB
LtTvKACqkhu4Im/rwBGrm9MAa8+GoyOSH1RS0mKC9oZkYtb4kZWugAUEMjCRGFh+mDXjyQbLVu6t
wjWiB5yLeYLtwjS3dE2h04wUaUdGamS38cgv4F6KdOhTtEiUYcyf+mHGSxHiYiSVJLSS0t+VLL2S
p8nEtL6Mdx4EurgcZecKRBDNjZqyDzlDAOUG/sEC6u8tbZXZ3fvG2PmXbF9uF51GB+omW1IO15df
1Pq9rSOPAAwwfaEd/2lto9es304k90vtQzYmMR7ay9hzjHzqyeuHcdLvSNp3GgcvurW+fvDOB/ga
JjY7WFqc43Fo3OFNrvY+Tcn9AuwVZOUA4e7rQn2cRCZtg73jzVG4JbeBiXI5NORASKCdPcgQSrLs
RGdj+kNBcfVwTz60XuVe59SorlDxupHvA79IXawheQdcI08X3ErGz1gIuJI2HF3Wc5CnNaI6m2vY
Lhv04vAK7XNIWQMtq2kMwhotaJ73EioAyvCt09y/CBJ85w+H0DUodcy3XvnjeG5tTWbQs6hBuMp+
mnOJuRn06R1+dhWjK1a+u0VuBkBQwPkYHkk3gl6lCqynGYm1EIgCc8ufzDeetw3mAhnRhXQeW0rl
zbOnfFyWJj+d8/uGgeziiJ8wzON/GCQwNse8OCXhhMUmlxeOsKKTYLkkvsOxBKHGnN/ZVNyAt9Sb
aqCf+J5qT70lImvSFmsLnsEBK/mY7u6LDfXc6phH2yG0n3n8C0tFMAP0sLBuAmFqFUiqsBqKcHu6
rJzfJrw6tbofgk7H3pt2HaoYMoYmVVYvmS6jVHDFuDahyT4sKt1iIqrI1uyU+ucYykP9ilAU3Nxf
HbW7DOpCql51hM0XUQgRdQLKqK3vhiT5fUuYIANXDzP/jbnvbdgCwfwdwx5+EahSVxuI2rZzIX4s
abSw3cq4cqUcGViEpTzsFxoDIHb9UyFN5UA48uenFAhA1rQ0PSeeRxIBGvvf5I3t/rjboTNBeU5L
s62ZeJVm65d9g79y9Jiw13278+nZiTy5pTeaIIdP0BKWp8FqK871JsyjzP0yExL2VuhEO49sLQTx
q1NzKOpkyvfp9WdNeGY+AufxToNlJDDfq7bMa8SkSb79qkNMje9RlZfQ4a1Gs6s9cNqRJVm83YaC
d8d93YNMcmKM5VzGJ7GncDsjOuO5QIAMKRWn47XAaffQ6wHl3mblW7psT6Pb7SSm83s1gIsaVTKw
ra7Gh54oA6E4brMisj+eYnnat0ama3eAYgPvKwc84HvvTmWue3aOs+dgw0CxbSw5bLkETsuM0nZs
A7rJhKN/IT35O2J9M4Q2P7Od+Tl4d/UvNpneYhcm+dVIeMBMCGTb4zgwTf+e1tRd5Ei9OTX09P8m
BICcrJUehJUphXy0D7e9mB5knobrGebz0pqTAe5NWXc+7kHRjxr85JP+Nlx5o0GamyFVuO974+oY
kF+t4v26TUfeF1bIZR0WKjoQIgesR+w2cuL0+Cc7aZQFdTfcVGJm2wItSsrZvNFktQF6nzMBbvdu
hxsPFZFBKNytbGd+hG1smixg7to65gYqcx671omIbVEUGeR/FTzJ0lzH71sYK97PnT6eUaqyY6Vk
ORMKLWLeYTH49J2v1bF8QlXS/pQyDvbIznsjto6dtrR8mMUttwHaR/fqgIjPrBFQwMgFMdcsbtcG
xShsDAF3ZOeVTsrgi6BrmBC/VkiGto2BegiGCPlxjxBeZEtn4975Y4s7be83UcgByHKjItLDXzHN
HlsPSCMOa5UFOeaHNQV2fXbUWtZdi5oXheck7wP77pif21giRX2+AIj3xUhwzThbD04F0NX5hEIK
BNy0tJBAtNdigFC2/i5NJQBG0v+Qi3vgydHcWr1oj11V6+T0YLsGu7pQ6fFzHZuI2JpGUjNZoGYD
QqMg3YlcsFtU4cZS5pOFfock4FzbrhOeI0+yhQLdQIZNRs8ML/LS7749ipFhRP2NXBOeKBdwsXla
ALxHzPCvbZoARJGpZidbIUgt4TMgN7F96mn9Uo8EaEH0PXC5880x3liXPwaZ22NFdWMZq1e2giBg
3T941uknL6NbD3AMkLov0hiJ7e3O7edbXVBI4siMJw56i83FC0Y4VoW/VpC0BdW+d5GhPPIpHTbl
zlsaT9UkdZyQzEGKsdSBqKuqQFyxMfWTK3z46+fK7b9ZZW5G1GJtLpFjP9LPsqdP1GHFmXOVZsVk
smhLf0T2pDYvq+0f3Pfa6aTGJ6pq+HBnZiKbO3LJKT69riK0Ul+miKY8KtI6kpTCZ5oJpBrzP9HV
fI+l/Zw+TmJaVElqGkZT7ghcNVPsYIo36BXNEcKXYPnhpXUuH7+WD2PYYtuJd1rhXyFXTkpF/qNW
GgZi2fMEpqWCrZiVoqXfenW04CxHfzsYjJy5GfW6XY9Z1Yyshjf2wWs3XeAOvkTxVAl9cB0nsFU2
2JMWDqivqpcBjz3vksSIZH2kQ5Xd1tVjKKB6IYyfOhHZTvOHKXU6s/ij0qRlMqmtNCL2L7MPvYTH
XrZgWSdNCDjQVnCbaK9OLW3/GfRX9XIMjeGdgxVqbw5itORM7CgX66SUcKvlEK4Kdz84+el34ZD8
eCLGL6d4KDNz9TLFyGzEakbi+oO/mIqpmnKJGaFNCT/bBnYnFkYV2/Xv618JgTh7ff58xeZD+x+v
CjMhdd8SGMkF29ODqIu0r6OfgKx8jKQzaDHRrE6qGVcT0knAfcUZHOOadolg6zA4kf0OO/umpYCH
BO4XP5Zo60d/fFm7vt0JDoG5NMzuriuk9NIBbtG4ziKny7j1IhtcJlqYlmHo0iDpWKTvatvFo0dF
FZJpRudOYihlIvn/TDkqQMojDGwuIUmHRc1BJdgDqij69p2namw5irhff1vuUXYlnja1AKU+D+rQ
hfTpHsv/n63XFwvmj6wH8iR9DcSR/ekzbrKLNI9F6yxOuWHdQbYwZC6qpAf/UWqvMRm/VAborXcE
ERXRzF7GzvU3Dt/wplphXOozj36ED/UYvKqPZ4t9yfx5waHK7Payu8a6U27tjxblYYqjdFinV0LE
Q9fham3npFtdDqqN5xRrtDSSXMxGWBJXawdCH6iz0N/JLoKyJpw892kxPI6GUsNc/yAIG1hNeFtW
4J9S9hlwp+4Dm6S6+3gJACQ8eCbDI4TopXDrkGEldqXew0sCnSa45k1GJQOkT//LI4Np52dZ1qc2
LKs3tqfK74QMM6rmzjdkKV5WrPOnpycMnMQqDtEHKsHOrqO8j2Z+cxhq84/lgEoa1M5/HIpHDsg2
9Hei1fIp+PQgmKBnoPJZqau16mzitjMfILRtbw9xx+boqDybe0TMRnYE6npgSt/vOOhskMymwQ7q
UUSJ94IGTO7/We8LZJklRtXk6/fsi+kNIPS0STw52f0r/la+7FBfIBwNsDm+/a9CvmaINnkR1u+A
cDpXMfuiAW8YP7NVinNOiFoiCqOiB1C3YXQQoht2CzKGqgzJT144iUyJYS/IZbUqNGs/LBh3cotr
qNRPWZK8mwltG1XtfQitykEwMb97tHS69gerbu7t/5wkGjY8IPnum41cBDd6I1+Z8OD2tQlitjDP
tao0Yeph7IcA5LWtaIt3oIe5raHwBXRk8Br/cs5UT4KyxINLNIG4aeZ3Dv5uW+1OaKgVtpe6A1xH
ZHcrxbYue8G36SyJfs5wHqd1cngEECJ5pSiGdo0z77B8OBZfUpKhccVJlnipIFYYVoUhyFib9wVQ
kOd8vhJrvsm+6HJbDJ10g4RiGCDcTAGpFejRccO1wsN80gicApGVdfFKkjCAxYOY1GhB0YNwJePO
QTA75CiO346rObjdRCwO/LE2IvI6CMIJF9SDfLkDJR+U+P48dERmSqe69Mq9JvNpyAQpzlZKEFoM
eiFjog9cL5vd75G2fvCIqwDH2gJyxab07nxLiBzoKHCBQmq/yoE/vVlS8VqYgRB53TGBKuhmNv9O
gz/MW2GZm1PzEimWfqGbfTc72hWUCy278IyDQMOSPCNnhOyPcqdYL/FNyRP4kRZVvuFy3SG1eK4w
103NTK6A4iglqhtyBvUGq1V/uiDBLveVrz/7qCxrwAEggFHtzoaP+vYJPenBACfmadOoCmy71qrb
B665e7nlySxSGBW4bRaNFu1rxaWgOXItmDTkQzyt3ajNIfmMer9pWxiaz3ZLJOZ5V0HfBtiny3EO
eOsB0GL5qR4cYCDT2HzHMiI2IMM0i3YOUeqQuooy4l0YUVhKSloDksA5q2TwPW1SDR8ehudhNMmI
sefuEl96E1wTU5XTn00N4iYcREBAeHs466KLZhIsUXU21PebSN5k2JcfB0/2R2VQR410fes1GQa8
fhbJjrHk8jRxh3jeQ5Ks7LJHhGjNgOjBL9rNTLCSb9hquli/h/aSJLAW7SVCzNAa+k2L8rdx20dC
PfbvzmP9/rh4KakOaxv3WSCERbRmVfp2ynnFwBT9jpbgr59oPgcKE8M5FUZuRA0aPBy3L9FB57yw
BnVPXji/9TM7GzCCL/fC4LciPEKrVXzqWQC3oy7U9Nl/gFhdzcC/8Kq/i/8RdGdBbBgbGGOT9sPB
lIO7AY1MEOSzD//1CCMWbxFqvdOux6ccR99fFlgnHL2qKbp18BVq4gBpN78LdRaJe6vXHpGLsoIG
lqYcXfXdLtAUtuTTqLYdJ/DU3D8uw/3LIj2yJ1wDfDioVjDuWk0/bnHQ3TLl++4tnfPOViehExuD
70mxbY3kHo1EEat1X18pEnv7cPrWxQMtXRuMQn5O/mt/rrMPd3s1Z6Q/E88KwQ9/eldWaxV6x9xp
OG3M/ZlOc2uVsxVV8hIVu9aGjgWR/rYyzoC8/ht5w7ZTsSL8GTo3CcRZ6Mwe515ZVlPRIF0hUqkE
Tbn2DoWDq7qOiiKQy+rKaueiZCuznbJdjgsCgesN12WDnux2D/aei6YxtUoABCo8fzQW9Dlo5fI8
gKq6DHFNJs1RR9BrjCR81R+ezjyhhBiHN/ZGYUkCxM+ktvaen/9pW7RihPeAy7vmAs4jpNvDZXqj
kVcGKurIEduEBrhPJiM1sKMH4Qn6oQfMmzoqDTUDvtWNRSw3632m+CktUVCC0mG26G1hfUA77vs0
9eUy02kS1K6gUZnTGwNdAnhLgqN7WPHyIPBMob07JQCT+NeXyBheKI/rg5IyMZN0+WekCEmXIykp
2guj1do14iKsVHeNlr4E7jRFe/2GU9VccDlty6KjRuKzAzSlNmE3R+SN+v50qcxzQn0nfatMuspg
/e0Cu1NNge8hgZpRj+nJmanmX8sfmiDdEmzpE3yAT8k7/GRVlR8XzOS/+NPdm0xVG7X81+b3VfDk
aAUs6SjMI9PQUEL8YRCt8AW2oV9MLlvy0UFWCTy3SRvaxwJlU60Ms/kBr2xsIm78aT82FzMTLPUM
TudGM3A3uRxHZgF4vjdPPKMAlcr6CHcBTQgn7VI4P6dYCQsm1vl5MC0zHruMTBlf0ypURZa0eeuV
RU0SfnMXZfGG1OSaqjXU6tjJ+Boo2ETBDyF43O6VXZ0/oP4WLOdzTK24EG9vbmb3DIuwZuDeGiM6
ZY/Iy2bTjM/r0EIs9zTevqAgJixfTLHThFGV8EyjKZ7ah1VFY1dTsQf8yT+QjYmGXuTFV/qEUGeS
yBa6RT3WlF41cCLAfai5Pm3ZgWWX6fRP9NBCKWrkzsorX7tCCbqCUwWCSnJtVnJqxdu/znGwVDN9
i524PRyZGELg277mtaZR8CMQLdi0qA8Fl+wUCTjoiS1r9Qpz2QD/eUG0GJvQ5nPzB/tyBLiJPKhQ
UUALJBPmlfolkzFds1Qdo0if3r37gFG+xGZlg+ICwmkEnIBXAU4Ehods5yyrJsPZ9Jf1sKZY8Cza
XH/nf9kqp4Fk48ROmQWkYdwWJSzWJBxxigzyeAK0/heOSprgrmX+RAdEyttOUWbWPRgpwV00UDOK
7iAg8UZ618jG83QoWvq6xXheUT3qzn2Q5gZmHUyOItJHf5XJKuuedRMAaiXWZ76FgHiTKnEwu6ko
wFbABq4AS1U2I72dO21TSTiE8u7a8MGJak5RxTXf1oHxuF3mxctTi8/E2Sh41Mbe6X6IIPiKh6K1
dD2hhZBpFd2O6JMs8nJzWRoLqYFqNKBM4YIr0Uo6JrkMl3jbA4GbMWgCIi65U7mqzV7iu5ULJbdx
ruFkqFPQC7d8qIkSzE6QJGZ2XyJ0IhUvStBqvfT1nKNrCjpVUr3VwBpJhPus0WtA+VmPgvpGpf2s
4WdVEu0ocnQGhehqarvM1a0rX14h2cGOeWf1uyv6BkfF4KL/BOr9quurnxvyOzUGQ4sGafguZRJM
0SwLzdhTd3W4u3EML1XqJHmwqtWWUa7S60jOzONLVxO0E/rBiekIj6jCzhnM6WWd6+yYY8Ni7v4L
GQJruO1tmaa4l1Z6WXhlHyL30m91P+Kn7UyCbImAg+tboTD4I4h2agY13MxfR6oHVuKJ/TalYa8a
o7cq8Spthgxfe8yBn/JXGp/XumjOG7UYx+jj1lAMzhdoVZEoEDCByqB92JpAhGVB7492XgpIM98A
NwIqOHp84MM5pN78k3hJG8XySRC0kbE8pB89nsamQmcFJdwsSmInMJPFcDtmrNy+HCN9MNSrGgml
Hn/NYFiQY3Ei1ms8m3vBtW20Lenozco/J1eeLdt/R2CHWiI649ZFQhUzc/veCEhZ+NqKAfkTsGBL
k8u1uvdgjqAv7rOy6nx78ylcdvmwTYIJWqen6W9vnA63AmBLkfMEY3KbHntZ07Qa+D6wLHDLe4eO
/QYFtvIzNaTFUgfmJunlAOVFye+kYlMLzcY+CNWN0dO4E+/URQ5UC2x6d59ICf7A1yhK885yzxe3
4PU2QpFzMEW1OQwCFR4oTack3ZwLd+3oPATOO/bulh3CGw3MALWZS5cVFiIqP/cRywaq/UJANDzN
oXuhb+wjSKtWofHwQYPZOWj/nXdw9olBKSXsjGZpRoG/bRnO4radLjpbEVezoUDjPzdLTK/KZRft
Qji8RVx2vv4AjFaxq+PPbHi+PCSPEchHf35tQa90WRRs+cRAr870a5B+C38AUyeMUY5s8unxmVcj
ZY5YhoEygAzdoiv7Hgv1N19fIiB9xwPNXFlU7i7l4ystZf+PVgmI0G3pzjGTdk5/w+2QPnTFQsns
uhvX/ljvxOsJEw+9EzjLo+Q9czfVC5hHY86bLYSIY+/4X/bHcHrHiYzobWhP5gH5TS1r0Yzd/i1c
JFdtbR99q2gPJvLznZo9HqHMTHoZ9mk9LfS6K4ShAutfCmilcAzRH4He3lVDNTbf3hJBxE4iImXE
drqeibmmfRqOod8C92qA4VcjJhhGYXGJuJe1+4nABQKy3s9wCkG72KOkTz8HiwzBEN6aho8188Yr
/+vAUCTACJSlf5NSb1YX0uRnImg1Q6BilbCWuSwMIOZTYWZ/2iexyRRBpF4uiRprME82iuzSTN1U
enF0aOiaeEU8UGR6+rqHBr3GL4oKYuRUfBBoOaPfJlMz+2sxaxAylOfpLjLplxvunoOp9iB51yB3
EgUUAmjziiiKbDgi+Vl8/7WeZsTPLVI0ejrj2B0tuuANG8wv9elYr9K8ZXe8HvtJ3zdJYig6XVGS
dYwzYsGD8AyxzRzR83UF8aq+plRmwEIZcnrc0FsRwbF65qTO9ypY0r7qTTofVwqsMP3O1SyPvNu3
ymWHBykdDYuU/RL8bnyFmmmMeYCMvr96rZ2VHcQf+Gneg+61LQOJae/k3DuOvRZG0P3gfbu6+5b2
CzUERUfXu8oM9wT+BHHkCGkKFDqrgrA/KG97thq4wIk5ibDiebhaD/t2uc7s86VsznnQQouL6HhM
pZPKdq4/JoKZXkjO1Ay3PbwBReqd151znVvAjAOePiRJnJF01Tk+Vf5wOf5VNUo/LqPml8PlO/PS
mgmLq8m+NUkNunqijRvYGN0pzPdyRTjzIyEusj2vChZBwn+9zR3dtMJ2L/SKQaJ4OBhe5Tgrp1b0
05gmjIXzmmQsP2KAxXICR448eNY+xtK6oxSjHOvFq6EGw/R6WiXjWF0Y/aTo/WFCZCkJMMirY8eh
wyHTZrqTRW9J1MW7nkXFeccEwBhQleA6bHeYeClieWCn33XUa+Heq082XuAo9xWJG4fkQFnaIMuY
rSsKl6yWt0JiwgiBUSfD9EXvfuGyd2c3jGGPRb+/HCSmzPHU6GvgWS+xK9Ajo+/OW+r9ebRTwiVu
fw/PaD6jPwQD4E52kykcrgU6xl2ENwzxWoi2ga5Q8939nbxvcB2WAs/BbHP56gDotPPPPs4Yzm2i
gyQ3OkLxX5SPalEG8OqjjrGKp3kuN6DfHUFd1neDkUUZ+Ql77VTzlUxcBQESRRVlmJ3sWtUOOlEE
MoW+kexjL11cw2k0QW3ycv1U7357RmWBvzyZXhfu0wMtJR+SFHX6pL2KU28cnAC2YS6urLFg+/l2
83eqaCf69t5FWatx5ut0EFBXS2PEKQ6zSO/Lv+vbCAFsYJ0Mz0YNR1IMHEZNlD3v70h4ar3M+XfF
3IByFgpfLcTfdL8yvQ3Wq1ChdNy+mase6wpS/dWz7c20Hc5iSDePebCubtN7ugAcCSXQgHvsv3J+
Mk+3zlXmeCSJp1tEbHEsxp129yH+h5++ro7pmG1ZpuDQlQ7RXIWsbWW7qTCXbGW+DaNA8EZ5Z6YR
GjUOg3w3CfllRTX3Klr3dVebz7VKty3aVj6fE+QbX9yhQkoYff7hzAol0N9kZTQF0+iDuPUgtJvQ
qJPK7ezl/U+vRJwHZ+/T9u4tTZItt5oSbFNGB/a9dkLEWCtH6FQKTpk+ZbzBFw0yn04wJP5UNPos
4YKK6zCWY3l0IK3RO+NrMZ0h7deF1M968B7oX/C2UM+uL+JZp0y8uy7J1X8zIjNd44DrB/DaLEx1
qRMwY+gZ4wdo055DgdiJ7wBuTY2vA8S+3E1gn8LXxNzHRZTeTSWPfdpWHUZUtPHwjEGl0DqwU0Tl
OvdMvXB6dUJHhjT4O9zPhmZn8Hv4ME3ld7tK0kiEiFOSPiZsN7QFPx1NdHMw6aYpYW1G9vcRjbQs
CQ56kx5WkkqtKGOpJYOTW+fUkP6wwItam2gsnRtMLAQ1kC5nRgnIS45UHfGmrxNHi69dc9a71Dvi
6fNRjBDCSckIrLqSLgbiEneaMRPedVWZSxYBkSAQWx8R1Qb55VHwyFOxPUecq/yUF+Hlse1SxoYY
qT//xUwJ3KQr9LemOlGpbbJC6NI1PCqYXS8cFUCEXNynUP850+/iqYy2DRs/+rKuXelVp1jxpW11
8dK4N24EC19psCzjVeZdg9izUGF4y0jbDx27PjPPqzBluKsrDWtGpd3iYH4NAQ5g/D7xtNejCqWN
/LyC0WETkYsoqwPOjYmH+sEJftQBMofjccP3hVGNPuuyfa0yoot2+6c81SL2ue9XMUQgBMxPb+zH
nV78daNyAXxobnjp50HNSiQF8SC2gjG2jc2mOvZYcvMEbXnzvG4gNIYbEfj3I74BRV+tIfyOlCHx
o0PxvFDgsL9ScNYi4NVkpHhJPxUdq0WftmTMdtvTKZpbZTu9yJYBcz4b5cBCExUDeTHUh9ki8114
qmeLkmKYHgPxoI3E0YzA6XozAifOsTu1lOnicSNZEGcHwrBqIMFhN3ikjmHDMKqhI4XC0ljnaEDl
+OhO4K122rXYgrPOPsxOT3eDc80jP+G11aLme6k785CGgtV8nR3Xur0//Rwclarw/g9Vz8gAT0dI
ZhOEmnvRdgYZax7yYhoguhh3zaSO1NTHFyIz8s+IcDUap/JxSaqVHELBhagcv7m7R8+vbgNbV7ni
GSBDrCI331MkgL6ZEwdKI2QaeI6XUmDeVl7MkYS8XxXcUFOUqIq4WFQbGMBjhqo0m2CG3a2iOoRS
GAV9E8aZC779ZPtKiCRwk4ps0EVFCJjkHioqSnC1BIFC6QE0LDDjsRTM+dtGfWIyf2LuQn+KKFmO
IZPd0nty8Txd79kXqnryWrES9V+ZPXR9dpX7bHq6zm1OqavJGnRoojCmvq7bhvHlrbuhnewzoccf
tQuzV4OSUBznnvnHqSbkdNKoNhAl4K5+9ti4OnYioywQ0XLvRXFlzoWrbTdiPln7h2h1inb6OKBg
VWNoV500+5Y1jX25otjzfMcn6deEYGlnMThblSKisyuRhHnkAXyU7myS7MlZbt/7CkllXAKUzAq+
JfXHXszvUTBFKpWyTIAF403vekzlQ0XifNFbc48hhOfPZY+NM6KkgWfdv3RneN/8ypDehQUgKIMy
yeeVqtwkqb0QtZ6zG7Zx6j0gisR+bRD7EalRrqo8Ho3VkFLMnb/jkQdPQLzueCRRRXc7A8m6CxFy
h77jeCPo8t23Dg/dglLbEC8Nzbsoc7MZAAAwk86+eZC/J0NVOtsH7qDxvzwloIa447/IJmqM/D/U
K/SMCf/x10zzZepErc4ES1scTW7MIDqpi/LK8zcI1XoPTsQqwD/Vpdva9RDNQ3rbiiLwn83gg8fu
AM1jZJWFMhaq74EFCFDTHhCZZK/CgNNUuT2/TmbAy+nWIgVm0JMVtM+aOswia9+0ZKpun/F0eABC
Zq+58Q495Pv0ulW9eBvwcZmLBJ3c3J8+EWiJ5chvnoyCw3pgbPCCZ4Ek9fDLfiCFfd/n+WVFcJRS
iKj7Hoxv+n5TiQAi7v9/JPfdIbmoGebYWDaggf/0KtBGWju7I5bUWQ8MTsLrcwO9gPRCSrCz4U+u
fW4qNFGuSrBZmNJMjOzskn03YprsmN+ahw4e3OKOuAyXrbqg4cI4XlQaEoVfC8DzfMOM+WeTinew
hA8i2UlvpkDv005chyLjDpU/Mq7g2Bz+0fFffdyx//hxS7ZLpvgt56XytIpaFaos5T8VccB9ccJF
SmWHgtJfppeAiYOh4o9VQ90Krl1t7+9EY6AuYbI6Q9D/7UWZOrZ/LMC0YBPBRtoRDcE1NtmB9U1M
uYYEnDpTD3oq8okuqL9Nn6TYUZgRM+Kx0LShSpN0n0rvHxuVL+2RdWvyJAWGeHDb10clNts7t/HL
yocGi6MToUb0EKNAIxHysnye7rns1szSrPETxaB4IjrTZh58Ept4E/DGWHAoz154GA7juIiKBXRB
q+JcJYvO3IKAwBtx2QLCC6BZ2BOtKBAOveM/dXhwCxYi+dzQaI2FZE8bqCnnZaz/gWBsUau0UPRH
ES7P2GQyofdmGVcbWUKhHv/7Vjr5jBLzb3O/MS7K0LacrhShOga/3Rdl3ZI6bZPYv8myq9HtVmAx
NVljQvR3o49Z2Qtbnwzke4QtpvXYEaCi1YGtgU78W07SVYnnDFI5y/NqEQqjX7Uin0Nl9mkwKuJG
uBT1B197iY3xDUgiEVs6WZLlgZjYVUdULLoFZPEF3vUnW36GaITgmoFPFZrXUY3rafG/QyTaacSE
9vr/bdhrFsd5n8b4NfuKsrqAghW6H24PRyEx7/3dFKQqX1pW6Oi6Cyd8RG47Y0CBDYislYGKbagR
KflH8KDTiwiEi7dkR17QNAK8BH2TfKw//mvULvJuFVvGVfEBkHX8f++HDjg7RUmZW41Ybst2643z
/esRltT90SxjM99PIyzvsRLCZ/BHGNTF4llbPoHpJBu1uMdMkLyxebM0+2jNrC36akSWjMzpFpD+
IWv3e7oKyeHOIXrjL4EL/L5AzupH9o62Pw1+KqpH1R0U1zhsDWrQUhYj8YCOq864EshzcZhT51E1
cWmAKpyj9KkPTYOXdP5xfsBPfcDRqNxL1VMYydo/KQSvLoaV/vRu4lq3PRNQgGakes3kpFUL8qOQ
0ydgcpMElJ8SBziLcz+iuj1iayZqZEeU3wJkEL/x6PiquLIJwZe5epE0QDkfaqKpekMUlGKzvyi2
lbASKTp6c3JXdF+YozbcSfdWb3pjmf43A9QtNriruQxcswcVPwNeZtX2joehSzjTDFd1XaQnKqsT
ArhwF60xybBkdXUaoqg3fr+Zs2n6d/Ylph1xiZUWrZP8lhqYtMuVcRHNv1gD7zl/IUO+rUKco+Jl
kTkVl2yedRAO8lr7ScmyeYY/ByGMk4z/xQUHbQvWwAtT+ne9smynda9M/Rp7xq7NBh2idaaYLoOo
gf0K3PSQILU7baJw9UUK6YTJR9qBJFGgiBYYNdzeGREqQAacI4UDGIy1lGtWl7LRjKdchUrp3Txa
Tf5ag9RB9hYhk4lzvaZU2dfljW1nvd8TWc6hPyIN6i2INR1hnrqrx5DxEEF+I4suKPT3QO11Fhnb
uxPEfqHL4boVFZDISM03DO+JXPRebpY0A844Wpmrr4fq5DqIg2ugHvWR7rH1tMqGDyHuP7ciRyjx
olgtAE8wycJQrtC7aQ4EvXAgOo5vLE6itHQErJTkQxkeeF51fY0tF9IS2W+voO2eFihc2J4p6qyq
4T2bwvBGURmGZ2rkCNT7Jzp/wJB6w6JqtBwVW54hhFYQJ7Ox7Xo9h86ki82HKvcPdym7hlixwwss
aQ3Y0XOUYs7MUU6ao/RsHyU6omS3fic6vrd3cAD3FCcMKIzkZhYdC9I90sg7KPMcK6hIQk7K6C0s
Zf3OFMZA8k7I4ch0IEggrRRuRJdKfxMqm+SpvVKFpsc35zOmyESqZsCmOisFoTirp/eZilddzrxB
3kXTFJcPBKHnQPMDaS4kyUtxlDncEcKUKv5A5S9Yvo10aZo7AyEbO9/RUllRgD1L0RQRIBykWYG3
JLYKgRtF/xx86wgCfuHH4dJFsQptM/YoovTD6Vr+2WAjcYCRau/kp40ldaouVhLxmunDKobA7I3g
+X4JQqJUo8z4PqsTd5mu6ZTzYBoBIAqI4k1hcOOQfbtnZT3FVryC65+3kOpGqSeXJBHvm/3rgfxy
Y0VE49S5YBuShN55knavVKSumWFfy1i+3NSImVSnTiyCDU8ArCL+DKoCesXOJsPetrGIHNggO4vy
zJtAMRCJLEakKosRuXny8jg5oyh2PXveqQniakCklvcJd8U5GlHIrqJctvKhwK8hGS8hvd3omkMc
yH0atsVewmjVAdpIchJeiL5YWwDhnpopqj/c+TDWaVPlHg38tQTWENf7ESC+ovA+3tzg3A2g0nYd
97EB1bcdg3i9SWND2ZI4Ji+NKo6zqAFRoPT9EVHVgVLOy/vPGGIrDjCzW9IuYM1nFH6FywKxZnAN
GMtx40dPLJBfcow4qslmNtz73sBiMXq+fQCBRo0VpX/C2DjajHTlmDdaAaVLDeGTT2QOqKd2zurA
Sc21sMw4F39gpR99NW22vdec4YodLoKlnUP6qfB/Iekb4u3UW8TgRc0Ksn3PjAU1dARCnTUc1X/C
HvTsC4UsdijQaFzhOh0en4s4okfh5TjXH+cpsINhTiXgiHRYf369lZJPFRNheiWdBJzeNXq2xQbE
2VbtOeSXy60Q5YEuOQpuBZ7aBv4CiIjR3GHY0ZlyOp3r10Q+Aiz2Up0fCmnQr/fs0NEu+1zuHvUi
GvNrvz4YUxZiB8WzMCHc2TlHppBujj/3BsKrhBKzGnr79zxmZbwg2IRbmSFGOANVcjnSb4C3Gvm6
Cd5yqZVyKJJE1u5EcuhzbEmcQziGm3013Ph6Erpx/4Y7v4KZ++f5xjHyS0uQQiYf6u0hKLFoLD08
CSPLkMToE1HCJ+idOWv5/rcWhHanE9B2jErqSBMACBnlGZR2bgXkRI/rv9C4p34iU/09MTHla4sB
sxoN3bTAHe2WvIqKnmzPQE7PSNkD94i8wQfBJ/POsq6GfZ3wNLxFdLcziDP8HRYvTbCcKdfnYNdC
tymW/FsIUFNQBWfe9f2nz5r4dImmpi6CNgn2KwuDLC4IrcPLM8cbZifJyi4MIZooXcjNcga3ETE4
PYJq85I8UHqP9YEaosyfJLOfH9APduPEDqME1eQehh+jclAJNY8/WMEXDq+Xar1F4+IgdsBHM+4G
zwac2rQe/LbczDgH8re+j9OBm2JatSqD0aXpSdIMXfu4jADhiItba/jIlCTreV1xB8NaxSbhjw3o
hrj8yer73iok+fRvB4WaurIFR2ZvOfC6H94qd7+uSrFYtM4/sowXiY1PRaD413998yjDNomP2OFP
2WvwdZvy4DOj+v+3SkDgn/hvrd10ggicu/uGU6iWRo+HWTEp7Ig77rFmkgHzi9ZCgvLRYoCOQEyD
R2+IXu644JhUw6N8cEHv/EPlfKJF7zqLLd2HRHHE/6lk/WmQy0guSLUFWC7fw/C9xXO5Zs7k29Ij
JVtpBoKbVLyZgng1yCWTfj6vTF10a0CpFG6atHSMc65PvQ4O2UMrUobo7rONtWYzrh+M/nFkSgOG
89SEyU7EPgNKwyGDzsl8Bba5k2jjyqXuKSmvs4S+C8RoN4j0iOuezvJJf2ZMqFv0QzgjIG23dCZC
nniTq+7APPpt+lTwDoxdBC5JI4CVfWogPSFDB465pXXAilBxAEPwke018TZa4c646zyJEffBLSx0
MSCN5EpIpgrU+2XPZxmB4Q8Pm5d9cb6nnvIFqQN7WPKEETG/tn25GnPTjtepHCUJtwip39lCOhP1
NdfDh2MA9kzWhrIezSbE933EnwSI30ubZxkLfifXDBgqFiDtIj6JCbt9rFfw2Q7I9N5NN/FoLk5u
ckJj7VVLFTodtHpoJAZtpDoLM8bC7ADRD8DrCElKgSFWAKC1ALfcu84PPnlOCMYB0LJt3cM8IBYA
UfAS95oWucoaURN9p14BYUgf1nszBjDOb2Md+CMQcNMm6IXcHy3pJVfc0PwpZAx/UHYxBUq+TGj3
hbozSNmihmzkEQxz7BuB0nv+7kUn/aBPKrcrhS8Nhcj8+fFPMuY+a2XmFvjFovtLp3Tcemtzvf0f
ayrvIrldszmwXCYhiJEVjo8d7PCefuOzuZ3ACY9v/7xJVGT0Mz2Zgskj1AEPsxjxJQYY4yRt7NHS
xyf8BNW/zXjueNytj+ICuodjfxRDlTjtWpjEbT5Km6KLxRTI/l56Uw1lWuFFnHP3CkEEFW+2u9HC
FwYQHushWfOZ4G+4MUQ6+qNv3YQj+XjIZYwkAM9V9MOIlUSQ0Sbewa24sPxklNNkH57/Tr+OH4D5
Uhx+Rnrh26Jmby74rRT/CivYDNypcHwshLW7lY1LR/eUyRASVIdeqERnMwJBpSWWRkSr47zgOH3E
uFHB9rEwUDCazf5WZDRlqjygUoH/BYDtd4mv1dTfUDjCDQDYq7jSuayecSgUToSUlCwfOAzP2Zlq
EXjmiEIJo8TLUvWDyWFza3Hqj3yALK9hRDQlb+n1reUNhc8nl/u8P/od5Rp92sg5xVng6/46M/9v
f+MnBZt5ijcugIowSJxoZrHBD9TLrXyqYyPXJJHpOsODskTH8+2Bb/kpbOuEJFHAklG5PHqYKf+/
rA2o55Fu9y+y7XRD7v2y5/RZjJUJQe3vxCSnQFa9wY4VxAfZdbLCCjuPilYjejT5cfkSVC9iFzef
xAKA1WWPptrhb9c7xRjEfMHgh8T/GcvQNUMeBc21VIV8s0sCqpqCOHuu0oZBzILybX6KfjHst/ft
lsK1ge5Z6gO3r5LqT0jVIyNz5UQpnHn620bcJ7NXNdBXmLS92L8qVYa51JvyVRFl/YwkuCRzFqKk
yH/wi0AMYu18pME+i+TlbkEf0ZywyvzKw5p/yprsOXI9c/Ez86yjFTC9AMLtSfISk5OnsR2BlkHu
5GPp4DAzE/utj2oLLZc7DSCCKDo4iTpYM4PRPUfZ5iJW3DCPx1q/J1I7krbWpIttMzEmlg1grQlJ
UzGuzE5ijRMgDhwDQULoOBN6ty3URtvS4OhfnmZXSmzsAKk6htQ8O3pHrpjN9d0+dcqmM/leSupj
w4i+qcI+uXHnlZDI1z+CioITatcQ+RJU4mTE5/SlQQEkxh/Din6Oot5iCokSmQ4Yw2KBC2eeAOPG
gcUzfGbx+R4MJst7Z27Z0HzGPVdyIIzFWnBo390oES7jQiPQbhBMUBh5upvMH6gX5CPhJV2uaA5L
FLp8HaF2sjjNoNUnG/ItYwWigAhmyvvn+iFSxyYKGuwrgOdbgNKLO97JnYHa9rNOB2CumdVU0kxO
oiUSuXPWCVNWci3Eh7VVfpaT4+h0b3zPxUQ6hvcKll1p7P+9brpDRSIdfITrAPPK4ONkpuviIPNW
4Hk5I5BEuSZLSgtg81YXavUzBUAwBEIBVO17V0ZZAG6EM/YgzeUt83/zxz+arss5+QzRANZ8zvPW
5XFHJff4E9SAItDWoPBLxUbdwCtUdTukQdg7is4DK+bpZ2QWJgrnR4H44VaSPJ+QOkQWJCOIuGYm
196z6rPkHiOFGeY8aNawRMw9ab521ou3Ad79ZjoIvv7q+ESxRrG+KN6lKRR3JtesIusXr7A3PJf+
SCHzk4lY6d91XMYFN3Gkx65wOCubIplW7AdlfEnqkXVg01WEZX2XZflflwDEf+6tJd5EYybr5Z61
Tv2SXAYMWHf0TQgfRVQSnHD4kN+bnFU2j6lfRGniD5hJ+D1sHkaa4NH3AEPno0OaBY0WphRzcMy7
IsEa5l6vZRtm1k2Ha5rdBlHtj0pF8TrAFrjWRJXiIQJDp/KK6ad/ZWUWdohJbzh5KB+8d/pMnxzz
1y4B+PQYzOl7vI+/0cOC9kuXTyLjNnc2ZnRtcuSm7vOwOWyOPhjBmHbm8YCv4xiTh/2pJJfOKDMh
bpVeGI3fJ6KCiPcarzuyxEW9aHwi8ZJ+Fy8XcbRN8ZREI7exPU9KA411ZU0PeWSUmrzSdSa4NJT+
SJV3OQTHIuvX6Kbk43kRne58RBFZwS0yxQoEIsF4AH3/5mgsE3YJ5BnoSkywDmcKBHmhJ0rQERXr
lyxIouXQK70nn5bGRJ1UkvQ/ssD7XqNyxjXv0pRQLbSGmrDkwczBOHuPDJSdru2vRuSBvYH8rMvr
ryGxyU5dS0AvWKq7tMrxHEPdOtFrdf6asLsXgqXlQpF6kC1pZWKbB4jJYmnUchFOwwcQVd9XGwnw
Jm8jv6xNnJNgnNcyhlxt7jKWCmS6Yj+thHkJDzWSpfvSk42hRCFY2UXarSwhkACBBVwi6ZKXL2ma
2QrCrR4nCZyLdwMyoLHYeMf6JAqVvQs1qsMZ8EsggnlFeXc4ShnMv3G9KZjVHQzAjmPx1Hn6UmMf
bZAr0os4BGsOtWlZBr3vQm/alxYHClj/+WpDlb1KOT8Q62tQCx24fHeiJKCdhBBLGSujWB2meyMN
JvIDqsLFmzdBOt6rFwHq2SBSD/YOi98xDd6TLCrjdZD6dbeJfl2R5QkWiGy6quHpRaw51xWKDtNK
ExrsJtv9FGLMbvv9lWQVXi6BkJ4CLYR8WgIyIMd2CsMN5Y4dO/V/vfMGliuOakB8vy6eKJwi90De
C8Ym+Uk3hvYN916w5wZ5YDsxZ8D6ChF//MWwHJsqgPFuXUpTxf+3Fl+6fFcLj/G9HfDBaCQ9YSmJ
sZpVSwrAzN3prCOWUGfFauzho2cQL8TJcS/OQgbQglTGIH2XtBobrK/k+N5hprxxpOFr5uscoNDz
iOb5e7Od5eHNQ4Y3OVe0ywPI+P9wdOI4TspGCSZ2GCVdJWHesJpiyDfiujUy6nBJi/seyYvP18QU
g60vlYY7XvB/yQhaORJrEuIVRT8B0kbS1xqyCFcckmLB2/GvjNZ9h3njplC0q/fQGtNkmYKRZGuQ
2bPVmo0CzzONzyQdf42bg4A42zOClrp19RixL1XpXv70oWY2VWARHrZRRHdvfKCqB6jCC3Ncrcet
dIBs+qpKbS3zPZJlDWF1ebLl2JtZVUJQvJ3T4RMt6FD62VYRB9Vc9SQEgYBEudgtBJlGbrqwx0v2
zzOi1VPC4Oq/7P30cyUCEQdl+hXbu9ioAGhwAiokhcYP3sMFE4xlig9H9mkjbZzqxmcXlAEtlCoA
Vqafx+nuNOzlqavBS+eyvWctTdrZo2aJZH+A+9uB2gOd0Bs3xCM/5ItM/CIOdsR3P0gCsAAU/Og2
9/afFWyeOjc4BvS72n+gZSkvmaYRi6euDABY0ZPQ0n2EaC3BO+L3yKN97LqTQQtv2JGwuCfck58W
MaiDx31htS70dVUvlpsOc+Y2f3ia29Y5JrxIKDWaqZ0AbPGojr3ytFDHeDxZFMI0YuxHFY0iAsAQ
sIoEaml3UVm2hQ7P9O1Fgk2BP4Cr9ndWV0CNvgFJdlTgx1NYtLozstmLz6KK1jzpuFNIEt3zLZbG
W3dTL6h2+TirYhA1yqd9Piq+k4cjYgzc9yKR6fWCgXF5h9kK+WcA9N4DBkImGAhFU6NHFJPwUMvK
9n2F9yfCKfb0PZ/qgU0TC1kol1DaZxVbRAcZ1ejY/Xkyn0RJt6gig+qJhqnrJfakpg08Aoxs5wBc
Zn62xfBDV1szhlQ+2f5RZdViNSKPwIDuv07rYU2i5yUdtfJCIkoA0Hpilu9B1w1xDjGcCwrR3rer
RSHguEyCBSj9sYBUujLgLc5mJYIBkEt403E+Xu8jySCLSmQDt653BI0RkEsILfYTz9f7WLf3J2c6
p4zo2iXvRhVluHnw6QX/jAg61nLReSkVqfA48/jF0huNwoKl2QlfjT0cBW5bBT60PV86FPFZHrcR
8oDzq4hfABRNYS1VKYoSlG4LgmjBUMApb2erI+y97MgqOYv0uEgF/gfQYgcuAeNKsHQb3ljTlT7g
4FNpkcZvPk9mNqDIDQzTZosbfdGqz7/KavNVBlLouMdGIdcQBjysEEHt20cl3yYr30QyzFULlHPH
qZubQZCDmFnw2QwXhbCYDoLFF5HjlJyPv2VGvEqEUVh9qnfharve06ZRgk89BSds5aTpDWbiVMO1
yGKsj3qupYOrGXqrd7lJAYZSsa6k3LGIR3iRKL8So2H/xHTCe82e73ucAfjt8CSeto6YGtfq1aOV
2wmDK6N6PAGtVOBa4nUfA7n6O5xxVYyFic8HJNAeXKjXK4nzxhJ+F6QFG5gTcJr3HfdYOw922+vX
OGCaySXOI+ITPmP9R67Y/WrqPE8tGmgMBJ4oW7iVWMuMaDRMIocE5t9O+HvyzF2I/23KPdJ+LVB0
0I/f6QrKpDJDLpQ3Iy2mFgORp2fy09wEW/lBIGRr2E3TzG+vtgWyevzz8PjtpahtfFer1dyjyH3a
Kw61pv5sMXpX5paKvDLGiUeeTRk+YiQgM9H7jdt4I3I2wiXB2XehUlmsGAFoN7zdskbEphhJF+vC
RnIJ1KZqjH7f3zPVUZEHLy5JgipJWqJYkg2bq74U91WE1U5+Gu26e4HVS70jbJG30hf+I3OpuH+K
4LAf81f/9omxlWHPK9A+EEgFqlPhCGXCtnpe6mClYQFlP4l9vKboBVD5r0/vSvgD68QSTnbOiHD5
NVts4KlAcEURyDakG/lsgx1mW8wgt88qRc8lyqw/KbivJHiTNjg7asPcu9ze+O5GRNB30C5My65w
da04i3JtQR+Dz7k77TrAaGKJPbdlb2LHVbm6PXa1oZMlzIQ9/OdO0r4pAgGwKTpTLC3sDgWeLdVN
M2lTAcQyHNypeOxRC5Mh7urPv9f/t+SeNG6lXSgOK8785vx/icSWAO61ddC+3N9+hy69kI73ljZa
x4tuivQbyY/M+K1ksxkQpwajcxo5TV+ki1KET0v/B7WVKb/4cmETyCpPnojkgXf7CopGnDMxSGua
/g//xz9pShcLtOPCb6cx/FEV11vNS38mrinlmdbs7n/r+WsFVRc1+nygdJ7QXlQw2jXXXC/S/rPo
3z3fe3uU+cFq5RTDMdv5xhdq3nOdTuCGMKz+w3lCxfE7ziku6C7Nl2n6rIgC9Ntkb8M6dgB+OGV5
RXJ/2u9iYjdWOC0E9lyYMheMGHhY5RMokg8pVPqxzSN6vzbTXIf7Xg8UOT1exeHQ+5sPUFs74rzu
27bemUo+SUQM5DJPGnOmCUSgpyNqzr/rn0WVNiDSjeSWSePGv3nqwYQTy6VAPIviPn13SPZGz7uS
MYVnRgF2NI83oLvhkNU70cjqJgSrmvcH4LwUOFgCQQaWEWRkpY3Pd3Pfw6v5z2rEaCuzr0KH8oRt
xdUhhsLD3uQ8slkV2Ea5ymkuoMknGVrun+hFyxBt3u9AZaBi56wH7c7x/Hlo/Q20nlJtUr/oJR7E
4F+l+McyRT3svhJikuGJs+ItZznk/zcgJVdVnHrD4OEBLQ9s2NDdSDtAtI6rdvuCAUO7JkBrz95r
hqSyG5RqmBrfGOJ1R4YwaOjMQ0H+OEXP7jwLXf/2FBvRoH1eD5hw/kDuY+illimR3lnmUqqfpp32
eCvkIsBq634q/fAvmvl23LGT4x60qlcJLT5Q82KCf/QeovitHeWX2tyBSS6y6Cxu6KpgTaQ4QS4E
nI9cK7w+e72FJUQMuOUfTiScxQlSD8Ehz5BZbRUgJnpHtKkios9gBEMiwK7zm6QrRlv2SKMhldql
XBDGYzyKDCeMllwO8mQKraFbWst1+z46todhaak1eUh4dpKBAMRHjYyoJg/TX7IyU1KGaMmfbAWq
a8hR/dwFsp7+YjVDw0cnmJtQaegploA4lH8vGFP0au73ohTe169E7NbQ5giE8WT7iLmbrNPMr+GV
PWoO6FVb5vFslfesAAbQ9n/VIUBQO35GwDs02g2rkydEsMOLfaOASMysyHbWKedb3QG3I6kZ+rey
k5pf/TKKT0LHgQTA/9VrmVkDJJnWKvzit468sCmY0lbqNRxptTX3RCHytBK4tYWRYAgLrbFTI1km
3laq4YuVJGvTtPksk8VwONDgKjttPKJN9qXa1tPYTeMBVSwlHe723D1oORqVib5IuYnHSuLsmxjc
UJDKLcpnUcOKA9xSPU425VnX98LqjnA7QWuRxmNf4LfIcwIj3UFNj+vC1GcdtNwhraUaCIe1Itf7
cUDmVin68F5pHHo8paSx8EmzSkjqZJDid8y3+NFfOKyObIWd/bSGu1ixQOTHGyJVJcLmLrFn6UKF
zYRDLPDAxr5gaC3iWwJaMJFL7lsSgFJGRXdC84a/4qbWbMUuEajQBp3Noy2e8uwagHUu256ws5vR
CKed5p9QmAKGXFx9nsoDLkydj0qbvRa04NoVCRiZRmeSjj9qkyLjyypzyXknKsVg6sGCa1S1YkmV
CcpScFVhs9lqKZfXpScGppzebIMlLOJaZZ0Po9nrOcd8DQyZdedf306eaDVVGnxIhbnd3xKYQwRJ
G9awEU1k7BzLYQ5vrRUItDmw8fAwB8yxF0ZBYAGHGoyBcll7sTZSrlZDBzXlAWa/qnX2XIANq/7q
jsaDv1dVdXXMT4N8UCJA7erg7TmQQnkEOfx7iXqIzeEXqLzUoRfXdIgaGB/77XdQBveB8UB6yxKy
UqICp3tU86dWYrn6bjks+U8+KbucvFtpokDjhDN3ovH9adMxAWu8ttdAeN9EPwJPVS9YZkos+iN9
SowBOlmkSCcp9McWCiXCE9PIf9pmDezaY78FcY4rqoTUnlVk4jHI5wOhymgNYDjmwRwIzL8EnB0t
1cbDxk9w47ooa0ajPK8zfYM+avHmsObibkh5Xh71Ms8stm0sGl0QEE4GvIe0tHaApFvHhYtjYtJu
rC1QMLYrZVHca4R7N4ilX2VNFWqUlrJeYspKvHwwwhpVLgqulhRLhbkZsSf0/hMA2jLog+aO41Af
bOJ2doftLutdkqL8crH4CIUgwIsmUTPsHwXLP2qYZXzNzeb63GlhtNU/uJqWFbj18AUfKPro/Tyt
ooKJEX0UPxgf7APTPVPU6a2TNuyLop152qPr+HL0qc56W33FoN7paDlt+e7uiB4m5YgEXnY3wFt8
sScwYMoueUFpFB9lQgSi+Sfpw2au2duEMEO44I7I0JhPjwY4/vcGAGs0/QWs3eLpp9954Lt6KAz3
wJSXgUeCKB8kfJBbGkeeDR3DRwuu8WT1giC5sceTbUt+17pWXnrZ3laltLEJRXRlxk1q62SgfYh0
+ErRSUqQec0fGd3F1e0nB3DTmYUHzqlEkN85VyNg/wJ6qtJ795bVPJcguq95rHuikCY2UxH48niK
DLBvV3JSjEiHfLJdjSpnmcPTtAf3dv9RapnRcoOTM6W8I7HSdy8COa9kKaucUFVTxVJ3V4Cno+Qi
YIQ5Ml6HBcMeRwM99AQLCZmfXPX/VYugELJjeRgn3zGjFdiUOS8FbVU+ShF9tXlxtRbKcX+izP2g
DYjrEXdqr9NSly/EUnc+S0qA9kzesADcl5HVc/16roWJ/B0g9ik0HZMzEfCseWynFQTmmB/0JuGH
7FkueWtMSWkmWqNXhV1f14WVzYD6lwyB1tARYPWoMh5Oz/49i+MsDP3Lsbx5lIQeZ60842Og+1eE
8kpgjwqMVLntr/YJIiHmZ5fXrL5RxbgCTgB6KurLJKbqbiN70YkNkybpX+vK+UUDZfkYxrKcWpn1
YgAv2uaOYLMVGp+PKttsSVUOXkXZNfl80Tha5vWG5hO6G0NgAUx3xTFk1nlwIld1fFtwYUcGHjnB
fw+nz25YE36orMt7YA8EAQPIjtmWTdYlvP1MOLjOu3xs5RTCQYbNBlqdSfMCsqpq6G2j2yxCzJV6
uUCPqtkoxnkoTQbSt81mtjb+UbIjKPDpI9yyINRAyDAc0zkUtbnrL+WZ0u2dvWXaaBNnlgfst4ai
HvesSoC3L8STAWHipDXi2SLY+rpsl3d4nHiCN2SxF3G850qSXDd4P3LXlGeh6otjk+FjyRV7wTEG
hz7uAmgmWNPM3Jdo29Qwx3WljFJpXld4JxHBAunFiDqr0Lx5VUo5c9T8dLvkF+63PkfiF3tu5iPu
sWj5gCiUizr4l5I/IAo+MEI27mDI9xxfV944Byjthrf9ckCt97sBYcsVwXei/DaQ7YC1X2qbsQMu
bQXfNK4Vwl0ajJL7VD2OpYSprYhJVbHCRfTIm3RgluA71vA6vrhVDx5hlcHH9Re7Y2JFAPqYR5oc
6ngFtTfxT2Wf2aL+s+aXzojPEGjIGEtfXEjt5lfc+gtsECXL6ks1cKqtQ/FVb669vDLTuIC51xQo
nUQhvX5PDnNIqymChgwdTQwZW0gJzp0bq34r+c1ZePvfUyMADxrKfY2DzAOT69I0tJTNpkiEb8c6
olb/qWHsYw6JAMgLsUa3RQhTEer340uQeYyt9sn06RXu+LMeMKXC4iB9vujdwSWKD7QYRqj2h4ya
GG2T5coUozfX39kX9gWullmEY1FFmu3uK9I6mMyzrGs/m5BcTF2dDC7WaevmSHGMix65+pKE9o9T
368MboYySTnInCaKpwoY8QI6w+ZyIBqGydMZZ5VB9eEwwPSjXF+K43Sk84d8dvOl+asJoOysF332
RnaMMqFdaTgIRxdGAj0Eg4cL4VbqgI9pibuk5t3+QcdZg8UpjNMFjCxfteAAcFxrblEDrn3m2Qjy
bGbNgK1J+CEO7lQ5RTJMJe57j8ZTtBnF0MwVNH7nRH6BbB3Y9sHa8A+GZ2LfJYfZG8OpPp27qrWD
AnPP7t81mvLM6v1g6WhF9TrUiuIXJ4zqnEpIDjVm+yDm11/agXx6+2xyhXJ3ccU+jhmhb/T/rkfK
M0Qtf1avjukDhTyNcUdEaQqkT80VWN1ANbflk7TY/g5agW1TAfChs0L+AhsEKoSJG/fzljoWRN8q
XFzJgnuPkhBTAbIhGw8rcKUxWDssqEf1bt3qiXX4m0jcwi/FuuT83QGn+142GHuLV/ZJ25KsORmJ
jPcqhH1yEnSKlelDm9ElKHhvTWPCn3/LtQ7c8CWZXYNBmE18MASlt069eL5Gk10tWfSe1kUa48AV
PyDp702yOhaCvZPOS6/y1NUgmWOH7HRDZ4iX7fwDEcNfHvlQWJIcNQWKKAmerUZkAkYPhX990KG0
+jypGwdTDutYP0huWCAMy/PZn9bwqgPAOEmKVkDObAYrpYLb7Pzr+dHSIoVL3tY06Sf5CLhbJynO
jTw6UFdEcH+aMD6KgaIE563+cz6vI/r5zBilR8jkyeFEwTuodGrCXjllQtJKTKjsT2D32wwOFoMo
OiWn5nHFnqKkpQnYPUQAgCNTzms5tCbT96fLxrjK0Td8MdKjCyzspMv++5xXHkOS/cPMR9zqMMIA
xAFEuwDqfLrHSyrntkT8Hodk8SSF7ZA21Pxihe/7OVJGpugzRUXsTAlIe7oH7WU+4jBuYVBYHeiA
NUfjw3k8LZW7rZ8+NCvqpKJ/PhbOdNJTowKOkl1JNXZK0CHa0ZFgHIHT9iT7IYJYfPDXMBFM3+eW
maeE9QueJeqNdYQrosWc0xLl2SPiD3B22e1IoKdG+h7eiRTS7KG42sPqbXnsPNgnMbGP2hGsWknI
EnI6M+Z++1/WUmohz1jgqty8jxzvMFBD3ISzCXapgu9KRWsZxtX1mh76a65XVtn5cevtTJYmfQvu
FdnbwZ9Gg0+TiNrUx1mlamgyZAZ9tgd8ZzMS29Z2ssy4/F5Al0t/GLPCbGVB/KaYfub++4khAUN+
C6tfettPbSrzFZtXn4jQnka5tlDZRmKRB+cw8oPb6YFkgMMrM96sVKv+X3Lv5VrueLQ0QywAEJE4
JTkBlLr94H/eIqHJcg4VrnqCb3PAGNFjqgYjMun94/frMRRzgHClCvAICqfPSAi6xgAh/2Eudm8W
46ZFxO/21LyiXBnYoUqqYSUXJoe9o/PRCWQFJvYIrc0+pNyS6+Y9M43xglVZCo0smb899IKHl6lX
hzj2hEw8NaLh6MuxMJBtC8EFyMREkvv+21GIP822I0KWRaGzrRPhGo4H2BVtSleOn/9eccA8u8xk
KN7swTGYoYBas+vYFOK52UCkAeA64A8PFmDt975EU2tcuHcRJqMB7d8S6a5jREKCutuymlirk/X6
PhWsIkd5Oh+CLFw2qi8+yQkH0WxDvLW68AGvc97ogh6hJLFYDahPsVdaERj77oVODDwiPS76jeDE
LPtAKf1yPfA5I0cz7juOBKGij2BxVQ21vxn2S2ypU7VCUgpXbMzijHYnWImMfrDknXCG6y+NF+9Y
x3t2LHuInxAA6q/lXVSWmdM7mYNjO221Fh3cDXft3Faw8fB5I6HvfP04hHV3tNQPt5tKCUnx/PYj
XMxwJq8r37XrogjgV2uBjvUf56IALM0gyDXe069gQtAwpHRdG2QLA4kp/aZa7JNbIlSqfsJ+82Ia
06SkJWkovYgmNV2+q5xk2mPTDxH0klUgcVJMf9GdcoHrwp9Z0R2EHTC/GWy4KByCn1ZZOeGt96w1
JQ270DpTXwh+ZnR1G5o47W2BwRfnG20g13Mrh4koaDUCZA+iEKMEcSG9PZAMuMhZr8jIYZzxQ6dX
eJ/oFMOYmuycb8fA04pA7BhtEeE8lz/KV563uV13Um6cv8D/BH3+S8YpmGdqawymCx8cqNLlOUxw
abmbVceyGBTfQ2kcas2YVvFz2TVLPy0QRoJfUN0KaPwHdqG2+RTPO5bBO01h8Z7F4UzKIEARpPcw
OIdx768ERnDVmRtPuiFl3PdBDNChGynFaoAdrLMhkIojBLshqqV79NXrVlnnoBcWrEsrBRIviuMF
8tSOOp3HAQnKH3yqcf+3BBlRGz5y3a+i+LbNIyc2TdIpzRNzz8WeN2vszeLmrf6kcsTFQKNcL1r9
QBsQK8sJm1Tojficg7MvyAIdnlZb6QQQYjfsbRZvhnebeH+hHQ8ETLHgUYPAF8TxRHKTlpBJu0Uu
Hhkh2Kw65zZf7ebJZfwnkn/m54bSylPwSwJx9smWxoNrqFHXdwgcagXMYi9LUmbsbThqC4ZYOkKt
wrBGXC+KiL5n8qpISw/rKC705H0mWTbf3VRWOX4QMiPaiKNgJbIg/TDHOMb3Coa0iI294/HFqc/b
6YnFW/4YGgPSCcbxmBYyqLUVUsbW7QxoXEIf10g90TCxic7ciCe0PXSLJ3i0zZxBwTvetbU+FSWs
zo4Bns/J7f/A339tB+WiGeXF7JUERr2ywaKQLGK1IbLytSfFLJrrbl7SsAUZ/WNEFesIP6naPga1
OWIyqVqfnm986AVpkJhBO7HJF50EEsb9mmB1FJhltmrHhT3UI8jtncjNtGPeZEuzLnKrOjt7cM/v
zZM4HQw/f4HKA+XExcBvW4phOhtEbSB7QdvpUMuoj0wF47CqGSjZ0PP9NcHdzCAf03UNwQ1XsZmL
QzYLbVipi+x2eTg31nVBM/x/K9KRksPT0F7+638s9Sw0yiGTy4fGdQ2FPmn72XC57CQdOIH9zD7Q
HfLDbpHV8lKZo6WIGmc8wFYSaLhrVApOJWwBxq7rbkTkstRdrjdr9VuRE6d6kVxUuOP90kWnwYoe
tL5tzmSbDZDXP1kUK2VcBxkR3eOI/E+8BRn8wi17NHmkKi0zgHQP9yW4Gim97ZhCOgBenv6smirW
7yrp5zG+7EiowWTqcJBFGVW+i1tv8ah0VBWb+Su/yD+llNcWMvWVaaXKR2d216T5l1DUPrtxcusG
5mBLqBLGHwDm8Wjk0kuaPJ/1f1bpb/ZKtivQ0xrt3F3wvWiMIxy1JzJ9p78HvIOhONp2Oj31hqAn
8Fwrr2DFd1EfGeymqPUFrwxPTLWEWxd2zyqEePwT1nPjyHCxT/WT67qEMa1D6MXohNbqWr5NHVVa
bO87Mo4jd0Hl6mZzUP0x/T0Pbwif8dyxpkXmD6jA3hOFeGsKMVTUe1sfrWM5qS8y4YyB2rNu5Js9
0XgM4jZZb+FrF0me6ZclDEVxsYK4pTDZ23AC6tyOZgySrpSq7ixIOVCLWfpvqDla/tyARsZ2PZqg
McOwEwMFh7esL7S32DiWImxAnybqfrcT++JLVyUR9NRCmvt2zIDvQMLg81UtEjtSs0NQl/L2kwO5
XAc9VjOe5BY4E4Pac+AVkjHTMgTVxrPr8KgQ8tpGy/+eE5Sak5aDBeA0kYcx/Il5xE919CoFHnmv
OUb4SpASj1/pYA0NQjujOS2j/UTG/vuJ35+YwRBRVkhOWiYgx2/t27YzRmyZKrVfOQkLFLzAl114
krZGqSOtAOoHMQA60Me/6iNWz8Le2zWl34R0af00+B3CXrpT7Pu5pBUWqC5iKEnB8j1HjUr17OjF
7cCWvjZnOYkOYpNaa5dNSaA0gGdX/MXAKo4flYk/ovGV7TFVXZ4cvnw+dHEi0tL0A7eHxmATQAIi
A9jo0ESYWBrSDfXcNohLPGlLNCmbUx2u912sYsIPl8THsFIM4oI5wBbEIevLYqTswz5LQCCSG0vD
sCN3HA3xjFz0NSODuqppi6BBbdIlxL3ETWMk8pPO/DBNByBAGoTj61WyZieMeoLKG+6SoMwTqVdq
FGq0d+wAb58tGkXNKAVB5NflMdxSsgiXpmeFG6W5xwU9eXUCuorPWBylRYQiqfVb2L7xYohClA9i
XLfbYhZOMHvICQnYSHgCYCbq+SV9dzMylYPqOfBtkU3fqlXdoqsVRKV6KAEJsngUth7H39tAtbEV
3iQ7VwvkmUKD1Kxu54P/ksDP2RUiKqLIIqLHjxUIsvTEIpgFffGUz96m2Bvtkm7NvhIXLB6G3GC0
z4lWZ5iCNPRjLwDZ1SjH2yfkBiTCkPzWOJEha9oeeMHT/51f2ZLrqi49pgr7WtWU0W65jA0wks5L
KgijvD2Be/N8pRrHzFYWvE7TGWV2gc3k0zz4fI1SBpyVo5CU5BiLMYTsq4sjr6cBD5dv1yYYSsen
7BW3Gpk8pSS7TL6P6Poby+cCPDA9IUCtnI7/0FodsxMrxhFgmwyVrPAvD7prSUuT2G9sprTcTehF
RCRHnsptn/fNrWLx5hgbNZrCGON+xi3isVutnDtqH7c2fpkqWVoKZ5DeKvRDldMqmhhg/SbnN033
KNQeEQsBPHWk8YLK1J+ULza5VuLgOPtu/+SKCA9XoWEokTo+obK9S0Sv+ZAss7Bagc+oSWEuJPI6
moZMRYbmlErsbyFsgHb7bU+ThTbb1Cd3lZce3eNHVhlhkjZOe/vgM4ed/5BHMQeuX/G/NoyePsnc
N/ClDYqwZOvgIxy5jqMBUReigdLTfHWfeoGORrlbGBLPQYYdQY5Gico9ErXjXOQNZkyDK1HvCmSn
3TuitsUjBcxIP02MGOezC/T10oMBoJwyc2sjT0VsF5PHqg6NdMS+HgPWydt/JFNTFEgUgrW2gddK
keeTMZdNdDCcOTo/TX185JiIoJSj17n9eKWtF/Sy473/+1sKpE2KetnXlAtkI+pqW2lb3t+VvO34
av8PnrhEUat+NxN2YHDQ1FZGorHWjHIPvE+0h6TcNJKcLkhB9KJ2D2oD2Aaj8Tghqfc263tHb9uR
aKz24GksgJ+6//jupU/sjsSnal2kCtVdH5/NJppleUmFayhC8Gokz8WN+FDYhIP/UXiByQq8VaIR
KAqwAjz7u9W0hKhH5BWWtPawpeyiQFXBViTnj19e7qQm2RFqhsltF964KRvVj0t0ZIoBN8Uo3UJy
FtKPbRJoSDSrD4iFRS7UKpr9BV0QWYBeAkoVofB5pZDKpzpoKmVZqUCzf/W7jBZVFlC1CcADcQ52
Au/E0nQWQ+1CXVaCp3eOjmwM61T3KIwK6o6z0c+j1HVGmQAIigmbjIN68j5NouFxP7yHNVXvPwDT
NSbdJW5o6X3ilMlnCcxGVL7MCTZ61cPcR62izByZRsvGBN8vEI5V+Na7SlE6pFwKqg7NDzbf56x8
V2Bjsl5ijABFPBuAzxcRlacWh3LYeWc5iN2aRb7Vhy1Vaykkttsu99PuZYP6ZAMyFQvh/YhkVAP2
O5wjzdSGqqM9am8OhYwedGnCKiI64dDjWJqNxbCBQlWjx7isM8/icYhRAnECCbAtqa8txR0rIO+5
QwB01DMBny0CK7hrBC1Ek3MnKMQ70txn6z7R4uVJAo3SxDOKjZqYFt6Vk4UJ6cLoQ7umSshqC5No
fDvVVvYIJW7ADS9aLxMzustZJEjSmFuSyT04dhWC+o4+uJRmHHfBaDsw0fpTsjLuWekrQ6Usrlcd
tzI94fgejisa/rNs3xr/6OCPSmYQrOo3JcqazvIjyGS6cpniZz7FJ5VSqQlANzc0GsetqGMu84/F
bi52MQh9yTJEy3TlSU5WIU3bgv3v4X309T6CoHJhRBvBzdA0v8upBD2mUG7zgRSlpU4XYl8NH253
roWOYHUfd87PZiiBRv5mCcx8BBwmVu0kHbLfzOPGVI4RgyH+cFL98hI3+qHop2oXgJTn4HIzI0OQ
iglooZOisl+r5p3/NJhBqhN0W/wqX7BGFwTNNbBb/NpOwDma8xcseG22QtZSrQvWdcCw13Q0WRSK
X6DNhV7NGht8GEeBvl/YFBuCir79VCG2W80Of19CNEYRuETWL1jR6X0e53VFLwLSq2E3KF2dHVkj
BlghVTcT+z9G5PermPUdxjrpSoeSfIN+ugBhFXvQ6jUho0Dsgt7SmzKj0XFN3faQybqf6AfkgA40
wsBkn8s3TH29eUfFyGgQ0xvlXDB6LlaAF/Db2X6zWrw9XZt9fHfUA2Yk6LoK679J+J+MkWMSUUA8
2D6Le9NtZkS/w5kecgXJcC32elQ5Pp5crTkZJenyHgjikRoU8I4HP3faN1GcowDLyELeS7y59SmD
0LcfOFbji0g+hk8bl7bFfUuHAwEEsWLiva6CEJTv4mH9tuIaGqINaQWRsQ6cj5OfnKkv6C0g7ai5
f9Z8Lb9iz2p8nzmksZhGinNUZPXdYAevTHP0E0z93c5FokLOFv6spjZmUuhv8ZoR7YvQW3ekFAYA
IIPuFO5XuGT5fSfgEahtnPJjNJnd2m9JIokmXu336nLSRSM4wFWtz+yOQecxumA4fXrbU7nEtLmb
K25HyZFjbQjnkAtXsHJ9tocNFTfXz9hLRE/469DbfOSPvgfRM0c+qxM8qkJobGgU6iWtXmslRtk0
6bIsaHz/LT/WdH8huFS5K375CG8vwo5GnRZDa5FdSuS0L3YgD8POb6V3el/9Lvzd6ky1zQa1ZyWV
dIdnwMwF93Oyceg8Qo6Nr4oYdPBAzMOUyGIMpV7e+c8YK/KmDU7hew9obVUxYG69wusjVe1d0gRY
YenrZ7/PRw9KTfhqGnK3AX/yg0RYbSuWjg7xEJJ0/QAXYRmmsp1rtca8BtRHmRE4+R4v/Tj6BPfe
HqnAe1znc79Mi35Zh8vgo7WvUvvZxqyfBmDkWSsZdRDNtrQ1FcEUD9VoXsC2idpGGAA2J/QHEL1n
o32nJ4TX13z8WtDwJOvYPDwWCNjIkH5BYKEq/pj1S5eTV+RwBei0lrgVX0JVPbjBleN1SdtU4McO
OyycPRc65rfailfXeiZ6sS+CeOgllbBQnOxn9guVDvSCzPF3TEGq0DbZPsdNcH1/Gy2/880aaVGP
6Zat7MicyfkyA0GDTSnAX5sKoza9gpBaLMmq1Zimr+IzzCIKCEaGgkpm0CtYQxJZkPN5KPGMcecr
hc3psSWomPe2jyXMXBqc9FINdOB2E4t8/RbaYyDFV8eGxFamJA3jQAsLGhMIk82+VoCy+xwG1Ujt
F/F1sY4zYVJG0KFsmkstepOPSwwyPmCqTnw98M2JEUEOSQio1D/OCwPv3DG+qkZyYJz+sw3qYuSf
6+xKZa3XQWEcFEmy29qC8MhGm7EF0w/lDLA9r7vdA+7FnrWiN69kQDbI+FP4HKAt4gR3QRf7grrz
93TV8F6g0r6dVr7cJQ09ibJG/xukpMU7d4WBR5phdkLuf6KlyLhXQxA5w6WULeahNhl0H1htWep1
J34m1JcEHikg8vTp4zECOvCelAygodM4suISRT0izXeKlzWsKNPQjTBRdHikbEQg6Y7M9cAOlu4I
/oy/Lc6x+ITbaexUtYCs/ia4y4VyKMceIHj+ZcgQrYpxQDWBPmgSe+ulwxIhmbghvVSken2g5XPw
ZOkEVvt9yQfW4XorZ5oaaNZyLQ4RHxgy65il0LlyhQex8dvwe7Suad1F01MJxAwxqYJyfooU/hwV
YOFZXI4hJRXFllY5BZZTIzkJiKsP5Iwk8XaOaou1C7uJmbFaRSHjYoaQB1jGMBIiwPkva4a0HMmu
q6Vu0rNVT0p5FWRA2MhTd2y+DD/gMaS4GpY5YyxntM36wredUM7RR6l35Slt3Y67i/8Bnos/oA8b
0OSwyMVQ0sOKBsFSW8hsDLlaIxSyrTYphcbo6afRNzY85aMVQ+NU1woyOchSz86+ui6WPYlKSzvX
Sfi+OJfQnNY2aIazg1RgmQsmr1MmmdFkfetUR1x5Vx64lrpB3s6B0ICD6TSLQP+uqiHMUMqX/3JT
Wqd1/8eFr5Lchd5sk25WQGBudbGT9NDAtmi85mzrXmBuW8AiP2j6GXTwU/znAFWODI63MMJ9TRwp
n+BHpRBwgKcFdFqUh0qi/RbCrzVbnEWaQYTicrks1ITdHs5zvXWtmsOasWsH+hy5YXZlDFkP2fg/
WxKttEgDMBKBji1ZfYRZqoAsFQUzi951g1cSHliey85KBKIrcT9OejXY08IDJSVBQ8iRydvMp4OS
rhLUVREqbC2vqPO52MaFFLuZuCSq0j/J+6sBWC8TvoaDQbKYP4c9o6xmKyzomhxowjt68YOI/FSx
5Bhw/i6nImjfuelUq/YUukPrvxEcKh/QnDl08+5di52F11gUWeTfELMtVyj63Vppn73U1XVSSWH7
CGOfBk02CWQYzrsYGrsTyz45kpZf9XUhluG54F5RL+YboxXfdmQc2EjlpF6n4p49kEnH0UPdUq2y
wGZeNLgkX1e695knG3BRAjwSzHJzy/kf7QeT4UXhSQlKzypnN43rIq1umcqJ2722d5kCNS8pWkRm
uwmTFhFQa9aqaS+pcUt+f/NE5wXHML3ALR4ZNm+sC5ag4c8jnhpwFNrqPxiA8WcJ1on/zxzInp87
pkl7Jp6YkLPhc2Yg+HpIEKyN1R/S1HuuqVLMXUj+zDWk88r+43gGi6+xVqK8lsDt54fraOVsYXp4
rd3zCcsLnzjQMFKGELsG4cQjN8jERNknEP4RixmfeKfoV6dyn76+KFSgBRDQE1RR0VWYScBV+x2G
BrEpjq+QY1naoAvM8YMuRKyZSLfkAnC50fCH/n3driIxgawKKfdYtTbZClZX+lNlDy5AS+SVUNJR
E03kNuSKYMqkgUcTvJlVVSxQZqtxCLZcfO6RuXHWU2eR3vGoroWPLYCBw2QHlbeaqzO1XcGlshal
bWYdNLZLWf9ithrRurjIarm2UoOJp4nZ8FJhw/J8ilnXRKbHO/hMvFmIXkn/OZ4moaHgCtAwMTeH
lAeSubv1EofhMvy8RS+SN1jPk7VgGR9rntDxmlmBR3ogUy+SKcASlgcynNuOfkqhVE3iGgfn//Db
vhd78j+EOEu8WxqLcqS+MHugd8Qt75Rx3o5uvhiWJOQfOCJxOePxfrRzS8sYpra0eQbUDHPuEUYi
+GMDPKLPPo+iCwmoj0ruozrs9O6EuPscz1NkpVjLsHWc98gpkylx4CIbTRoE0l5ooI1E6Mi6P8h9
wQKkiXoTcFiQUhMW3dmKkeLtwQpYWnHvewfqqpdvH46Hl1NzLYrbWifrqKw/wrTRgCUPlGqTsYz1
RqFuR/xWkp9AcOsg6rHi6F3gH+W/aYCziAIhySgYci96LIXH4eu7BYLB88IydFgqeejl6GqB4vW3
I/7lGVeVlTCainq+KTAC38qzQ7NRn631l8xvAI7QHz3MCRqM+nQrLUlV3oaRSS1FQ4ZUFcETNWeW
RonCOJmpzqwvdyYXWt7zJwzDdUuVMntyX9UN7SS2+jJeUku0FtPxUcviu224wWcn8NDt2FYpWuQt
R9O9FZjjXrRz8Em4uA2OZbokTntvbp7bTrkQZ1WNkisUkcc+RDlmTmSsVCiKMs3qzDk37pPNkDE/
9vC2hWwTudms1dYSpe1+/bqcn6GMnc/Ld31zZOUG5T6z8Abwy8foviRzVQ41fNPgqu33BE9qhLOm
DqfOGcWQNy9fkoa6HXtmeI90GWdeeQPXcZAic0cKjhalC3jVq2M0BdSYAlvURlX0aw4IuKuFOWfX
KiQr/DTpcik5yNmRbKdXxjdj+0IPWTjT325unhR0Z9sDWmIROtvG43paPAWjuKOn/m3LUap8Dm2g
g+Ac1knBedfjUYBihA+CM+1mv0q3ZfyPqFuohD3hfMjhe2ifKWFoB2BT79CaIAdOGrBGd7v5MWCf
7fi3zxWcbbM8yN2s/1lfda2bEMPRZ1BBxVYLaQP9FN6aYVCVxvrPFqJazoQSj+gFrl8N2W6Faudy
h32uLv+gYo8p+bF9Rsn0E9HXH20uy6+is3p9C/pX2JC3Dm+OFt6aZVDtsZsD1NoquGQvOWgdzf9o
bJYogWNXKKhIWCviTN08p3k90noJSQP92gEpHpPUoPKoRi5sjHBZzKJffnWzUSuj7gLxw3h+GI4o
5XO0ZAc9z6gKQUmvNeSWWLtpBwfqyyqKX+DJeOHWCSSFY3znKmi/Hjeot9bmunGbirmJHzI3xwRt
U7IzxEYrj50DWqlZymL+G73/7B7pRhAooRd9suv9+gUDMLuIR7/ctbz/OyWAIuJdoVznERwYzmGk
lVyMK0xyJXbLtFlUgoumE266XvLs9IHNWtQ7UUx/JCoQhJ1xgKeKhRgTNb9WmTHCc+ZAGW/4ytkw
ime5aTRBiU5OsTyqY0O8xTTntAl2wOQs/vj5QLO0JvB9HK0uF8S8aevffpDYTIHIdxGq1sucEVe1
KLzjW7uODnKcgzjrivZPzKcDoT9lLFzM9RltAqKn4KOTP1Sabo9lx8trclUr/wgxr485msDkcPLH
UXQJQCDDvAMzzvSzk8y4nNNYhN//8K31iTi2Q+QJt4IEy+jfzIu4d7g0APT75KJgVUaKaGdLw8lo
Waovi/HELwTcLplNA/m3QncrBWZ5a4rBOl7f+blyVBgRtqn59jmk9YimZbv6nM3QxHUNJluPY7XH
Uyjn9eRJK8PQw9pb57Is/etSfqof1KtUMpajljkiqosXIiZqyF3C5FfmEKCnCWcga0UmSRpMFzWR
OR/Ii818opOHXsUxKL1bpnTq91bG/t2NKMTeaJu6zjv8WIZ08+3VSyIyC+0KJgwFAm2t18p0WMOs
vRMTvRxnVIrZe/1zvFr7RXO5PYlEpkquanJH8wdApJLBxmMwb4fXvc/3HmH0eLi2I9BDNDhaqJqc
PTIP25j6Nn2S8o/3Bq5P3hhtN2dSYVzS7hpFADW4wnddslWcBOVZ5jVfkpTPxLpiGfOY9kf+ic9V
0C5tc2/ExIkjIYPhFvSIv/HTVgR0XdOvDfldKGOxKF8Yj8s0O93sVML3gIFwsvzT28plnZzNAypm
HuDWQZcXJL8P7w/v+v65gIxaMTtQXeEAS+Dl1fsISDBRVdWQEjJE/kSXFaaK13dZmGt6RLHhBZ4z
YRGgf+kcmAxEOp00duiorNzVdWpwlZKB9PgcsmtmucZ3NfC0NZe4RYZ8uEvao05iwf9/AVoot8bS
aEAo+KLC7lbrHA1CWiflr8eQjtstDksjrlI14u+Cl79SdLbkQrW8sPBHjntjgeHfVHcwYtRUCM0N
2bTMJkpuQTMpmdBZQIpkfZVRJ+mfA4Z6oqxJKT05vyzvpCOHqy2G/12G8UIuG1Pf0RuTB4tjV/yF
oUmLGwUUlvIYoB59sCNcUmH+qpQMkA1rkjL2/ZQc3s3utnxd2P+FuCiQNn5WFtBRBqtaFD5ngjOx
6bqU6Ph6nRzpeLdAJ00tPwOShYYidHC50ODqgUUsZ+DIs1opNKHLgpwpC1XY64yuyHiqDEbVYL0P
e3DccAwZseFKldQLW5m5E9qxfySn8/GEV6etKlKCHYBiGMHw9GVAsfjW9uvQpM9O0Q2c24taUM60
cFwOq1znVLnHhmlf8eFEwRelRTeQeub1vUlWAeq8AGH5E7IVPNzvBEPbIMcqxqiLY5RfFK1witxe
v4VUY0ik0FbNdMz76BLLHY6IBWmwgCQ6w9CWkrnz0+hwtbcTdABDz+NXMb/8dO8m6Ppa/1ofDLIM
+KA89LDhvDPJhmK/1G97yv5J8NlUG74W2FHMF35uowcy5B5l11VSqCqJjsrOhFaB5ELoeKIUe/Ra
1ExFKk+xnMKF0imbgQ5yhfiFmvguUJ2hyDLHo2aBQVn6l4jXSOlCc//nFnEXo3MWzoxMEcYxxmk6
KusAEfoyx9Lrzdfw5sDkBqzMBiaEBOv8B97r0Oehr9LUx3Mete3gt1ErAZ6OdkZdtMcBJaZM9UkN
8N/Bf97Vsj6ewXahJeZD//ub/7HzRMi4UxCvs/KUCWIwROGYXGGRVO/ffUN4Lkp2Sf74wQu/9Lf0
kGKTc9jrdU2PPnBhwGulCweSP7pOXkYH1FxfCqnkvOivzGgxqrNWqCdTdmlkac+0j39JTp8BD+r8
oas742qVXXlAgxcBffokeJlxo4TFYgJEYJhbw3eFtS5SBjSCKMPUrJflvirpWjPWjyYGiBAOelyL
aVKDL81/R6N9yxOOw3bWq8hUUT8E9akS924wJQmRsNb+Ql6bdMZVYiX6vHHLoObO/drC9pEjpr4j
p3BGvMqlNqK+EPwrWQcug2VIZhzLDkF7CA3FlzA1QGApSdfEpJCugnNzRM0QyP4St3NShyJfjNIX
N5cvvubLxYpnhagA9aPuasDC+ZaI8lmUTqSwRTmhClym+fIxXAowz6IualGBnq26OGaMikqmVKX9
Q4mIkFb/OykCuwMINwFguI2dXdlE9XNIVWiKpt/PMsoa8/TPgPytjMl61ux8PpHcvgZvm89LsgW2
RhtN6vtC1PT83Xb5BUstMNFstmggwlSk1p6HWNokPM3ORR6DP8AkwESC1DKoPxcivL7o80CwBefe
iD4u4ez036VPm+SHA/t3IVhG29eihqJujwWk/xm4KmNdkDXb+YB1wm+UUmou+uZWk1K+4ZcAy66P
j7cjMMDPCqYsQ3QNb0U4yKh+2nw5zuFYvSqSam52DJQbFo6JA98hIhFVC/Dp+2s0IBLP59I3yheL
tCkL+FWfvDEDTAXfvPYMTrjijz3/2Sq54Yqi4KG4fOd/srtN+zVQL6V5cNAkz6xcXg6f/wJ5TDk2
FJkL+mf+HlImZvNEGxICx03AkzZa+xoCpTSunUD6yVsvo+RRZZfMQH32XTtPnVCOvQthRl76hP/k
OLlsFsxU1mAgGfgsbcXb8rFFNzGZMbpMDBI4Eqkn6GB1lIY2x53yxcQRj8lVHvWsJuM6GJ5oEoG2
eDess84zohHqgsxJvNmZ4/8EMUnWpcM0H+hJKMqptuMcEk9G9McMciO+0pfyYzjeaqa6y4Vj/uKz
EeWCOb/IvkyUdzWGP7knCg3xl6L8e6vepgjXT/PGa5PaHu34aXtjJWkKuKVumSrTQ7SBHFVx+0nK
bjALOzaW+lVpMyeGvD4loRKMGXd0BzdY8U3AnxD/uEHs9UqFcYOcl8GaS95sbKlOfhzZTzLqijKb
HZMi+fGnF7JM9A5k8ffLb0jVHbBogEjpKOJ9EQyS98L/3xYOzfO7ZHK2KSVyKB/O/aPkxoU4JECf
x3YhTPt7LuwpsHY1Zpfg8IXplyNP18soJOHYTG+sl70dwoP0/Jmtt5PfW0YhEf59d+PGJNKF38A/
dfSrzkoJuoZ8NRQs6cQ4wi7/B6W10cttAKGk2QRw9FFJImWx4e1dpEQu/H9t4J1L3f55UbCrcOT+
085yHEBWGTnQ/VUiP8oTeyVcQc1DYp4kV8JoFrYbt09XY7u/wDyZF3fAo3Kzebj2rbm7GqA+3jhb
Mqsv3uodnTGNPi0Ru2dGL2Z7TzHVgAu23D6C2S+tijPhEoe8gYubtkZxMyLBhiMZ6o1TvMQq63ks
elw10j35wmdMFwTHhM83roOkj0Wdmz4fkJlll4l5N5rwEu1xR0mXyZ7MR+Enjc71HCaCWALL1f0o
Cv5i71kn3CIkoeTEqs515VSZRnvfinHaLZLW4/HXqwSW3hDUOwbEI3vp35gtLgweKq7NbgplG2wY
w1SIPPaBGX/043C/a1VTkB1Lr4JzSzda2DTMx/QEc6peywfGUwEWqcguRsieiEOUOUYQMPOYHxHq
YuvwdtBHaPOF2+w+U6hjXZb35unj+OCX1eoH5/Z7i+gTyFoqRZQNkuxbhehpoThlG21WCCmqrhfq
e/9FYQBHrI/rg1PVyC/pEyCxSaMeRu1S3s7aKGBVp46Y1Ko14/swZgO+gE/2k20rWZx8V/y25BWe
BkX5ntECHLz5EPK6Ja0Yxuw2rJ2JNcU5fOceWbqDYaVh0spaMiGJ3kg2FW3OFq7wJzgL3/WRMYfT
dOd72T75aZz6iQ1AyrY/gfWW3Yjn+DIgveUWBut/lTERUobUjLi16EiKjeCXBwVtwbVtnNbX1jpw
OdzzZU/+7W7RFvEOULBUbTWxDCHGcTIEXDTQDk9uXOvMj1/fmBSYDOXGKZf0t1+up9AL0a33rX+B
EJfT31upXlSIv/PMRO3uNU+tb2VZnt2M8WZbPgOqMl9dYLdo7M8oCx+9mr8JY7ODsZ81zkBab0tb
cp7yHBeKYGZjFO+NdVuN26ACm2RD8Ze2WCOmfi4Q0wF1GhxCOlpvwvKKcF1h+RAyaVCtzS+18V8d
RW67Amwd2F8m4Khl4uaHQaACzWVMQnDquPPUSZ9nmjGKa7r+8u82uIS0dGI4jPlBvrqG84geK6zO
B06HyhjdqILsaIEpeOwQh9ifKfqKqg3LqhR3fJvZ4BI9ilGOwd8IbsupRKa1wxiFGpRzhg4djrjU
QKiT1uGuTE2/2wjFl3l+nH5l8B105vtMZoi4OLIbqcUca9DESU9ltHSSykYUZpLseRdKkzrR8k1h
ZQNtPGP/3WOJtK1GtboXkXVyTTO84iG2DwK/7YnQHq1/Ncs5fOPgGCZ5WLA2LAf8DxjgYvI22MfC
MjEw/THFPCoYcw8frJeBAWRMq1n4nG+qcuwIum6GwGRxUk5Gj6lEwlnMSxVVxYIB7jRlYWRT1e9M
pnoCB7IKo5mYSqijjYruaoUUTpiYphZ8alL3RF0POZ4G8IZiYwsRTAOVs4yn2eJV+WxkGhpshTaa
3iBED2hDwRZYCxk+icDK/2WjH8GdUagzk1VV2Q45bKS8QCzvYAG2qEaOamRLbxfD4gW025NbEo4U
f30G3LtDtvebtexp9cG/RDTNam/t8FROIbrzcwUuuXMKKyfBvUuOVKc0x1zSFI0M2xg0s+rfVJEa
XCZWTW+7/xRnFd3Wkcrf8G8UmT+Xv1hlRtay4PweW1Ec6nOYUupZ0+178SOGoHRhn2DCSDA/G33P
fhLCKsy9y7LEwpnG8HrrBmjUygLUSEhrZcXErF/LfS+3wL690lsSr60B0wogQcS7Lm9sqEB/eRu4
gYcaAkzBa83SHnIPrWBUY0afwenIwdA+W3p6pSNWgD1mRXfWrAB3ieEbgFNNQ/bWVVHZhoLfcXw6
jrTsFJndgMlnDf+ciYHuclQuYRsFNPE3rJ84wqbK7gho/kvgEon9FzrvSK/KJdd/rRtjtsmSYmD8
bra6iK/V1X1bUwAzTEd6HbwdJUBnoQ+CA4eAX61G7LAJu/dD7J40GCU04mveXkrXfOTWXk1glzAb
L/GY6c7D/FUAyHgL1tOBlTT9niix5CWyB4iUGeXt4njdk/YoHaPZCrKUhH0nWx6x/NBgA0IaCVez
YlhthRZa34QHFl/v2NgLdDfln3Vkg8nYLUswy7VTRb1BTwYQRuXiRXmPsXFx+PSimIexg3Rzz4HP
WRjs+7xs9JifnUZbXWtEPqENyLPF9u3+ZC7byOeLvDUOuAhZpZ5MLj206lsXHOymPFqQRstp0mkA
+kcyscxn4mHlb+UnbvaUdjNkllXnf6MkoTL+qSzZdcfCGloWS3TJcFtI+fisxFLJIWAfeyPvvndk
+VZESKlyEyPFbEUcej2MWttBm9P/SoBXm3NHSUAiRoWD87/y45dtzNJcxAidjJTgiLHC9LpSpIvR
cVT/FexI0TXN1fq0bGETN/jA2xVRmjg5opv2sJOwTAX+jNetdqO2nDfOB+mYOya8w0cu2uRfx3bN
0m4FXUVpbgThWM9RQB3QWEyavIH28mbhXczbUyV8vYb7a0Crfd6S5e0olPQF6Igdh/inOk+1ojjl
DDmbUNVYty7y/KuHcxoNx1AcaW6MnROsKXUjNPOAnV9nWCdLblCIF2qrso2/7PoXANy+eX2QNGlm
aIovQhhd7CRjqk+dPw0P6Z9f4E2y3Xhs44asYbyHxYmh2W5/EUriS2YQAfal1FCpt9D+wW3telHR
38uF25PEbn6mF82UV3w4j5Eaidk7Cy8CLh73Kqzw0Ogx7rTAwo1IUck5csYUcFwrg0CGG5OZRkw9
NRHjsCKk9sfARi7DTZNR0yedRkOG4bXphsisiIAp2kXTRiQW+np9Py+odwEI18B/GGhzn2IJxYX9
7UWojoAJXAP8kMtNEA5iXhGrL0J57iYUz/m/r0BBWVKiMSHTbj2nokfhM7r3zZ5h4YrL/aonaB9m
4WBQNqZ7g0U3Zrn4xS1Kxc7Un6IXWTZ21EYOmMiWLz7s0m6a9FU/BmgF7NlAXrlfCtcd8gvSgLO1
mUv0JgIv7aKLsrC/9BNt89bx0epic3eWQlYKfnObkTWolsgqLlidG/czMgXUOaFfngio63R/XPp9
TMLmBmGZFF5vaAQbLOlMav2ZxMVUA3ySJepPsQdwSQCMYHdMM8l3MmG41EIkRYnHlxfUXZMRP/Qj
rTefuzZ8UbyUcrhzo6jABars++HcEyUdP9T6Cn8T6QnU5kMRXlsCPWu7aBoLmOZo1SQZEsbk+D7f
NPMTKe7eWo8TYdexqyrDVlUPg8MNQB4r4/vdayweI/tRsRjoA4W1Kdmz7PXtbqRPyb1HAB+BIqNf
51vvy6y7YAfIIqNCZTSlnDnu66AERZJ6ct2xk0mGE4dn2761UWixgaP6AVbsn/86dd5Nxitk/1vF
1IfJt8lqpbQJVqHobK9DfufKCLnl02duuklKj3D3mHhYZM21nkWMwTYHKm84V1ZCFewKitCJ52K+
pwZG6Ew04DqfyPpePv6Uy+y88UzY3Og3EoXyWPEOxTkCGosRUmf5755KnS01UQvFOedaLmSh0Y8W
77BR1r5n+OyD1CkvM6+Or+8FHkpgfhv8MShhaivr+An4V1h68/5qoKORxqbcgRX1UbyIG+gbJXOh
l/LHU9ApB1FdsaZKlSlW4JQ+DqDysjDjY14NFkfXF1fXBgkjnwY0A8XYP1BLucavFPQ3A1Bjgla5
FPvV92qyRunzjh6x0p4Sg61p2ZPKgZoIJHTu2OyK6lEy3mnrVC1vUkuG734tFEIPCv3zdDZAqMIR
AU3ByAdrU10CSAzVU5MfBlk5kw97c0YIkuSj3u6BF9fnYgGne4C3KDuKMYp04EtA58CJmPWjwz+N
dD1hdnJHN/fYWoF/Q/HvAe4S8F7/Fi5lETcIEwNaftrDztPZ892vzTcHVUD++A5Fp68V/VhXLuXG
Jlio50yRjZYDosSIHAyBgvb5je6h66rkOU+wZCP6MZ8DnPNQlSmP/PABrccBGNNdlfvI3o3UwI5y
CVPwWuEMRoA10VU/Wo0yqet4qWhnChfvHSzjXio7XdrNGOjm9UG98MNHYNOaY6hhAPvjIjXk3w3u
VoOETJaN05fOFDKAhY+cw8zfN/STe1uTyaZq9LUnVxpA5HKoL44UMopsZLU+VryM8qNUem240yci
cudYXQkxpsuNfTLTc8WEhiWCPA8ba0+sENsN2smOVOV67vn8JQhwDNDDOJ7pIQZdivT6+x0As4ed
dCSJhQ734hxqMt9x+CzClVfngEswhzYhuzkFXn9AroAPKzDYe6NQqU3KrBGKtoQBSn6UmgLhZXea
5gtaKMHZ8b3Iq6DC5XzWOhRzOVxWqL4NnV+VlSdR0Xy8xsf6S54X5smQzHNTpX7XQQEFsw3ndLJm
ndplF6TQEf+2kWVu8Iro5JRktX0ozETkSAmxQEUUhuOj/jd1uIdnROAUHOn55LZtJdknzEAvAAaq
U20wJHtwIwzXw5AJB4Q8GBISXhXjCa6DvQ++1don96FbNJtoYrmM+JDzrzKE2hFl3tTRbFhuZKed
02HkCAZ1GKdIUB2kIz/pVBCrRwb9PjHB3E6IJMWN/tUU5LC/JLa9OXIhQ1gZ31fGPkNiufZeHtQv
fBT4DfLER2FMxkwyUaKSn2zNe256+eIlGahevBZ8fQlMczcVMDHjt5IJLQw7g7/mk8zfuJaGNNP8
7vSxFtPDfBFKe14hfF9P0rZE/2ZaVsS1n8HzzrKHNDcQW7J8XLQUUlqt4Fz1yAS6AJR9uQzVpyzg
xB4PTI4UdjwWaEn6HsEdbsdpe2hz4whwSAQDzFG/A8/qdgIr54TDPWm519/1c0UmBrSUYrT9iIj8
z6TfYuLSV5iOHhG5LEhjXLJCjygdQEECVJEugKWwqBa6s2aT8O5jSHGBPmVx68SAkFuVuWJfIwZp
N7dRJg+rjIbxfy0Hv4jzS4jY3Z4TlTbsdr+4JH/orA8GDbebCa+y9JPGxR+9VzXGOlLT9v9Xet8n
ucLtDoXFkQTk7y4L7k2ZJWO7NfwHEB30+hcORwEAD/fWZd42wg60yC6RH1KrJZ/NJ/IqI4tDkYiO
WgYc59ZrBo3G6mDJLNeQM2CzyUzFtlLA6qOwpudsMjKFOwM3lgA5Noyj82/63QNXN116h0LicEyG
0Ck0bEUzUrZfJjSv9xK7Zo8t45TXH52pe9XAKAqW56pftuHqtYNph/qbPNNp+latK+TgIR4/9wbM
7MOwrs58SzqrLEwAEYoPS2Y0IC2V3o9BGciMSDHSAJySofhX/URWRQdACH7WQSF4idX6TOYWyR95
TO/+UKftqmOoFJguU9OsKBnrNorvnuqAA+h7ltGQYpvUsRDAlv9EFAdEkoKBNkEbVoOMNr5s9dx4
aSMhFqFifj5L4GeVcOtFiQ2Y68pUyd+9unU6FpFexFtZFRDTDBm+7AcJBFEOp+BHETOL48ZBnm8v
fLWX+U0VplOm93u9Z/v+3/2tFmCX0GYHlR2QNzI4/xIojHzELnPsbbR6qPszqOjqNhlnRmVcztck
OQXOQZ/DADZ8RJF6FMVvpyV14VJLs5wDMJXOwVlLhkyVAnckKkAIY0hY4SQMO85f+zmtgJQ99RGA
5et9HKriAmqJZ1fHP+p+tF3uuUZSJFJx/X0jL/hSIswel8Sm8+IiLX7a6SYsP3UM8SihCtZhL+x3
ikHsr++diYnEPer0eUfm47vNjG3hdtzJ0g9gjvMoxqZHXdMb2wcJPhNJ++VX1OWDoYzcJ/ZPf/yP
pN6qUvXNZ/A4u+CWnU/Sw7yPqdKW3LqMgp+qWaTdMWpgqymsFC/EZBRHVeifbzXjeCutbywx9US4
dfGr5RU4FjnqvY8BHsb9Ab2NicVKWNu0jB+mzrmdHTbBLtp2mxQ+7QgT0WYFpvyZ/1yl9dPqFiHl
ZHjbyDpn3lFdlmR+kXCanhbSZkh6GFrucYyCbaJIqJt5YhX4GF8NUUg4mbq7lUDDWRlfYgZ/3Xec
nF+QwGIvK2yGUd/3lJFPtgDotdGEI2lo0WdWxES7IrrC1pZcuq1cnaSNMGU0cnzjyIFRhG5+AOLD
+9n6BxWbFu+knhUYQK3Wtif+LhoDdUfDNn97p3CWyOLOMn1umIXSnEmn/xrwuDvsnF784Cxa49Vo
d5NFvCvMpP4irUci/0HBNDihqJWgI+SNeeMqLqxFHBxnlJxJul1N9u+eoQPM/Ef0DxI7KHu02D5L
6pEcN1F0eaSonBz23GeLnN91liwdJpl63+u9M/8+D1aEDYhjQA+OE5Fsyqjb4R2qW6lhg+uAbq4V
biz/PltSPyoX8xQsDTkOIETasNU5MPmDVrjIWn0mRyoJTsMCJKHYUF04kgLcnJAIoHuZL85ApFYs
xQNtY61AkLD7jDV/lIbBVJxMTv127u/S11DANk92GT35hV2b+iw7BV3Ydc49/UCW682l70VEK1Rs
II5pjT6E8kIGcN8yQ4buHn8PZXXwPD9GB+lr1x9Oe8NeF/KeA1hbanvV3htki9V2neDSQTm1iwfw
P34S6C0PedBWddUkPxfEUnkhapjuw1CMnfd6BYGxHgP94c6aLVCq/vhhZ/5bmR4yRgHvEN9cXY3c
gZEaQiZXOJp5mnTITbu6cQyLh7rcuBN3U74Z6LpXmo7ZXm2RN3tsLfS1hAAv6E6ABKNI37Y418mC
1JQd7zURTVQ/n9rm7bVqzcBnxrybvLSNzI9FTMMim37+r4y0DhNFuveu171WJuQZyms0+2VIwzqN
VTC3INYdQOexlUrAdSfeUp4vQEDT8/PgJ8m5pjy78oWBRprNnUygri7FaJ5Ycnn7yJuWQlZbEqRt
WurGoQvyj6VlPDl6qjTW5t9FDSke+Dbh2wtzyfojdn6I1uctAqkft/CCUN2Rm/LHvPB1P/5PksVU
jOkdl/+GpHvZeTZTgwuFKTwCnHCCYMya1aLibHU3qktyDlK7FnEWYJa8jzdVTFiDNjbD3uXBEvdF
aIe5GCu/U29w5hONVFfa3oXqyBm7sTay54NWeN1c7+CleUwXfFFAWMZ8HlRVXmGN+omazDt/DkaG
mzogcTeYH+Njy6qWMtc4mtIkniAaqj/LGyNQEJlfaDn0ykcQ5+aOEtkyIzL5h+AuXVx+QlF9PxTZ
EGdhfV4fL3XDsv6vFllq0H3c7i4oVHJFA5NtE6ke9Yev+vBk9FqzcbHkeBp1FlFD8PvFRLaGAoXL
uCkoNWoRXcRQZP/M7vYZtWCHkOaPxiuv4MhJV+uhPHCOkJhpgNl16G9y1y7NowaHLG+QDN7UWW87
L/iESd3rS8DhrLM4KwHRGDlxSBsF/+bTjFalhdbZ7LyxDXjTvfhpclJUPf2zxSBcu4xO1O/NhmJu
eMIQU3YA63jp/hoiZK6W0tPT+iSqgLbURqiKT4y9z4i6zdyfUHkJyCzVYDrFD0nvLpZSGDMCAfhH
x+WJBEmHFEXUE3F36/xTo/KDVcAklww7KHL9SGJyD5WQX6Wgsody95JSledl7juWaV9eAkN1uXE6
XUk2ZeHwuuKLaHP1YRvDNO4WSkxE82barkNksLeD1lvIsJ1HLs7wGDDDp/1/B8gGhAnJOZkyEB1K
pa60hqcg9M/oQKf+xKVOB0/RqhgQT6yy02ukwALKjU69wIeguDwlqVD5JvCbVBstKpqCCYpKipe4
dUu8KBDre8UXEYL/ZLKmT8najYQB75NiNDurEUFBDvzZmvVkssYYdav9PWCwk6DBOz6UR4Mnt86a
iEzflqd3ezsEuP0I6gM/Tu7nIzk5Ih/LEXkHxyvKqi4zrTD9ygvX50ZDy8uzTslvkNUGPY8tpBtz
hii+cXTvCP0Tuc5M13SHrugz7efC0KeGIXf1WO9l+qh7Z3GYW0tdDD5TxgyjzEWSXMCDuF9ReCAf
Uam/157HfZySYRJf0eabadblOJhZhDkTXDFfsiTDIjJUh3gvcqbuP+o1/YFq3pa3pBeYhfmmpUWh
lkWwLN/j74ot8R/SLJijK7VaFeSvinZqdPITYX/+DXRX4ZtW64YUDq9u8h5PznsWlqkx7krme4LS
Cvi1ZI53k90FOu32iweBqFrG/IKaj+xbKFHke0s618kG388fwZt1VL3f6I7/Gk/mYOUeQQCZBXae
cLQ4/1IWRd/KUxhJu2L9IZBWgSI2SE9WGTrJYqCBta4c8Q7k6ogYYvofENHacg9BtwIvzQGlno7/
LJ0gEBY1E6UyUUwB76s+F5P006FxBFhJIoK1FwOWVKsUu0XTQ3dKO46x7XP6lZgzGZkwz/8TOPWO
dIDLXdMeX2xgKi7vBic/4k5YYWrA+pt5ktuLWI8KwEU5GEIc2vduDYBDxuF9yp4WXOKEED1Dzu0J
tw7rtNaVBxbHWaoIFtFHNjSj7u0+3eAe09YgqEYJWd3avVz1PzQfzOUBNVIOhGBLLeLFexmuDYwI
do/bzEaP3IZJsl+4tf+vWvYwLMRO+YcvYe1+EvtcCPdS2pJofPvnaNBxCEAYpLPkOIwYryYke5MX
29LSB9bM5+eVACTuaQcAevc/JBHFkKGJxtnJ9TsMNtMKyIjHx7WSuXsNqSoKAIVEWrOhGuNp9EYM
pAZEKmpcp6SfP7B1k46HQgbwSHXOGq5DQbyLhOTrlNNG8pIzAOzrcPhBXuKcM10QHAF+JfBboeMw
+S5Ao7EC3NVLQpjC5HoGBkdtaxtDuDStUTGnbklBLv7vWL4HGtQHydhS8GfXZpLltyp75bRDlUrE
ydlJ5zCtFwtAu8FECkAWfoUD/qaG8q/uM/Y6ky052aOI1d4MdZpHi0tDU2Or6GcFJXMiuE8GxRxl
EeyLNStxakr5eLDoAdYCalGve3O4//nn2NBaslL7+uUkR3gmVeQ1CLNMI7FYSbbBnVe66WH8a8ic
XagiqEwFq2DTDVUkivBxAwV7y5wd6z2b1VQxJRTrGoHJHJZDpRflyQiGZxhEIR4sWQiDsH4cfAK1
pJoMRWdm55EHm9PWRhDSBruJYtcjSfMiJ5AVCMXNnXh3h9CF4RSz3P9SHb1JGspOcgXENf7kyjsW
nDhOsQ0k9IUCiyV2jEVDL2cdOeNRWrc13dysevUrUuDdZWJL0KR7b4q1k6lE3/W+z4jl9pc9Y4lc
NP5u2gsBLpQOob/rNsBeP4t74nPwBCwctxkiyPx9ZXAjVXFrdB/s26YUXxmcCPN2mQMLAlxGaQdW
rU5ZBQ/HjCC8vv8X8YEE22eZmWNHukypX5h3whZrR2eY68GuYvE47ryD2sozWi1I7a+UGr2i/zYW
KWaChIg4otpWWCBhVQLNWXbsIBhf2fcgVw4Mh52MyqjXvWEC0/Qn978fpneRJRC3LXnYKzs1ZogM
LbmKSiyiUqLAlKrePrK8fjRvw9ZlLrpDbcCuBI4nChvSE/b8g5PCWjjZOrGI6fhTx1AssAWihy6L
rUm1izDNGCwsRwcERiATsrradojIw5owMYCCZZnbMeL1WUyh8mGwqkmoaLbnH2tgjUxy9T8VmHCm
KPKNdHCDUT9I1ipyKn9c0CXlJDgknM7jADpn6hqz3hKqTmPf7BUXOE6YgT3T3F4vEF7bx4T3JG9n
Lsz47uo03HR8Hz9MUQWQ0eZKoW/3DM5EIAUB8UUxjDHDFvcQe8ZyDVhQOqQCLbKL70tMZo5fTI8S
fqHpqIX32gikS9PayCqTszLIBBw4X7ewLwaKIrBPhfR8VU4DZGUHQunq3fis+4WEWPRf/m9iNOEs
ijXllWI52L0uvhksNZeEV2cFqjYqW+uRuioEJA/dquH/T80xGenQJQVxlVHVj4OIosbSsQ2URFXK
PNKIVswsmfyU01MlKwwo7wSl3bjZksGLp5TdrmP8MTb+qa0mi42oCoS1xEgawgnOq/gQTC+m5X+t
heeVhx7O+Ur1FvnWPJxV77WvH9essu4NC2YngbiTIOBvNywXTlLCdygAeqYygATBSGoaGdNC7JH7
L5K5sPLcc114J9jLqH8/FBtVZCvmY0AfPJgmkLoUJ04DFCEqK7mQQa88UVDF/jiOvdFTbXRapTMx
BxOnXOqcuLCypsG3BzT/BD9eFCGENKFCpAnmwG2y8Tgu7b9Al/40zfwdHrSQUIvMS6u1LOy88n0w
NOUSalW3hr5CM/JBXET7vqFzOJBG450ZFE8MMOHdAxllTjrGs0hwZ2Hk5fgH9e65uzkufogfclhs
Lm6eL8Ne6bJ6QuSGKGBKPWAlvCH6UMtCPryUQflfm6cuPyGR/qoZn8eVEUYqyA3B4egTLOgCgB13
+5eMBAhJpBUZnUhKpyraXq6yQawka+cW4NxKpVRS189gBJM7LH+FTiwrZjnrFrxuWmd3WghjG4Pi
0vi2c6dUFzeSnkuUEwNdv+kTL+t/4HrlwYH7qxWuPXN8zPv6PvkVC9byYo5XGfXjnpJFrAmiKDoA
YnEyodidVaBDqRp7N8BGlfq6HdzHOIJRvGSgQZwP7ZwlSNasVZz2CQy7nbfzGEGCbTBexblGFv6d
fC8/+qZbdoaBWqZwND2uQTDfduYrLtlo1vXV2QBI9MYST0ANxEa0DM3o4he0P0+IbXhzSu7h6O8r
TOBHawxUUEakU5B1ikOtV7UIpCDIHmKc02niJXbVg78muIS43uRNDsSHf0Z6xC4SzYy+4J2eFOEa
xgJ2tzTexyzDtxtYgTYydfQj8hQ4qYSlCtj/FB9GmEKlKt3hyW3Gj4+rzOqsEL5eLo20pnrgCg7q
yVeBxhRt6CqgEDqj0PuufHlnAz7QA0+8IsBQl4Y54aUt60fCMse803mCQ6mnQUzshRUfwGDoAZ7f
zYSMmDzmIvu7ncb/5Uy/3Apw4KpHCYwlEysa7jozpALi5MYOhTMEmygPEuIbEOTwMZnBSxOmll6o
vkbPNc/u5qn7x+UMoG0mMqVxn2XvUXVxyAsVRWcgAZdkN7TGi4FnqIQWiUPpm+8ll/bvmGB9ilUl
84wyRVFMFEokFvVRbb6Q9WmGj4UTq/MDouI3ny9ljpxYWQyjvFkQcOI3Iy/qiLyKuBSEqOvsht3P
+0PJAd8pHVLZ3pQdPqAFHU83dPmBEolS3oVPG9yvB/jJ9O6NPPjdwXqKvTpOdAurAEoIlZIrV/nr
tUGtz0sfWDD+rfLmoQhq20VzNhWKVxuqsRuis8sIIWx8Qf81zZEl8USlW85SrQR4YjNW3j4lshpS
CbdZoMPwKt8DyVBdSobe7C09FWEi/ReUGlW491SVTS+zJfMKwDvWB8Ow8L3FIeMfRoqbFpqGEuob
FjtkmhuPiAcS6/SeVU4bVcuu+AXTRzvPrtT6WCtc8B4RKDS2y2XwMjaHSawiKB4kNLKknDQ9HwfT
D5Vma/2aAzvHFUoJLufnlEyeiCJ2NfvIFiYH9MjPMM9ShY5vN4AlYQNW8pSTx7PYu1qp//DzjvCp
ozYJJFbHPOKRBKrBa3Vurye4WYpenk8XhdHdVUxZSOqdQgXe38I9Ns9RgbokOssXrTUS5znIogVy
hDoGc04nmeUiP2Hd7/t1DXXfSnXPtcrJR/g3aeOC9CKJh9Y10LI1fMqnLC02Gbc+ljoTbAthnjEH
96nX0okoo2WPURUDNASRVS/RL8AMmVmlIBW0mUOKxKmNRJ5UK9Us8cMN6WrLBeEKyDO3WJvP3pXM
aA8pbYNIBMCXm6ILQn7ONwTxDkhuToG9+aowXlMBzakF7WXWIPCxw6IGtF84urlZyeavPqmdtkIq
XRf7lvZT5WJYh2D/rCZ3pmJDI4vAnWDgy8Wr7VsbdNk16aCPsQj8g57XK3MdtQ+o+dIz1e09kklD
TI3lAt0CfQmgYb8iz9ES+RwQIFfm0ZLA7H/oZ3+nAy9Uu36PiJeKD/SUmMPilcmbrsbKeHy3H4My
E/hF24cH1JXTycR+fTCk7qr0p5IhmhCVIyJgj2gAPjnLyLPaU6G3oDchL+aBgp/+1f7Jjocd8nCY
tJ4e+Pyu5Ahu6ZhThvqvE6Mt+kAM/JeGnDWuFez5kQbCjaI0rkgGObOqz0w1w2ba47krbtMN4dd5
avOE7Q4YCH95HSVBz9umb6zILePI8M1kPDGbTgMOK83Jd2rpgYYrRG45VItxXxznsOQkfUu0dOtO
w2+UvElmo0dNPKJ2asO80JBQpbHjwaOkyWhsTpdUfoakT/PNTuUGuUw26f4L1fkFXkKI1O9ZwrbH
0BE9wxmRk/h5SHjmjTxqBcp8BwXzppbEC9NIREFQp/OcmQ0BO46RwRdYTmU2Rp2+uFigG5uDSRbz
Hcig2qQ4SGETkp9CCBNEG/bATZp3GckLPuwRqyWYqlyWrU/pfGDgWddqbJ0jJTmxfByveQiUHvv5
KPLUUXH1IdFD7J/7Kwsw2ECTwbMQ1xnnIb8jcaRcQ2s3AN3qjvaU73mIxcUInMqHANMrPb4pPnaj
eykPqNFkj9JR0YYBebZOwRuf7hI+aXnhj/3IQz7jc4TjV6Eg8I98RH8MSzh0WJ5ubLVqB6916de0
mjMEkNeJVfo8tjZ4dRiI9ASpj7WAFFoP388iLZzrz0myhgt9vn6KCVSw0bvBFARC6uyv/pg3A82J
lV3q8ODT78FqMqmUhE5s4J3//nCKZAIl/yMW7UpJFrXp9OI2phpMJ1KrFG6gHOSJlmNPOhErVTFV
ix7aK2L5VaGUojKp52Eah3ziyX/GXQSsXgzmFkizGoP7SMYeFRNDYhceFnvoZVLY5IWe3fCX4Hak
LVmg1bQ32nx+7Nw5eT/3qWJk+YOatzjTKXKAAWI6m4ZaNfixRPTHZ96ubjfnq23c3TBsQ8yqXSQ6
qEcSgdKtDtLoV6hE5VyBmDJxIUFiwyJn/XWDoQ7vSk/gGi9SiyvTVMG0PJHmrp8cNjZERIgLjSVZ
QNC4hoPToXt97bP3SJ3pJgqrWZOuOPC9yk2MNhEJClNK7cSqz4P3Vuq+XmMsWIgmgDyRX46K3Pgd
08/SvobfqeUNViaocPs5GdWmBThYPYs0i/EKlGX18g40JqJmoSWfII+tf810Qz62RrMTTHH0kZ6e
+RpV2wd9/wYYPuJqrLq7rReiUJTy62LjU1Z+GO/Ymn/6zkpoAXETcJa2jWgmBsED/PAjCiTY1zIZ
MEL51yaGjx8YDIAgjg+jcblN1k+Zj8dySmYK64vAUnwJUFUqSBL6YwPUuj4L3ReFJO9jdUynbVCM
wh/ygBTLi5ktgtuJtSxVuY1ArWpW+qdnccxjz06cVz+7w3GemtI9QZ7NW7eDZu2DIFIVse6mZ8Un
gMm7EMk7RHqHTQj6ypqHa0KMvbb5U1LCVkEJcEO2fWyYW00IY1tdG1FA9u/wCEJh+AaygoMwzdBe
/m2GhJ+kFqkNEcMO37JKdkvXnVPOIUqX6HQUswbNzFY9M9wLPrlFBRocldDKXpLb5anE17crbJ1O
kDAAOaO/CRAYdDX5kaB4BY74NbHQaxdMXLadr/ULUMPwWrRxkDlDqlTkJus3OFvX6TkOItjQpBFI
MvRPKDpM+EAy8UuYgWs/4ddDQlxp3YlFqmxqFBKWYgvv54HquIUYdzVlr9/QjU/lla9iqUkwJT9+
n5eY4zZ6iJWPBzQ6XO7pj0q7u9ow73zax5BNcrDJ7FRyN8YBrTQnQzPg1+nvho5AqHYNA2twQFTe
Hi8ucOn1HU3mSXn60HN+WIR7/sh0sYJr2hq/N0+2Q9V1eijRlmEfzgMlerNqSSfOmZZ+MODRNyaG
2x7zSSqSF5+PFyvtYkdMBZsNcnyrERkpiOeRH5PsicJ40sAQYv4mjYXwT/7sz+jEJ7fOca9kx52f
1cXwxB2hMK0PO33tuHFec7+AxBYAO8Gd7g8VKIeqCOgA9o8pn2WVE9Kiz3bdjjaythy66Cu/GgYQ
49CW4NBG8upVLm4f9st6VUJmcyB4arZApszdoyhk6aQ/z4FC3I33/K4vHzdWx07eQ13+WROnP4XL
lCUOevciF0xP+j2WB5LM+xF9I9UHifNwytdQ6zZsi1FmQTb+h58+oaJDJmXjQjglQhIIRp3r7QT4
NYs1oBspfCZi1nCfaSQJ8/lUNy8RUhXcTFJpWWRkn9fwECHZrdrDxw+ilXqGoSb0cYRCL1C8YFSe
TOJZLw0wPfoKJusHahaZThEcvQrFCJUFw+C2bokAS91V4JaUjWACMs83On1BnZJgFiACMq/Ab1C4
Cbsglh004qeCqYzSxfyDD0EPCpsTertUTUGAzx5kyyq96z94NZhH7Wbw+vzImqplGtaZWWZD5bNK
u/AJ9xviY9yNdeX+iLrOPW/an5hBNfBXEiXAn7Er59Ytw9Laf+StlyeqekKUnbe65gnbT4xgfv9s
yoiqSEcmYVQuQcDzTOLISuT/GapjLfCCJ87Vi9XUuQiF6k8HpZQuwZ0o3YcYTQHjm8juD9DcQ1ay
lTxMiJElF+EWLb+97fC0LY+mUbahIxtN9x8w8DLpjzZX5AJMCHRB5wEyp9knSuYXM4D0tnfPlBc2
YFhnceO+ypp+Yql6OOgO+HissPymA3z39H7g2ZSez3rtla6A60oS3BQMoEBFhWrw9zAyyoDt/Cjt
gsOXHzzMTMnkdIVGcHl4QNP8zCxbTZelBREORF2GrtC1PY9j6sSJw6Dbu2YjmS36vFvdmB/22IUp
cs87wI79LGvQAIqxWevcyNB5aPXcB6aTTZxy+/5Z8tXDYz/S7sAEF1WeF/4oTVsvNsbfqZXQdP02
sYxJDimCe5gzxQQQED273r8aET2FTCkqn2E75Kqx4sX3RaxhAExw+0HwNeDUf7h9+6sxZB/PeWSr
1AaVUXWc4eVQwfYMP0ebLfgCaXGo0pnZ09UACeYVVo0jA/k0eBiv5rDDX+1Ep3s3BE0MhpzEQjTF
ycJZGnaJxA9FrZ1zStwYElC4xTfLfekj6veUQThnd4zdmXfBH29O1BMoKWIvZ/9ovu4AoAYxbHZc
Q6FvIGxcihhS//biWM5TcJyX2lQoDCLmG7quytFXMphAJ1gonc8uh1SLvzPvLuClzIhxjFoNpK6C
/zRfzgaQRdonpXkp+zL/vl/P9PDDdLkH9v1WfODUHty7prk93VIL+Ntd8prZOcl9C25VQkFkzsZI
Jphgk7rrsSzYVPaDWTNQYaNB3mPcDQJ+Go0iRVJK5gzKtmPD7nQCSBJnxdzZ54jJ6jS+8P0W8+N8
/MzGZdipkc1RY5uhtdubTmrZG6PGposxzsvZYtzWSAh9Paok5MY+1u2n/ulwBt6vk9lvdX/SykLK
Kc3NbA7OEwVQI87HGwrbdocTweBRWCa0PRkqgtSuO6pDh5KlF6UpC4dWw4h2cVXm0buKr8zg7NdO
32qCfaP71LqIbzJCePs7gS6paIjlsmKOrxlNA+6cgp9DPL0MgPDbOy2Uyow+KSa43oOU1PZZrRPl
AK5M0I9jnCWh+T9Ehwbh8o231T3ZlN1w5xdTO0Vd6N/1afjWsoELpP8FgbwSojOl8FdZFAo5yWA6
vJIou+JVJjGmIHm+rVym7W1ZgVOsCISyQejyawhykddNGIuAzxIyR/qVCJboNGcJP0izLlKzumxf
W3Zd7B55yt7q+olYC+SsqP8bP/O+cpzjrqD2TqUmZWLhoOTe1G+rEVutCHVlHavTZ8k4LBsqIJEF
p1EkqnH5JEBn5Z0Lo/BcH9ji22JdY2tvkkKVmNgVoDKPpXBxsu79iDa/h8vC7KbzfvkVcMDLC1RS
ejaKVlYRuSQX/mS82zRnyXLNeeoJgSyLrgaYRCzw9bide+GBZbxwQO4UD7KO86Mz+cvsaP4Fw0tm
1tWKBXRHyuenmc2dsi/Y+axcLE21Ps5gKnqSxPDTrcHXyUkHjmmJ+PdmgTXTItjyHoeUCJwUegte
RoHR433xEox0JYxwMoVZR2fw2cP+ndEInnemhPlkkUu+iVTAGdSKhnPZhl+yr25heq0u1iaXBA+6
eqOJw0iKLXKsUTY6xx8Rz37UJ8mMP1QMPJDp7IFbxCZ663q8/1OH+WOL5gwNBqXbIQu1gkqoB75W
tlZaVHUWSk/yoDPrjlWsYrS9Ke44QiZRrf1oiOhrDPy0+CMAEoHsz4XsNVQroQfuTj+pSKjplrtJ
wrsP8pJXGgd9mf21gVeUC6o1U5ZbNsAjxCql9HtRPYiy8KY1Z2LS8Cf2gcX9pQn/S81KPMJWfnBW
ZkT3twZCSNuly7KYv4MwO2DykP7hbfkcw4V7Dm47cysinsUqgjfFDuZV3LBuidYhkmifWZ0syDsf
9OOaVUkvz4CtmodUWWnRpEZTcU42exbWcmpSFUk9gAcgcMgaXAxYvq9hj2ZqxJUsYRxrDY1lyjHA
X8H4y6Srox5XS6d1BF7kOlHhlwTgY82XzPS6KPSckQHxqzi2iZSRxoH5wqiryxdLq/egeYSlXOsA
XokN8sXUWkrFe5yNFE5IDGQTRzLAQcF/gcWLMCfH5IWRWdnAJsu51DV408btNpBmbznSJO4w4FIM
+iQFiD7wZBfcMtmOL7/er3OEDjCousVJFK1CRp+Srg2e8h2hJIFriMC0OYhPqBrGqlAhtt4J+zoL
XNXFwgq9sHksXWgZekt1cCqrlB5jAmUr6CuTu5+7KkNjEaLxp9FViNUWbxvCMnd4V0ZnNmyet+Cl
Tr1KX/niwjN/bmjUkbgcsLBGyQlHLSY54cJtlFwYlYXEuHKpVUQIOpQJ8vd8T2PeclXOfuk3CVam
uN47NQc0tO0xALlTtlBbjVxmnsZvFbMCqGXU26rpA7Dc5HYy2RgF439suFtw5DLgtKnya89F7aDM
D3QAwmNN/36ZV5Vvy3bVV5filpiv8LfXgMgMmjLcXxS2jNezBlNLsF4W4yXdxHbwTor9peylupeB
YUK6r3B2wYYaJkDMupMYOtHz6/tEszn/tNz87EqfoD6lZw/0nU3ohfaAk5CwzDBpG4inmfwIj8pR
wusv3oOLz0ewVkHNhWiGwO8z8eQOgV1sXzVuaCNtFgTHjXBxej4tJb4JqJHoFxbyTis70Avgw4h+
XZRbIuCu8leFtuEozkWs1ilbxT8Bcpl8c3XpUQf9ByiyneKH6yGCrhG6YsdGozmyx3blEM2eeHRN
tvrulDNx5Iu5mfX6nQmM9Zywvogo3bvT1EVXyxtDB1E7kj4XloZI9gHdc24SqDfhTlMNacg5EjXa
32NmawYfgR1a22a0aAvLXdwzCoiby75RUAnCrVtE9/eqd5MoPacnWITh+qxtgCtbJrnamiktDlHq
x0+lRbukaddayow05YSM7Hdca4lAtEyr5Z/+f9fz5AGQMxxYrs/dBrMet1nIc/I8+jUm9j2IovdC
6gLO6BK/xj48NoRCeljXCtVed0ns/5BlUPF8H7OQKTkifv2/9mIutPfdmgwWJcAcqL9yrAlSpKpu
il5mdfKoPxG1+zfDQVOeLOId+4W4Z6yF/OAqZ64T/Ss4cTDd07l9pqn14/5ci994tNIsdOQ428Tf
D/2O5xUMgB33my/jwVH4K4yAqLdrZbdRyUPYQkkmScYn+y1D4DbBEKav3LM/0c3PKjACnypv/+va
avaCGcYrP5kyQgwUew21OqG8OzSFxvESu8R076vR9elkTllFAxfA3u/q12lGInUn5B08qafLK3bw
ucr1ljX7ronBY+FZSDWw0qlPRrtyyPhml8WxBrh0RpH9GPTo8ZMrrGbzxSXHHTeiJBCr2AXp2lrm
FB978qkMTeQM4wx/eHz4OSz6ppdQo1PYTJjaSl0w0KSuTSpMakg7JIhvPPANuDNQeBjAajrE8m/v
4SLehulJW5EGrRFR9KMOP577p3nos62Ls0HorxYFy9okNjuWYf37573UDICkjJMf+jzzsAKC51zC
fkMpDoTZVTJRAcJ3q4GIMHiTDIji5B5bfL7gKOSPXNEV9NC0OxPtwaQh3RBssZIvTmaRQyv2X7/v
QWh/QagrOzkhs3XjX10to4cUg2orTRqVrx/uHii5vxmC1Ld9tgder3lO2H2Jx1e0dMg7DUtOAGh4
ScdNiceZkhth4qxXLc2vyiHfvregjAtldMJ7/OyuoMzH7NoUUC9QEKPXwGtDBkHTG1fglpLKtpAK
SD5BpW66eIbzePCyVtQAOt8bPoDDkDqe6ie6v7ZVj4O0nbooZeF6Uk+NQAGeJ9oPgaKjVDGaLwYm
7hZKqZ8y1ElyTnMFtH5+nIPfvaodghMH3ykHg000tissUrf+2ftyrm0nqSA4xi9Q5YAmheH+tFFH
X18fAsbn9jJpuay6kcxv2z1K8iiA7zGfZEyyzQC0I7Ceiec1HEfB7LkCbt5wYjm6Pyocp/8rHw8s
qSqGtwaETexNoGc5ko81sqdrXV2zH4e9d2FduCDL/K61YRD1GF4vU6CKhzrprd4Tvt9NhkzWcRQM
muxyPOojw9SdvVGW8E6BCSv8XU6B1Y+Pe38yaAswediWKkLxBNkHRq3VmZSLbLZvTt4/1dMnLpeA
rm137thF3gnXCce474bBix+2sBy3ybM1PL73ND8iUcrZciF2bEDBg9GwIp7NoExGSgpEppebtYJ0
u5917RQaXTsTtY1ilpoOO3haLpbSrgehdOECScwi7VA+aaSsrI0NwKbz1EVEvUr8DyfWbiYsx2bt
+hQMjUxKltwtHJg0C9QbokaZRWQ/EjBqmJXcaMOlppVJVycmz9sYUXriuKblGxQ4+PbqrVF5TkIk
lhCweleP7v7Ta1U79A1e0ACbh43c/uO53+PEWmFGwn9GONn3bsdsIZeoTyU7Z9+eZPOznPzbYb4f
Ak+hv9NCDDlJTI/A+V61bv/nK4bX8Gqcv00VHbqMn6sOMUAVW+a9GBhlCmvgnFb8EyLa0mhi8uzS
1np0JbFSWmCYIRVGynJauyCz5rH9OIikGsvXeMQb0pf/8GegmvSvrxcBX++s2QZu6E2j006JV0u+
Kp+fip+UlsHGv6p8F0Gd3Jnctf6E9dyzRfXx+zpK/23v3zm7AikrG3IALr5czo53YAkjWUSSO+UV
poTHyy/uv4KXPhLPetvoVnBRC41XcRuBjX1iz4YibyS2O7ulhX5lKLHIubyzjboglV2sVSK8lykm
pGmDasAUeQaJ4UvbdD6jj4dB64/4hzQ022Okz+ijeRy0crR5u9z13pSsDjZwpkozcQ8aOcRZP78D
u3AwDq8/AtnWOR5bLo33aURHnvAhliAb00rzOQ+MJCrfW8Dt2C49vPTO87uEYWGL4Tkaf5qv397N
C8NSJwQcfTWAXJ+74GN1kWGWbPdEFnGVQKfx+npk0gTVoXUt5TP2zkp8mue8otTi4n63TQ6iq5Yn
1o+xJ5iKGcE9TngvWF90YZyA+J75HF7zwXs4vTKhhqZHrvpOCoMwybYhf6v876l75kpkkAgCs9f9
H5DmxEye3gV10dLhlEPJure2iImmVdPvCjsWrlybMDi3g5vwgkRt992sW1jiInqVow8Hd0vJX6Nr
G1mXtcqHjHjdVdLA3MZDmfUkZUVVjAXFFGL6iVa8bXRPIf+AlcWx2iqHVeBkauDvgNUnQREujuxP
50vAGlMqk0IHouVztmUKrQ7yR97iN5O5N8gFneG9WKDOgzUdwOspuI9VrqgjHAbgDztCY6nPq5vQ
nI6kCBpTdmCVdrOWpe6++6o1JJXTR94BNlre65iRctfEvqqrDavP+Kchm0yjYWQJ2GE3lowKQoy8
jaenr3pY9V5ZCFjf4vSyfyTFZm7WYc5TPRnQugjgbvzAoEuoPKtXJRpIWXvI/PJkl3AKKsyi/Tgu
a24Er3E7bR7mCxaf96dz7Cdp5NCA/Kh6/9Um3FOrSghD5hNs+o2Dpj0aJqwYKHTgU6azdlioPxwP
9EGnY+D0Vr/5+Gw4wWZxMgxG6Q2qaSIm76BHaGR/NpSzsPBYtFMy1zcEfm1QVdLWD1Y//ezJTHv6
28FyiKYVSYVbetEHzOtzAWtx2wy+74NTrwm3PLYEtrdveiRoGb7X1bbey6PWW+xkJbQVeFNxS6s8
uiwr4YGjiK0QuDYpkq5aisvI9574LxaddCE8kqndnSsrkXwkuwx6RRFAACWeDza0aeByTPvylUS0
mUovPaYVnyuTHbNz+jkQNmKloFOguGOy64gANI7KccroU7SG4twvP+Yb1q8iVFFZiE9nPTlHu5F+
9jrfdte525OAOYmXWAEk1vvehcTdBP/cfWS950V0ki5rmvoy/d3MTdCwqWytVHh8cNIylHaPPeAm
iyGpXdc10OL1ElOmF7X1dArko5NvYG+UdGGfk1jfC6DVB4ImDaEXasZ8YcOW+u6vrKsCAS0ruKOt
qjZDtm0JyJlsPG79YWG7T4uBoa9q/BmcZuKTLVB15LJL+H8oxlKZFc1ll7pLP8nYdXKYVfWbu7ee
RHdzqx+i19eA1sC/pWU8eiw6VwEQ2gRebtl8JG8bNvqC58SXQy4XxLFmyjsA2PHmb23Ok2DHo2vR
yn16CUKeLw9GusMk9gvuZsDwx9v00+oHj5z2jBZEfC88URTfKiDwRo0mA1RrXCS4S98k/18SInTV
0mgLz0JVXLxlMhMVHFtDVPVDTtaVNo8XXvpdnJl/ncH5TvTMQFaXgRSaKvyB2qezgTzVpZ9GYXpY
37A5EydxCNIaf1Kj/cbFSVeiC8DJer4D+NM/I9kRCvuw2NQCSH76lWNkZGluBulbSKoj8ANq/Rsk
dBbkvPLMsVAFCjfuqxxX9dXdc4/LdnDFijJsDFU7MxLXnG8qBz5iqaQ6pXOMzI+XKVnDFbhW/Ncg
+IrM/QrM4JBTvByFJWx1mqMt0h8lx/JuksL7YRKVt31XwDL9UODkrrDI8RFa7IsEuDmrsXAEvu1B
p9mqVezJRgFoJPrge96cmVwFpDnGBXAw5l6xswPEI3VAOy9X2YiOxkHSxXS3Dpx/iO0qr5/WEROA
HkU/5uNtwyRLAdLYedXOpuqXDbB4yBLX1/UXLYmQqgoUkFXEiCH7FDQ2/xeSakW3hh6wKL+KcrLu
vmzCnyDOXyzxa0YgRUPQEx0aPZtbbbE0yBFLr41wmVaeHq0VPaJwfQuMphO6/uQu0ifqXQjkV4XV
GslZunYqxWEcVdYBiguaFZ/btEpAOXwvEUCo9irjKgB5FiYa1kBWlhi7QW/G0CoJYyROGAQNG8i+
tBiBcZoY/D3LQ9NwhF76I8fwYYUQOmFjA5zKahOwdcjFXLVagX4ll+uh5cgQcnNm3yIL2hFhKoN0
yQ1bdYtZgeN4IkuaNGcXuqxgKuMTdyTeiMJ0Cs8mNM0b90j9w+bBSvbVkq8Lr4ROO2IlnuxW98fE
q2nvYEIEAgMMn1QhTcysZmAlPkG+SDaB/KEi1dhGXQfOFAsSK6gNeWRMvPTn9DcQfKjKmpLMY0tC
dPGeyUE+9D5OyhxKgYVGGrZ6HUCy4LAFajblB+1bmU9+JCzZnK0NmR6YCdCxiWCvqTFJ6vnC/nW7
GGi4PdV7bqk4kfq5ChJVk8q6LoKkGEZPI1wYDi/ikJ9b7QZ24XnKebqOAmrjHh+bBK4IE5Fmh2ss
Aw6DHOmeGmqrpphyqTgw8I/pnS+sQq1YhGTC26qIuKbcl2RaGZv7NzWaMcsxp9ebA77AUTuZe2v0
wl5ECWw7B49CXe+Z9iK863IjQsKoR9GID+yYHALyLyb41oM5beFNVs2TiyncB6ynd9bsm3TLSZBA
AbSOqWXNM/yM88HsRvyxuGkfqdPWOv6iiLAHGZ68SI/JOJHA0z9pqSpBXmSFSPZuc+tvJ5FRq9J4
gKrktRlIi44wnSJyWbpmcJWHj6Rbh65HXJRwlaR9czhvlpQSwnw+Cmear6XbSg12cTGmX4kS+g0T
rrpO71Qc0EnWzMbT0MTxwSFwpFgGykQrMOTNcopTWxVl0/Dgh0ng6/dunxkU5/bcKvF+UR3i/iV8
cYvK9JsPQ+By0ROk654kNHrXbQI5uVtnmQ6dh1E9Dl+laxB3YLN4IfcqchRids3xc3OQ4gNJfb/k
A/7uGUxrr+SWqss6RlOhAEb0GuzK/9xqEkBoeOxm7GcTo5kMss+DW2kmiDgQx2TamclFZATvjW/q
UunruhZ1jTphL67Eb3EwEU1bGdQ84BfuY0EhKk/GskNEn8Onr7XWUomk6qT+X2K0ApfbR6QfRf90
rHckvppz5FvkRKEHlZ5pFD6+KRJDLQK0iZPr8Q2NebJ2IpwyjvdJsKfBRyNzIrjibRvjzZNgTFIg
qVL8MeRVaBSQnCqprRGQAf/j9Ln/BTQUYTp8z3zi1dDn0ClhL2n6ABpYrSFbe06aOJeVNPDyEMWj
AGCuZfNGoPjwHwNYJdKspeUHFpCCli2+u9XmVFttslrzQRs/vuXXCvtz9WD8KWPIbpipzl/vTJ/j
ZvFPUlcbUoJSupsJe8yG3SkrVznl0tk8boPHhd7lUdaz8JCOjZ6NwF8QIKUNW6cTsf1vSLNE5ug5
HxVG30owDmkQEjBfzdsEStpKixtbUA/aT3BK1eHR2v44tNcw9YAQYJs2Fne9Bqu7k1k+1ZaZa8by
80HzGOKpnQt6iBJwzWuxOqCpLUoTvy85KiWmRC/RCJfeItQae7cxa7aHaUBApnykht7bO4Ux0RNw
45yHLV0MqqMvFUPDbDsDZCSXQtUBa0fATQIKQa+oStqiBgMeJrbguFxu+1uRHNgXn6vPXduhLOWh
iU5ia3EP9S3D1FQbxC2CkP7Y2PUP59zGIELLptNBZF1iYroWLp254MtEqVskFyxSkQQHP1PVQ6w1
5bCL+H/9rLp31Gs04fwP5BjFnOYj5aGQwoKnjQjrVNAqWF7PRHmcUm8oWlBxy84WojZFtxxlU2MY
zbTtSn/YBd1FMHYuNSy4OYYn9SPlHvtrPRuUdE8uja2XiXpfKor5ZOV3x6AkzzJKR/tX1VlbB/q0
1FSmTmu1f7UFpubDNFDX4SFmnBow4ThLnkPM2xsj5KGBZw8UhUAcdo0rviuf08SUQoCIqU/1WPBf
RL/ucPO+F2yaC8Pq9LdnIF+76GXa5+EZ75jSJlBQxUYstKyepXqxZBerpOIUFCakFNFLfYHZs7kf
FE4FdZ2GzZQz3Qc7VDZWPKi93LNOgMclIT7Lf+XFtUxCL9weIDbWwVZxx4oaOsfZZUCfeATz787V
oHjFmLPCGvUuObKCbXvvscYFEDz9r/1SyT4Rxs3e2pXt2PR4N+S/OKyA4VQ6I1JoeOq4NUcQlhi5
I1wFcxjULbTZYcBis3qAzvAoHrDbOabQkHvMSWWCu3NuIyS957fKuqb5cP5lUAD+25lWWkp19bje
5x3SrCQuSfChk6BZhOmc3BZ+Mjntv2GyytpeaL8OBdNcrIr27MKfCJWmMuJteatmVGXkZRbNm7az
qNeMEowprPT3sGnluiqzbxxdEXRWqZ8wZnHo7Q1mv/xZERuQj/lNWVaCl17xlBOc1fHZl8JXruMV
6yZTm4TM/+CFA9lbWx2sIgAOFa6AVgO1Q594yPcOZAiVazCE1HVQePG2k6ZpEggv8UVH4ERg6uxs
a27PU61LFGygKUpmQbLyhz/+Y4nHA1agorLNSyPfP74Y8YCapHK4+2io7aTRKGc61zvRAwRlBAyu
S0YPmxtFhmxHnZOaWaLUf8diFFHBd410LlgFevQBG2ohn/DEwrTRAi53Z3IwqBk7VCbEMQEFAqSL
KYgRPNBLjnRwIovC+Msd+VCucbIw1muPhj6ShcMMeScMWPq3Sz7HbMnNdAJVYOIIlNdmJ5/srSoK
ePx5Z7lOMpSba+4QETcqpfRCgaFzJjVJmw56zXRqnDBCNtpqoC1h09VqOFDysmGhZXGZFHskvCLE
F3RxdnYahz0rlimjbCz8DqQPG3o/s0sXaVoa4gFH7+k3t3dEwKLuQgJiuIKTBRD9c8my76zAX2Lo
Pr2YuDwm5lnU8PN1IgHSUPXEqu0aBpqR44ZCheeirqcFtxhmcTEcRkAzkhv7qJIlhRmwetWAdU1O
P+Mkh7/JbnLVdXzhO/5DVG3daHLO+ZbkNjmtL2xfR3ARq1jdR9lkWoFSZaDcWjQhL0Use6r3B3Yp
aF5bCodLVbnkqk34JDYEWbpscm+pp6pQ7ow7JKdqKpyhfQrp0mr5atusVqf7896JlqL5c5OPZ8zf
wvzpzNdnR8sBIYMCl90pNGaSaAQKAiUr1RCGxdUfZnM0lYkoaddhuaqnJIUYdKzF2KuOHFQlVlc3
rpTVlv4rSFu5+ebzpZCLPqEc0z/J6OOTEnkIHYRX45mi8FHPf4sgDwgjJw93YRM93UwifKK9NDct
kMHMT1vsAqVxhN6dXoJwzDwbOsHFko16j0f+e0OkmRSmPyoSe/a3JH05Qz9tKtOWQPN9+Z4zaN+k
8BaOc78W5SOXmfCSPEk0HY2PRANpAj5xdZcgSbpwCaMMf+dobNeoavg/83T6ulxYmQbAYP5NseNp
LiVj6tDsX4K5OAUMtZUMmNSlPywzvnzrIBrA48VMVHTfWuk3Kt3gmJF7qtK4T3DJmoKUtz09SJiR
Uv7pM06EAXEZgSHEBfzwJ9yCyUAgKvkK9nVSVut/7f/cYixJayPe5fB99mm3DrUY4Cxy/bJ9F1n9
8TvX2HQMM+xTrgEYb3dTSLDH5OIjSRmI6JKQ5di5gUoJxMoI+EQwAvife0zA7SsaKNkgj1lzxMS4
THVsyufLai2mY0eafjyiS5qrknN2TxKSp5VLAQXgTGufNNE/9ANTnvDHSB1+P9/E1i8OAMK+d/uI
1sXiOsxctezO9DQwEReYNQ8LfkSkBAn2hRDoxGdtjkHxeJmMv5FDylmIeeUWHyr6T/u+YQcLoTse
bJq8w7DX7Gjslv4C4G/EE9eVSVgsLM6xkR6uWv5iL+6PCEPSRdBP1AHllXStc7Xtj9+uu7sVV+b7
xKrk3dedAhoCxEhUOAeb+usxpaxvoSuDVdcZlPpl96dXw3rePIaumbN6M2Btmu3BzTgyi4e8o7o4
bwgYWu2liUZlB3mGk95UnHGCYBn9TGO2JSqJxCVdQhkc2W3U1G3eVonwFQ0oZTLtFYoKjQMUGhHG
KnGNCWHRx3CuE6DaNJ4XdYBx6C5iq8+8m1LO8d0YOnY13i3YBNhO70nlvYsik6ioL6aYFVrv/a2U
d2/3uzOdrXRkWFXSOHv7o62b+RvBteAgTw1/c8PAwoRBTlmUM+eGII51qvD05MLt/LUOY2cU4E/w
DIV1Bmc1h/SxR4WpcGx0s+O9CLDDdZNDHv0gZXqlgZahgCVdWfVCW8JqqUNQA0EjcdcgPQAb68uc
pjulGB9hJianp2jEJT1PPoffWtQnKTarJ8P0budhVypVadzVmKPDxzc+w5x9/i4tT/RNPis9VvSH
qi4rp3ppbvrsTasvnjLjPzRwq+sIo7S63RgXSHu9goqSA3j0rdM9JbduDUUtgykafzPAFgoaGk2X
vYks3d4ggzk5KgFXQuBKXGGJAKWU+3MxPTyLB9TzW9orzRLnaUTzn2GhgugOs4b5AzJFQxu8qkku
Vpm/KrWPboJ4IxbD/E+2Q52DCkzMB6fLCgD78hA+hK/+cOvPdIf6w5HJd7WmANC2j6BVYns3Ng3w
FVYqruFN9vNOvCezBKXXoS3yD33zkKvzH+zooG8Jok9LMzZd6RixlQAkA0VPL5ZWvJe+1H/jyiUl
lkEGSD7llzt83gHHZLjmy+krscTK9Yd+zD7NYmf1djD72L9+Mbsr427IQnOAVbbDJC7FmUWawcJr
KxvEe9lnW2EFi0/FcKDYhiaNhLwtr2kEj2U8pLIJsBEp7aC+TLr9SOj2ylLRLXdtBXsMoiDtKRrs
8ZDkF4VXAs4eVnWhFCktmB3+a1gnU6CbmttEYIdUulTwUEe/x+3k4Mn1oAF00H7KwpzcGgetemsG
HN/3nPDiKOIUOS8TT1c2c6TdCrNyQ6cq+2cjr10ncuRvzqMXmAdunevmnkIlkqny523d05E7Xx2i
lF0RweBn5TF9rDa8Ld3nC/RsX9qOs5hlV1vI4XNF0pe6qfO5eapwHOsr7ooSaSlZt/8Hy93NSxX0
AoPS/b8UI4xrEN4Tdj7+XdPp8BA1SZr8ieC7zpHf124FV5lgd67NcB0HJ7H/Ur3sdpgV3vdb2l5N
CWesATqX6mOSx1cFncSNbxSUNzv7oNmZU4JFPiR/icUS2UUO6bRhI0V2cQ4PZjR0he7bJNa9THVR
50BiPMKM3gh6CZSs+XJvKXKuyrE8LCrwychw13bOSbJ2Fuy5iwJX+kTy+JJh5jDF/6ELfxgdy/Hh
ChXG8U6Iw3pjtjLFPR3lTTXF/kw4brFJ2y/+2lNGg8bsjDiN9j1Zy+tVRBSDrXAp96MbEP4xqzFh
59o/qQhR9+YUfQE2QyM8cFCbjEdIlLpybYgcZTV++56psnQExcOcrtob36M00xvlkGJWGIPjyGh9
jOuDpxj1yYXsyBJeRy5cKZy/u3meOwRdWP4REjTvlgYYknFMzGzGHA2ihULgzkEU/ceuA0nxl5C0
Bwwv1bg9vMUWoa2xFGmRdH7iGNA7sgHNzjiS3DVZPfZ4MoL8v2AizFnaBiwb4srgJ/HafRiROyIJ
JF9qHFavYBtwDITrztB+WsLxn035WEYswItudIybOe5djnIrcB+xVWjqn+ronbd47E1fpm3RCUBE
2L47DOEuIvm+8s1Ew9fac7snmLMYuTTeqWDbjIoyD46+u8gO2ojyyywA24R5G8QsqeB9yM7fYtXd
VW9waKD0ezKSr9sGPmkBUGBBtGlDgh7h2w8bJV5BMqjwf5CQxF7WLsE52pDLM47p6RYa9wg3kLFb
cIV1D8nFdfT0zo9+zEuebZaG6UHG1a9DmD/EgmtB8Xo59QnDAHBnFUQs9pLaoPz//fd7qM8JRkOQ
23xNSUJtCbXS9G2wZbWM1VuQtHcXuudSyBaCD/Hby3/OVMmzVuCXkv18CsiijFBEYnKzFmiGAy16
NYPR7uzc2vhYwg8HuEgHqKqDhTfoj8PZjosqvPnikbIJgtatyKbqzyh7Le6R9QPPsgiMx2U/oot2
E8r1F2fQh3xUjzR+t2A3UmdJcL6tY634DUaCd3NOU2J9bXG1zST8xuXjT92VGP37F6oToIK5BrCw
tJx8QzlD49shmgGOwgNFOg8Sz8K9hYTDSEXWoesTqRS/8vR4aHk6pDh6gX6AFOsHVg8ih1XFL5BE
+dwpx3FmRY6UZvpxclmbb6HknpKAiTvcuE8ZF5dhQMBZOQVljKjlrx0FyhKhvCvBDCPaDtTELr6w
9RM17Cz3CsR/mpYshpw9ntTMvGFy9RHKyGkrSyJ3Zp1RUDUlgr6kC3iLNbHie7VYtNFUq4lgoRP8
0E7lhpfYxCSyHYeyml6f6NNe+LphfUkOYnXs+RuMNOJYl8/Uug9N2ewfi6ydcj+88GX2Y4Pzq0Rt
DwyEkFjzs3dEUDxYsKdqMX2Kalnnj1sQdtPB8O6IeBsaUIPtbm0yNJHeHODdjobW8MZg9m8bmEEX
z1EtRmCyfL4B7w6HS9+0lfRuYku+kdThVDWevxUR4k0zplmCzz3KNrsmvliJRDMG9d4OmaO1a1BJ
tKJ6psU5dPXoRbdBHSP4x+WNAyGoXgv4YSFbCAK1JOzE4s/SN+cvKgVWRyJzt6rmEXRECI9hNK9y
L2JVzoTo1dW1i9Wc3D/YDE+gLKHAmrZNE/8vpcZQ7nsnxI6ogRDvD3WgLKlaqD8WkoNWJaDqT0zh
whMqaDbCZroG6z+jPDpy9dgjMVswuTw0sgc498OhSPy7JsAlmjAB362XTkg3BXFXUki5K3OaP0HU
pztJtg8xAyG2Of0DANJNtwokx+Avg3srjaEoyzBI2M3lvkYTX/aFAyx7HCp0glW+O5Z+2qeRsiv7
N6ZV+yoZjlEy/X/Do5eHOvuzwNmkUfDpwJFXfIObis/AVp6FHzcFY5btzezcDD+g3Iox3K+jN2Be
3KX9Rv4j+LnBocVgnieZa+w6sTlIrDa0UWz56w9QN8noiVMBEES5c6Kwc544iXi3q8dKcMw+olKY
NCb27LkJXBwEbS6tAl9Ki9+3Wi6ZBGquQyraBV5jddwtAjM61/PzO9AsLhZOrVZfr6hmhFCgg4CD
uOBjznqoLlE6tnelZxQT7mK4GMMyE7GYNPwJfFfIY2I/QuDcimy/MLeohODUUlL0TMsdDi12NVjX
rRYQou6X8jUw92Xz186BlvENcQDaI7E4P96y9zJMZMItn44Mnu6F3Qojl90sAaImHv4m1P9gUc9c
dyZpQBOkv2CPp67lTL26E3u+SjIxifGvS1OQiQ12O+HwDn/3EHLOBa67Swd5Mnawg2BcBAZkxBgZ
ILxMrvgNVNGa7Fsjepu89L5+W4y6ML4zVA2+tJ3cFQW9RX1iYY3r0zy1rg+LpRntONXzIb7Phsp0
UeL/DjprFnpBg2ZuKSKYpENo6nCqlKh8zkiehlURisFrOPHPUFjxjfwPs7VVkpWJclX2jVh5yW4O
Rt2Zfk5zccgUhB6MxhftNPLmCwl3d2++ZIbUfaUInSgQ5WEesSWsJ1sqIxdnsMOTImpoSEhN42Mo
ELjXULsw2ycdyMiTaLsFOueu+p+vR8Jtll0gsfvqsBnBQotI370Qy1G6/P1setyxzAJSgjznSJRk
lCLAxRqAHDZWTWAWNUZ5qZedk7NzjtJfUPf0zNSTzn9bAytZhYwdOpxhXL27rWZmxDSLPnxeyBbK
B87PvDDSrc5GhkcmSFPBUo0eA2vFqkG/GIq0lH51b58VEWM0HFSGS9rGB+8UneKGgvpAYyzgowEf
43g8Kccm0dCtmoOQIUgX/qVlFArFWMFGTVUULDjDOY22nUa9aygiA1qE5Aa42L0XOPHSjtSG6h9Q
wa4Mq4foiiXv072FYrv+9WHAL+acll+D2IpIAjjvg3ceiDl3nsRLtpCsYo40GVLnab+IHxWE1OJf
dv6PWiuWEEkU4IlzyGHjlGVR+J7w7+IfDAUe1kHiof6gSpo34LaStpjuMWRJI1Ldztj5BKTQlWSU
hNGsRbVqm+NqmTckhHKByBUF/a46KRf7YWnUbQVtwJ5UaOcPqEpYLkmgQuQW2MjQqnyThNzHqA0u
//mZmU921GiTcVNrYN7ahyBmeaPqQWSG8Y+d4CfERrH5dDpUy5tYgjDyXWgIoAyAGo/hYhCj+LfQ
LnFfyJjNA/ggEnnO369q1IUJtWdGuacR+FNTluiNbp1aO39uBqt1fPtig1cxBpavOccilje+wuct
Oi9ZzFn54wwjKlKuktHubdtX6r1iu/aQuCwXyMVjrp7YIg+dzXNREwleZcqk8Ua+iLtIlK5e6uYN
I4tgdnCmD+Rwy+GP3nrgp4SgkYS73SzR8NncXFvS44FsuzglEjbh5PZ+AlB9wLLm746EQ77B1WEU
r+gC4YrVkpcHpZzGuMCtZUcyxxdgL7e96jRjl6mlxzv3r64wpm0/bSS6/3GLme9vOZagunklocAR
IunGTI58YXp96RCIwb1PDsEpZhNDSC99GLHtJr87cYTxvNIH8w7GBd4sXoh/SuNbYDO7RX0zMUxL
36Uiuo8L91f5hGMZfMSc3PsWPb1hVCtEDk1IUzMZkxytlz4U+oN4sfW6w9tVfcasfTboKJkASd0B
Xt2Uf5su/HB/gJ2CifMWVMQ57j3nYOXV1WcUKhXc3mWxTfal5KdfORo4NiXdwmodmQeB6nZfokDG
Nhs9gFm3ohe+3FbBaC7qBkZXGil8ZLUGFqZmeZlPFnWqkpy8Z+ebjCfESMAbFHzgxP3tV8dpYgpZ
Yg4Qjo9GXSvDjsEljxr5DGZHZ24vFuhLNW0QSFMA7ZM1VTu8/XTw+9C5bvLVLRWx0vcGDZVe8jot
AtUfq4GGUzpAITxY5/vRKJQZZE9qdE9Y1S4uWcLGRX13ZZ1v5ZLV1sp/5AP5EG2aDZRX/cvqJ4iC
SDIT0ZbKBV37A+mEyrLXV8VmttWSYLzTuFy9uSuTxyeQS8OzW+ok3NAArAk2Pak/br3KmXRL0JNG
pJonO9VCczPcPO6NaBmCGPLUnWeBdm2Vp/67JjvIIpsyoXc/Z5r6w4sjQMED9BszJqIThUoqN7QT
6bkGpPmrPFXooSMV/YSSVIOlWcWt84pLtM2pY5LN/2ppZKMCUjQsq873i5zTizynkA51atbO8qvL
cwHqfrk9NjAVjrU+wUijSu6aRhYfbfCS+EkweYABrCjk/7kwz/8GtOnnz1FhBOFJOfHMvKXGh45U
MIfm4vIA7HfMVr9U53sFLVtkll+9RnER/7Iz33uGly9etqTUjcAmleqDwzkEeDUcnRfVVFx39GCd
JAoDEm/x106MF41muVuzNRnAIOfuG0VM8tNDWUZAyzplczdeUxDMgEvaz3OJg6Hs0n4PhtvO8TjV
O7joQEfp8VemNXe8hXa4HtRVdKUPj7rp+2cP6bdzrNof1iy8FdUDbwz5VD+HTzjwJqY1+v3h2CiD
/NkSRFo/Q8eMdbpNwnziN4TYP5K2TxHU3/W4OkHHyYA9fJJzWeapL8J45Wvg0eeS++QC8UEZo8qt
LQNIm2kW8+wLPgGG3oxa9TWxzj350pWcQaq4KrJEWQhWtCysZpnu9hgEdCAEqT7DuOOdyKc8qIbt
g+C52LM/14CxSXrurA2Nw1q9BnfZJbovBfyrGUfeMr7Gm1cVSWJgCDql5q9SdGVFPGHvC93gyk9Y
PdZc5jtWrmSBGoYyQz81bH5wneabVF7CB8HXon9bXQBiampcZXv8dYETNcF7n7sB3VdSPdAmKCAE
E53puQiudaoefkIyeUmc6zsObTInf1f+ucWvw7YQE1zXdcKT+mpyC3mhB2+mnmqAjrHfw2lvAJEd
VyrqxKXq+k3d8W/x/ciJmV600cWLxmwPDj/N3nYbk9Zd78Fq8j8SF4qlti5JbE4LP5OH7DZWWd9/
augjOxYLX3hPtZV+uCe2yq5Otc6rsD9kM2dhmi+Irvzpsd5KLm8YS1ZQ+CTcZAWVJJzbJInbyyxV
SepgD6JtGzv85RZ61LNGy0bpPdR+o2vEcPxHcJ0E4DlO22nKF7fwVdPGXUhpqaZ8A57pLnYS8/XQ
isipOCWA3fmk+JKsciEx/erys9h9gJwXwDnTswVuEhUCT3ALgvjCtCiw8v3N5ISXhiGpMoqNcY3o
X7BJRHWEfXcYwEK4zXb1W2G8+L2BIXhBoxNmyDJyZ1q2bnwu+eJCxUySWwPP/WH6N2+46pyKy9Ti
0wQsSVgGwIcxjlX8+HGxg6HyiIVzkcejHcsaqJrPy1WYZYbG0C5ysEKjMiTH/SU/Fn6p+95bNxSW
bsorSh7ZlEgReD/tPBjVXlwUGv2hVUIcn6GYxC6HhPoHUru+diWxhJGEg2GII7zWgnXbB3Z3dYTC
3ABJ+JgBOiRsE+zcqWVMyM79bJOpUHfveRXbj2q18YKkgsz5fFGbRHeNFQai25ejcG5Q2TK/Txyf
5FwtZNf/EbIOD7wcq5Gy2kD9xrOFR1U31sDs4C+Wdel7lrhDMNu0f4AQ/nYXQUwp0JYsm2iLsNCS
gN/3XJ9UZNq0GQtjcjSPq+o1HK1KWjSmSpEw4gPGQeJJSq6Ike1SFZBo6Hl4s9l9hfSY9tkNC0fB
e7nahBWnhqgWftDiFfL7qI+kzkH9Q05tQEZNtpBA+zT6BM2aOnN2HbVfJQLO64mcHAI9VmWufXFI
L7pM3fp24QxgM0xMSzr4/lgoqQc+XoRPmIs80OpNxDGLgMWI0Lih2pMGFlRqRYHSxKI/dhR9S/nK
kAoc6Xzs+YvZXRkOZ1fRJeq9ajLb1QCZkvKp7y8NBTsZbYt3j37rJSY9Naytjx0alDB8Eqmr6ci9
erpxtVgMAEoPiReMxon6X4C7sSUZW4bw8pg6MMkR2rIlH+mZigrnY3ctTPEEXcj82hNNhqxAswTL
dSREovRkvbT4OO10DetXl8+c09Hm7HnR0YpzZ47AO3j5WRFGzM7s0b9XqCQFarrtk2vKLq3nZngP
j7n5V7FzT8yNcbkI34ktWeW+zdFkzCeiWdAV5eNCyaT1HZMBk6VK46HBwHVKd+wDxo4UEPxfFRPQ
LpqhV6bA2x7H0sJ1BctKlpeJWFkLmOEoUf5oO+0kHYeynOB9G676OChWnEI1lRW6nvImJaj/2SAm
c0U9lFeu8HlXjYcaKa2nT12SaNAvIYYFuSpQHoHu0Q/w6tYUl8GgBohlqH/wTcyt6h1GtntsRvt2
JBWNdvOvnpY1TeAPSpevOtQZXRQ84u96H+wC0pKpHJWMDwFX6w/VEipZrMb0vtmHVJ4Oaz+JxX0b
vEaHynPPY6llekZFjc6u3DCvw5s+pcNp1UoGdF23IsG9wQBBWmsq4JZ5ju+YIBszbAIkAVKkxr+y
PFumugCpMne9m5npxQFkKLuGz3y8b4zvH+KlTEvLUTMBKPPnIHXHbumiJ6ae3sFej4rmfEgcqfbI
TgVebdOXQaLJYqxdOKNN2PkVPG0z4o+uO402V1Spdoy3Ttkul8anAKt/cKsvp5RrF6EQwpFiiYmD
EqVTf94KTFrmU7HJ8OINvX+2Gt332HP5ZGmAuBS9F6MGE+UZskvHyeiVVIAkaRM7j3cG6SG0sUoD
aLdqp8mI/MPml8ACzbVI3zsUB+/HxAaWHSS8O3N7atWWJuQU57VlPfbeTJjeUMBdjmILkOcjFs/y
W9uk6l2kUmdedBP9qoOeKCrJp5bnqlvfCdTnkUW14FlVAypl7CMCRhdk/I2akZkWrd/3va+0P6YF
PuD/mUM7UETsUVPqz8iMo06f0N+yLSrkzdmJYEOwc5yyStOJV7mrIN1Cuwd/LIEKS/cvG3IliiHl
NAZFM9ZBqAoeW1ufP4/tFoMZyRm4VCWz3nXdoZbOOpHFC77HDMYcAj0+gnKKppsZkwcGKg9NAHsn
LSmQBdmFhYvUXIYVGBoqol2ZudHm1K4+pxSkiUNfKxF74H+lxqn8l+Iya1ksH3wobzH0k7yKcZul
aaFvj5UEUAjwRh4zt6jPF1lYao7NceNrUylH7HvaOB1NfdIS2cURnZjpK9LX49D2HrZgzF8A5LDV
nhdIZnEBm6oI5NLiwoCO4ujPbQqPlAdQuEe4eSbYdjn9AdPuz35WOxaH/uXZORMJgD7tDZDJwFHd
vieb0WUI8xr0iXNc+O5tuO0q5axOYvvNhO0xl+ZBL4rO2ledAcPIS08fnGbt5F3RLF4hsyMqg2MG
NbW0yfYw/nla6tXnU50i8EfKsLHQPFRk14kbvqL4gZIGIrXJmsxYofvAs9JoK/ZtKdo1mTs6wWkg
aNMQr1LaBvFl+OeUJEq+whP092Dd+QehYWKP85hnHtjS28+yIciKPHr+X2Q5s70EHs5MUj3aWO38
Ttus2nj1OC76bnXwdgiEW/jU5NxNqkueOH0lVmrvojgJQUu6n+jHqFSutq48jrNDsl+Bt+meX53D
Vs9V/g1erd89OgSCEoiyrfA4Rt9sYSap/Kj0CcCdxnXTTYQa7w2ZZBxiZlJlH96O4EgrnGAHQq5V
fLDo6+HmxxdKZOg92NZTHKDL4bCVHsiyfuO5TBMepcsHibj/HN3rIwnNa5/ukJq9YyyNhY/FXoFO
f4XtRFHL2wCP4zJF3oslvGdYZ5dCzoVNBOsPF62Ffp5boLpauJUw/KMXe+D0gP0L/lLpYWhukYXp
I0SRmYWt+9eAH/4NzKdMoGQnvaaew9JScJL0WKAkN52YXoyOIvHPQYbTaYxP3iG1hp0nKzQ81t9/
RKBTpQZwhsxF/oeIUe+k0A5RYgkawlhjmYkBUutJeV/6VHqKcj7PZE4AOg+LrIXk0sRMXkEPK2IV
k/6FzRyXuTyG9Z+Vc6G4Bbn/ytxAl9RabYCa6BxMDLSxgDx8n0DlZb7ilseijz1yFy9oAze4uLV/
KUV7TLg77Rwa1FSPMebGcRvMyv9yRqL8okorAnyjySwri9EFwI3mN+p7SHwNLTWSq73A/F6t3dWD
b9Qdz7D1df0B5aZh27/5lFc03VxvkXzhCZgLKGWKnUDCYclOBkkBJfFNr01552JWuN7gdnhSfSjh
FacaJrIh2LkngXRR0IZTKufIKwEyyipyxdZY4DMRDokBI4wOkzgTWV3SzYeiLY4o3N6Q1mvd166y
rbvRbpi2+Rh6BGLhs8uz5utFvg1Tpp41v1kLmaYMJc2xz1BdFsVi/s06NaVPEVIFkkkQepQza503
FOWfEbiuLALlkHlEBoLrBi51OsI4HYLzvRciTL2Fim1/WXclXUq1gyzLlAfcA4wtJ06HZfAGTj2v
RHdWudKyAp7JdQV3AQAD8OnDWLo7rtumR4BLdu96yo6yDbn16xsXLyxHxhWS0fs+sMvu6A6ULClK
7HVO9GynukH3bRHCOA80MZpwwZ6Q+5BSKjDpvAKOlVg9hdbPJt198Z2TgozP3fFn4wv4hLH8SuCw
niCRyzWZ35nnnkJ1SR4O5Qaqe89L0Du0excRIWvI9Dl/sqWXAkgRpTBc6p6e0oNf4wZzFh0IENeA
2XsOOTJaaHPfWotOk5AdlwieBSoyVGJ9sYo5A9IU55qOlm9tqr6G3znP4Afv6I1C6CHIcH75DCJu
vZeQX3qer9Q5X75oOAo2hJK9sgUsyNTynqRQIIZO1O73THPP99GR/wjbJuuuV3138/4/2cTor7hf
BpiTLyn1Vy9Bv5/6iWUtvVfS3cE7pgEvFy00blwQHPOTohjBwRO/JLyKaNqWIP/u1tvVtmVJmo0m
IFxB96zh+TC7xHy9DM99YmEA03uDwBETBdOyU0TSmiOhguwC2QIKfkqtooQYw37n+lCJzRgcx6Qx
84KyfKtDnI80fCQDcJ3DyCT+aMQCR6TV38B/C2A8g/Oog66rKDYquJb4IoiNe95q5RlWx0Ut51s8
1VEikHU+ClBxYwZgOrhmWTq/qTOpPUUDuMXw25eTHc3ZTJjUXP3fwp8R59sdrnVuPDls2CwTtqD0
t1JfPWU159yvHXDsS2rPoqbL/putpNLTBsnmZCJtk0xMRu/0RSStddL2E4GDXrhlDlNJi9vdfXtR
ZvYtxSj8e0KfhX99goePkbioZhIeJh2gyyH5gclHdLxNH+CmS5yQsQomTbhWbAiJfbPPaVCoEjGC
OFTb0HCJiaR2GIn33bnd2i6Utr2v9ODimETWCygAVdffWuF8ZoWVoFmF0BaGjFMXnyqzxOIAPWp/
I0RpEuwLTQnq+OwR/o0vM/riCBN5gXqFjKECcLp8ZWNIbtZJHFOGCom8w9cd/SAn4mxufk8Eezan
DbYUcpv5GXzrepvr+quFaAH/Knr9pxcbbeGFCdV1sj1D3Uatbwz8nWKxqsDvabS7oLpAG89wNApZ
A/nTLI77zaB3CISu4/wgQ08S9P3BbJ2Fd2KburJwHnSfUgApyTxSGlBZtCctoPFEJzfclQPKYerG
PT6jDmBnmAYS+Y6lbtDpNcXwqHEw5E7SJp+YZiqo1OtU1idOaUCtmatEOOP663fw2Gkm+fb/DCs5
dJfs4K65iqrYgB+NvE6OFzlMvl+KsYKXwEX+/Aet3W8zYQOMnQSCDYVv8OFFRYjO877yeG7uYXsw
mJVXB8WYCouIQEICAxZo9CU6b5tYwrKseXDWV+2dBR3Zvbk6zKmIc8D1xIlsKrSOBmC3NEI2vcLC
BdO+Cn2SQHMbwfMP8HYrA7Yg+9ljiGmL5q0JvropifyW0o1wYocGXdLrSZuxVTWPzbYTxeuwyx+h
tkXZHJIwh1NhA9FEVeiClDhS9VvvXBlkNTmdwdU2DDQHRSa4hkPqcrX2guwbmns623PKK7ERE06l
nxj7Qm+1t6H3R5KNHqiOFm+hK+wMt8SOGA4A3nWtUbLbl4kkrMm7N/6uNKqGU7PrkEM3HIAhUg9l
o9PqdpB9DcHhBJJa+duC/+CJbl0Ve/9BNHOyqqwyIoT+AfIFlLpebaeb9bngLMRGEGG3guiWzawK
1S36YqJp8udzuB9P3d1H704RRA4v/VJXWku1O5t41JgrEukAEeb9EZuuDaLK6i0gsTl14CVwZIxF
P/iDfATaQ2MJDJzY/wPNhwru1RATsaHNVEjqNSLv0yDkfkRL7gObABCO630per6m6+fcxYS/AcLd
RhB9VRLV4AmG9+27ROOoVItFxL723geUORkHPU7CAdHA48PQ9LMMKEoSdLqhzK1LoJdGCOriH921
BopKBVEVwo7AiRWI+zyuMhCDqNlksM6w8/Fsq+pb98pmYGZDpDytESwhx0wDffhp6NQtBqeYoVgK
xduXFCxVvFDjyLEwPEmZXFHDtBSzu9TI9RDacRQhmiPbKaKN5lgo0fpHe6y5ahYC0jZtSHnj/WBV
niS7rQAQZn5SHZthlYFVJr7xFnKeVCbr2CoXba20KMmhGj6ePZKH8fCcJbGRAu77JuhSKRfGyDcS
6df5FYQQ1ihwVI+VfQPi00lOBF7/8oi2D7mJ9FQSLBnW68Y77HQO2C2i4xyPkyDKvXr72Y/3Ro8l
ABHCMIEPvzBmb0SG0On7mDAOgptmblSgS5t2RzHCRJGWSy0GeqyIVS/iNv/sbelI0j6eOhPkLa7C
oCimRuKdpZBzycZ+QRfUcbgfDGHRBMfc06ppQiUU4h7lJB2KX1olMxot2Xg9O7aaqmMiM0M/hawQ
WTUrtFJQlkkWI0TS0hrUEunxk3azW0qzKcXN6wXLy4HQAepIoLptlB5n5NaPsntuZ57Jd9F7G4Ue
fIXkSDN5Zfaz4F40eIpu7glxZxtGUpp+r94EMjyZWa7pgg/CIOycwiPa4S0lgZF9zHrb6CqSFM4u
cnp55oYGaVEi1MQg8I5S7xxr5flyrXXoROKSNFsImxt8Te9hVUq6vjR8utMkpB+SPY5djTyaLEse
GZBS5iOx4V2KWTA0nMmNjrHA+b90ocS8mbX2LfGD15PzXr1WcdZ442kfAfjv35+FJge5HtrCkyID
HfW00M7G23QWGI4/XKDzjwOIFN0b2ciTconwPMo3sd1jY3WWcsVgCTICS31lHrW5inv7OtPGpTQG
YSPYhN/wR9yeZhHeKYGk7rTrepyATQ7yXouo6rTcsEFfHolSiAwJtNavf14InLBkSStYH5SC53Gq
A1ME5uFI2EekzDHcphMEMY5PC0mqEZFzya8pS4c9VSkIcfJ9o7rcAjs9NhqOVtwsltER8fNBp6O+
RfyvmlakwyvAdTaklc7E9e/V3H1ettGrkztEWwJ9XPd29C7mEoNWGyWrCh7H3NFKF1e2fsqqzvSs
fD+7eNZxEOqdalaGdyR+gnVbtQGjbmolo7tai28bU19iFHs5JxSF1mDznpFVLqSHyTElzInXo2E3
e/bUwVP/LPMNartA+oQ/eCrvg/sli2HjaNw++ZVHoLkK88pCi4TJn9L7OC2Wd0LDYU634eBZM1yS
Cmhis4OG/mDUTRRqiAY1G6kviyVCk5qvAxgxP1ZBK07tTy4GdULcuoBoR9q/L21uWF+sB1tsMNHC
MCDaxx8It+E2Y3QbkFIW7e7lQ4gGKZGgder2hQ1QqJSDeQGrLHrmQlgt77M22hP9iwYr+YlTv/8z
VVIJGvgT4ZAppry0ik6MDPQdDnnoL0uYaCda8Sd9OOkWiRLPvEFRbB/expo2al48gln2Gzea82gT
pvTPAlyiVsPQ2KQXnUQYEdetJwRAX1SAm3CHy3NqD6iyu5jpAm2A3VlXq5Vxlhu6mxYZcvK2sobS
ooAk94wFuM3A2S7rBE+MECR6sTI5Yd7F3of4+qu9q1GO0ktIynkNufEXUiyf3Mu94a8iWIrcRmki
2nb8TqohPSwBjsTnU6g9lZRZdDgB81qCUFj21j1KY2+LZhR54RWKkMP19PI/oTkp4xqlEnZTWOST
HtgGXNQRICGOpeMnjyQuI2H6MC0rflbEzs0OGDvH7sUJXC/OBQPDCKB9YTKouLm5og7ZpTqRge1B
Ai7zqwCObna4lxRoZLoVfs0ugsHWQyQL/LqDGH1aBbopyE4KUueIXzGzLhuW6Bs2g5K+A0I+Z+rS
Rp3p0LrLEKGgecGWXGjlfPUllnS2vPeyMc4ExIFmmNcM2eRhMBLu/g/s6g6V7xHRZWDE+z+R++1v
knbvQ73OjQe9aY564aZ3LNrEdRYxxzR7hieiHIN2hOicsnoj2Mz+UW4OjEdI0+D4Xn2wYWk5AGPd
4n1e6TA/893y8Kgp/LQp7JHrWmKprKqqT1CQE0VhyUSvl1bEf8kGLqQXWCjaGRmZcgJFrgdfMlyJ
wB3TZpzPLxT9iUVMLrf1f7F50r9XqlDL3FsJPqJiw9nZEnsukVjSTU8FZls47tilzrNup3TYtPXN
6t65yu1Wp2O3SDYdH/5xAdJvmLD9gYsvu7oKJjXN+mEDeK7MAxvSDTTXimRY9/yQdusqomHASwbV
yH8bHpcZ9yo4nm4Dk3iSi5F2NKicfkVAggaSexDAKybuazt3GO9KOk84cikqKt6RVt91byAR4pB+
IAjynlXTdBSkpvg/FFWkJczjWAWWbXkwexKszvMF/S/o7zzAY4JsPfJvpDSVz4lBgLwSqF573DUU
bCjmOxncnA+buzWxL7nxkdhon8wVinp7y+H9XP4EotbhMRd11f2toJeNYLNlg9ScPvW1L44/zmrG
pFA2facycnxlIeiius8bB2ACoFdEInfcFQl/3zctsGIz8nI86STnBNo0BNJXLLzAEVdjrNOPrbLA
ls6etrAAtlr/art8ILANh3s6iocLNLB9PZ/AyefmhQWkH7TepI44Idzjf2SCxVKBxZsYu9aILnnt
4DYsdADf1AbBPRl2FTnvwbpLUYj0Glq5lNXUOvu4sY1djwJWiYgyaV1LjM1neUUOMTvJK+7Ngn8R
HKNZpfhf094364IbSg4nFc63YGtOIJ8DuDSpo0uIKBs1Jt83HoV4ztEs1fL/M+TQyO04SROB+TRR
f3hol2E3n0elgPcf1ZCMwZp5KK941/w2xEPn7wQ00qk6HLAMFtGjbGLgZH8ovHlP2eXezhwarerD
YgmavCXPtmp8tQznLpbHum9mJcPu4wuo/BOfcPofpGvq36dg3hkZyoMmPjeUSwrkiMa9Vo0Z6+ms
o2O6UcKQVcX1v0beR4tDg7QvHZyYaaTr8R2W54KVAJKbmN4arDz1ioxDnEIgKywmelUoCYOf7mIl
F1aWAxO4tMmtNSXTK5LhhQJlVttFvLHuCBXq4uNSqW+v9veCvE9b7a0ffT/3Y4UxOBoYkDcSA56i
bLXWil2XvFu/En1O8LjkRqm4deUSA9CGXdWVoUnhy28KZM5w1o5xMACYJgIZ/oY4Af0LOAzWnK6g
P/TqL3oDm6WY6a0+UuKQtsxhV7B0y5om3Ul3L1tpwZ4lWr5004KFHnoCg88YPr2npLFiW/E/JnHr
POXso5jDgUbUA0RYPnFXHNpff4oUhCZXRo7F606Gb90upmoF90XSOCSpLWCBBDRZlug8FBEwfaPs
rYz5J0pmbZe/ljStX7uD539D/2ymDV4S6pJN7aoBi5htqFTcaJ3kcoNleJha80iLxPCkzbnD5yUU
HYdCMS0LxI//JtNBlkcA5C4CZTPX0Tw6xOn8fpqHhhd6j7do8HoAltZC9NBdnfFotyEKWl45Gna6
5aJmJJ2eED8TPrO1HVSo+UUZ7WNrSPI/OY7AEcIc//kGs0fWJYkDrLzAdoN8AQSv2D0eOny3gZSX
1OKPS4HiU1FZOqIJfMco7eKKJ/6IVhFSeNbUm8sxDxZ8LLbYCgX2Ys3+YlWYp3WlaMwWrB2lYg2B
RB/bG/Lujho0lCLxGHiaJWnK7ZBUIB1yDp10hD3v3T4dbf0XYwj2+uPx61+2xQ6u4Nf4oJkCGGsg
B7wpz25ggButJx3+r4zsGol1WhTq/dwKTFQyNzO3NR8Bd2eTfj+Iq2vy3t+ZSKz57atKGfAM3l2n
ijIYb264tdZAGsbF1sJOL71rFvVbiOSSE+6SNQkdGoogKGtQM9EzCjY6PcRtRL7hKJNlLiGvrCL0
psc74VxURqG98hilULIRwPYb3pZUvwGojJ03pKOveQtfBkVJNZuqY5hO4Sec3QrgiCryDlK6lvP3
4j8xaI9gEx/hDFwY53Hvo4JD70RH4bxn8gzNViG2y35jb++frGuejPKDiFnpoh9kYkKD5IgrA1sH
NnxIDDCetoVwetPfcBWO+TNhztHhxm/T6nIRF4DZQurNk2/MyaJwVPk5yiQnzqb/3j58ANcRHY/H
Z7XnnT+7G/zAkGpTYaqfw1fFGC59pvYfvW+ygyZdhhKpXbga+rip6+o3rzD4lBWJrLLD/9H7e7M9
yK9P7Ik0PwS2q7CxvrMQr7TkNCOFrtJFozC4azLLSXc4v67G36GVq36qFwgJuzzLaqb0qOWZHqQc
ubVP8jO8Q3FpbwtGkwjtAUrvlCorUMf95oErAfkZE4+wbwZ3c2gEWHxwsGjwc1OSFdP3dPRfjTYU
j8boSni76kb1T69KTJi4oEyvdqRkgUEBl0sYFs94JCPOzs07Vu7h57as48TPRCsrKBRaAzzSidqz
BuuLhxRk8OtwIIeOifLlorQThjl958uqZ2yUEoR5/OZsjXXT5+xkQxccVmSIHse5mgyJyWDuFOCy
Tp60FsaSXEK81/DTqGr7idC85Agxo2XfLSt8c1dMxxyoBJd38NQNzQGFh6OOGsaaIA3MlJq2PNY7
5UCUib4d27r7fnw3I/MsYCSK3TrNjYIjNL/fv7QId4TRTB8Oqg9F2ytUSTbxS6GSgNUBFI51Ey04
6rRKBLizNPGgC90PgPYLT2gMAe6fanoKHfRjedjHi0JWrVEu3KkRWcIz1ZsF22Dr+4AoBjoE39xI
5JNiTA6o6xM6SpkzIf4x8KjDDTrUaTofHUCwrhpslZCn+xfa/R2NKl1Rc351pHj5aLK/TfwrPOO8
9jQFH3rfZ5XQ8jrXCpbsJkWcMxpfia66VhOizABOeDLLPSrkksSuolBpJKE+nKfl2mnk7hqTcxv8
0SypUMjrqP7yF/W2PYRpVf4R6oEdTMsVzyD/XEib5dP5j3GXyjHW2SKoSMBPDXZvUJTacEw2DPOa
g4PUH9ACvnHaY6pNyLk07RkN5C+9PuywwPshAr6TiSmwRPuP4aYF2zTEW8Mm8N2o0Dcy5V4KUhNt
KGQ/O0yMk3pOiMkJeRVr4qV1AKKwYtE+Io5Of+uXDB6o8j2zn0PY9RvXG2fVX7owk0LNjSqj70Ii
b8hIa8aWSK79Jx9rX/jrmqg075av671mn1RLzGoZO08AQYYxdeDj/yoDMi4VicLN5dLn+Bk77dr1
U0fFw6Q9gU7B/QT/G8PgTdhxadLaGpxqAEnt3Bdu/FxX3vyY0uDHCwPa+9KWE7p9kkmiZwE8RvZd
0dtbfDq+xpa++eG4ZI93ne5VAk+rwjOKBLTWODTHntiHbtthJaG5IMX6nl1FyT68bgRypXbY1wPp
cfZBXtG0iLy+yA9feKZ/PK7GySUdSv7PE/L0xXg0FIVPcZtcEKiHg4DHvI8CWr8CmfLMD8FV9P5p
HZF76d/wPYNMHKXC6A30wME32Mwsvqa4E/yaTNgvyGTBpyrhoB3Bz/ilU1LcfED+dYdZIjBjuopT
9GrzZwL8H1NNi8GYAt8maRYL37P2tHc/dsFBaomChU7TWUlANTZ2DEX3JMhtnOCqycutX0xZXZvo
n6676kuQXri1viVmkd9CoUIUXtkrc1VpN0X8ft0NosVQN9Atk6S+379EPgP4j1c8ONRPLFMoF5VR
DRoubVWOYWKF5L0fTI78dluMllsJctX3CQ/czpb59Vf4y1Bq+yRDXFaKuEzascAqlvpRsHHoOH7X
e4KDw9fE3XSMe2AkFhSHe4YYBSr/okI8XEzAVvDSurZ2uQerhXQ5Gob+0784XYTJtMKQnoQwIj+M
cBX27hoEBVUHZwcFzk6mzG5VUMS8jJOzIqE3XJvti5uuMHbKo9mGAY4JREQ543MeWCoqjcikeZda
SuWcDs6A71vt5tbQTqScDPDRST3vQsbMhsKUujhCbYpvYNI0VV5iZbnMMUxmxiiuA9iFHZDovq0G
0D9BScocxkLYFl+IRpxlkSUTWZO4J/lBMmgQ+EsIPIQ6WgrKJw9LlLhK8rn+2aoHHLIVwA+2PdPo
dcd7/ifFrh+3ICg5NU6OSirNrDNonWMK/mKAtuoS0TDl+bdhj4g8aN3vLg2nFQwaC2jwzctbhIy9
/W38in9wYjXwVZWbGnBkVKL+opBmpzAk48ZOoOIcPucU4hKkn0cqI8x2fAtBaJ1Mi6MNDoWsnc1f
BqKyJdn5w1wh3FCZdw7Hop1TPYrrktxmDgwqOi+uBIBU8ybhkI8a/tcNJ6wBnNgjLSyeDKz4LF6c
IHySLaGOT5QrZBW0YhZZVgb+x2wE/0/q5md5TgZ7sEXyIgcK71mQz+pLORM7R++Z7r1m4gyuMyDv
kf2ptORSgxR8fTuo+vlsoQsY59RzadBnE6mRCEF8haramzJKjRADPMvL+cxnms+PkbaWD2w1hD4T
TICekoDHbNBSN1sN5YWWchtRduq6NL3mHC7WECX2xEmj40wrWJxRh2+INoNIqoudh4kOZmfmbCRX
4HtdPIOmgAlZV1xvBnIRxS/7UsjwaOUxfN3mdpoSfsD1gA1608E5vpFiBOEyZPVvDHTNN2D66zJn
GSqkp/luKuPOvgxFfG/27EuWh3hQJWlvS2+oCGPxFur0adbkUSAouyXGyFwD3xHFvh+YadvxquOb
5PMakiFpclijJPR3W/9pQc91qamZATqOkKG5slS2EK4xIf9G1jOHcgYtwNrDalYarYtkVZentB3o
8OgPOt2+13qK3MwnITCgS+Hh9u62EluPrCwWyYuO1ZrudkB8El2EiBvOtL8AEzuY2eEoEq6zmm0C
Prw/j/hf/dJU8K8IiVhdoQiIg3HDTHQYLQGfhNzwVDXIs6zM32Gh1hatQJq9wyzis3DLrRuy6dev
K5U+iKEsZFakx3+JNpE1Y6XVaKuAk94jS/70e0oa2ZZQ90g+XBgtwheKiQK07PpnKEY/Ar0/ynBz
14bYz0xSUjhr0O1txj10KjWayHUAa7jDD4alf5Oun6XG8OdyNe18H4xS4fb/MhT0YZxaIOqwWXsB
mXpp7SpdnzFC501EP/Y4RXUgFL1iEUW4z/28uoJB2v/oA8rs5ybeh5xCTOxf+QXpB0Kvzrnqlwhi
K/QpQGPkUMhrsc2N0jW8lt2yRRSt+jRVV0UmDPKX+mSkTsCmfiFgn5xKjLV8onVEyUdP9x2TIeW5
TzsWmX5rtZ+moVzd+ZjPuRISIN8xGzGxS/Tv2os3obUjlmMuihoNoo5tl9eX87+u11X+DqcaNVUz
ckpO6zeGh5zl4DOoAqxO/0g8zDe+KvI4sEkHO0pNhObJiy0us/+US/rb19gtF4PQCeLRl5LqQBNa
CMhsby8YR4OeWkGPCUS4+eri9XVJ3kfgqW+mZSIVT9tAtRrEyufmIbSQB+B9hve27WziN/qHmLjx
b3cBqCFARVMq+kfsPm26V6QmNx6lGXAItnRfY3j2bdrjEoA73ICk0Rjj/WsoOU0H9HLFesPhy8JC
hZdY8ukX/pPIogJ85D3NrQtDfzb9AK5qeYIBWEMAUgxazSfoio2VU6H0NCUhA/jH3gUe7FPn32gy
0OCGLEBNd7gCGyiojOlqQbOs7XiBbOglFfzMY7bybW/LuaZjiUHBQhNLJbuWtg6579JQkRDa8AYf
KiYSefdklBhtO0r5s4F5/tT2XiPao0nOsRYMoAUkLeGLAY7b/UrKRuwNsdTDuzxlQ/muIAHU5IDk
zwZQOjzzBwNNQ+jUPDaE56BDEu6zC82w6osVXicP1oQ2CsFxACeVsRjww7Vd2Hvkfk/wpv6eZlO6
yMZn1SuDcrFk/iBT8fHdzfzV7vCKiJNLUMK8MI/H6M+JG+AW47Fz26S6bDOSfEyRvaCT3YDFm3Ae
rjbz+Srn/l7hKM8PACQAckLw6iQGm5CczeTVuniG3pOumv4dXdnbv5YZEZlISUaw1la1eTY5T+u/
9Cc4rULYJvTzKhlCkzb7fdsqF5ChRZYMpkz+V0BIrFJ0tA+AXC53/Ma+o+7K2cEQnQs7jixIUkHo
sMDtZ6Lxfg1ixwnm6uxNsp+w9Jp3HufHHSMPOLG7uB/FTROJI0HGNNeBrVSpqw/+g7V6wVOGsy2N
Rb83OF3vYzCLNTHvS5If9aJeNhUjOc/XfRmXLj/PTQzHZZkCX/WsFWK//z4NEMjzOAYu9LvjI2de
MoWEdFVqNK4jUxIQl3tkuUH88w9VkOjPsbfDVKzpd5jC+LsbjI7tZdzL9AhW9upVokNFsSwbiWRi
07I/8BdyzP+usc58XgSNtpDgTBneOqBgqwv58M4aH0qLctrOt++gs55gYLdW3pq65cGUFAWAgzSq
IWCMqOlkQDmy5kcq5FRk3GFp7LyNeAE3pxtx0WkrJLEJqo5mFMZZ100g0O9Lg0/e3Ah9d5tJjy7D
3cKiNfXWj2OrjvBd5tkMxYOplP7VtQp8nk7Jfel0vWlk/FjiAETzGnsqBTkbfnUc2nqJFG75R22x
Ua8IaU+mi5AwK/IG2n9YONA8VkLt8cz1tHq16wXDCtWaak6c6e1fG+vguhNxpDrKBKQHVAnuohBk
DCDWufDh1IpqfUDY2nRoDaZ/4LO77GD0mEsBDn6AzgC+fqZIINg3vFhjPTiMAI4HqrkfJj75mttk
7UB7KT0zhyiTFxmRHnmR29nrNT4yw003c04hzsBBQpagdsp43rycQLyNwJ3LGl2EEhFT4X8CAcZU
z9vQ6fV2Dlm2GpTX1RjrXJFXjdOucDP1o+Vm34nhLSjkkl8FyF1i0aP6MGzHko6Q6FImwHk4RBSz
ceCx/59eo221nw36Y01+puV9a6f/ACo9r97ZDn1HOj+NQPv01/DafV5hTfQtrSM4BHMpFgNvzIDs
QEE69C2PtQbAxVAVnSEyhYUP3jD0+6JWHccXHtaxMCxo6rtlgH4lC7Ms1FmZ/NAYh2pDF9uHW8wN
Bp5mHWTNsMNlBSHG0WG3G7AfbsdjrSsEnZM1tJ/xekSAae8IQpA6+G0hgBfCBwdRgS0olhAJvTdb
3pM1eVeXzrjmGOq/ReBeb9WnCD+xLKJ1yv8Ec9CWc7dxMrsCqBDDpQr2ZiikZqzk+1RKD+quXozJ
b2qUX9UpyzDSpKz7nzoOXP5RT7uKMJ1wxI+O3rFNJ5ToRZNKMFpkEBYFeVqYKLdFhFBsBjJgzCvO
ooKKnHcMTdzt4ip5/6795b/EqFBowR3r5nUpudB943cKuaShw+Bef6pjsrYpEsvpFNFKc27dclSZ
+Snk6ZICJ7AW1CDnbsUQKhnCVG1ODAcUQDXk1Zls6A95YvomByu8T31FI4b1kJ5wEa9HSPzZW6FV
Qn9BC75yADOPAY17JgLhqfyNC7oun2oWImFpGLyk4q35H+Ne67RcIMiE26RTWJgcdEwkyaCk0HIH
AqFNTCBTfMNOd+FtqXQMQIRkf/vrtUfUlMyoB9M1ZTjNlKl5QCMhAyq481ik5BjNcRWURR413Gti
ot8RZQUtMqQ8u+VYhos9+2ewFV/yns3jaijEoBqwEbFSgMQHjs24pIJ9hp3KcuVCKGgzWFyNl0Az
hRyEvlJyOyzpseJJv4K/nLWxLvys38Pd8QbvTO9FYs38xbgElEqTAJI7VU0GDUG3pDsHnWNAfZMD
GJbYxmn5V12e3C9+byGx0BY8SuzHTh2aqFSChJjEOwwzRMXTiCODHm9SGfB5vHg8DkzE86pJ9JmQ
J6toZZppp7N9BqAS7oxtCMKaVmBzKeZnYhEPw5Imi2B4fb2xfE4yFAvss9xRKBy1hV7MRoPwVPtM
Mz4eGguYR2e30xeW05eobOdU8QO1Ngoel57UL5kBzyFrnwg0cSEbyqd8UOEwZrnru8xo8SLseDs4
GfraK5rqSxlOG6/Q+zKGGlRFdFLmNSoYUruO7W+w/mHWEeifxlSOc0uYrDRY1uc8voXGNd6lKYmU
pIp5l3jNzvy9WonMn8YjY60DNWGnpRuB4a7xWl6J/H0jqh3v1ruUozEXaYivSSmZd5mHBwXAe/4Z
xiyAeZWdRLHD6by0zpS12LbviovXk4KlPGnms7uPVE7Z4UDRcaqUEBRLfZ1X78BtFxM62lZgOhTL
m+4mlHSZ4ioYUw7Yt2WjK3seB7ULVmaCI3fBdoMtkifd91N2bIjYBp6ExAUST+ylzLyU/wCje0LG
XxCQKBU8nwNJ5SzryN+tf9ENWHmfiVaQehItdz7wU2dWMELPHmt6S4IDhSzSjVr1HFIKVMUSJjfj
MNvNIBCe0yzHgKtIOUef9iwCinkkPiK6sZDIxom4lbykMPDGO6Gwy3YmBEiHxe9/yHpuwZ9klx2D
H6deNXW8NaPwysGl+zSeouUfy5xF9JDOjD7srthPFATDKdLlntEa20UcLhNyGv82Eh/cnYKr5Lwg
9QbyfYEInEwmQ0uNz2K5IDfkZvRIZy49h1E+Nsb7Br0uSsDX7AiIYcvfdJyRYgxWq8LkBkV5KMkR
Lrwf0JT7WNnr3YiNWmdXVJ87UFuAlichWWsrx+VrsVgmWcP2Cs/XbZ+T1RNhY7eA92wZj9mBTCdj
JKh8SMeynIFsf5cFKxNRN9iz0r0JROTFE2QSF9sIv376GpgghC1QlMRitEvknzzJZQtFUX8rs9EX
OyGRBZWa7VboqAcxUFk0Aowu4hafZYAT+cxXwCJVJTr8SWqiGaCZ5htam50oYa8531o9Xr4gvjCM
WTi9o6YDLouob56BEcFZoQ4kQn+fzX/u9sVDTXXf27IjfpINb6x4cEg/0ujqZ047Bd5lNphChQk+
rSb7A/Rvvzdg0eQKKYu2XzbpJLJWMMIZBQ36ru55GzkKLPy7LSwZhQF0HGe/PJICLRHDVqHuUM1m
009CF5CDJnNttXJDAUbC93FWEjNgapplgZK6PN8xlqY1gjdZkX/LAQvmnvlhapYpHTLkYgVhMsnI
Qjgx1CJ2rW7wBU1G1DrPKEwnaM/XBwLRXpalo1NWX1KoAgBdFjYB+5Ihs4J7KaRJiaWpHN8JZ1Mg
YQlu4Bxazq8L2pk/7qPdtPhy2Aaf4bDr1oRYe8Gz4apN+Tk5Tq9K91f/BJgLI+32MAxuCOTqAq2X
06RUhNeqBHd1XdKqQLiltcl9ii8AGJNKL5Xshgj2esYLG0o51CqgDNiWFWf/auQzOpL6LjLtYWt3
bWucNurMgUkg7y6VdMpxrJOPJ3lMbgSqp1f84SW0ur1krSN+g4K8jBKwHzKzVe5kKfc9Ty9FXdKn
31IRUT8dvpwy3aswB6ZwFo6ol7+CiumLyuX4ml8KP84WYwv70VSM2YcZnK4dICD7/WNRjnmsMjz6
/g8ozo2fLEaXuWuXUbBk7pdBucgeX/XXXwDfrPgNdMj4u6HVwy4SrrUpKByJeHfqOUCNHSUq63S0
NPSncg1eJhRx6gRryhrchc/vd/K4YGJ5M158PfdSInV82EKMVhLas05ZvXxrpSsFt2MamRHeaKhg
o6NBMwEklPXxZx9T8sBqafGqxz6ibqHUllmOoyIIynzoI7ZTUneu/gt7fP/OtJTKtPl8lh69CitY
c5U4hBc+Nb8FqalSegMxhA3dSfytDQ8c/rUPvnhfnKavvPIZIny7exMHTKBQh7chyccm0qrYb55g
jkJDkxfYaiIo0B3ZCr5gWdhvEZGI7F5ekVR6jT3QKNB3H5SrOXob13/CVhtB9fgEcwyb+kZvGPVN
4tdncnmmLKi0VWMQAJkF2TNz91vKWmRNF4w5A8Ed/4yfOPHSTuTYhsEeCTcH6oM30WFhddtfWl7s
aVMUnruheVPWMIyVNmZT6wU/pe0HRamxNk4oPoHHCah5JGFWiOzq3Y3YlWKi3ViIfK5tJ5Yxusls
lBQ659N8BgqaxlJomXau6w7Nr3/t5hbxlhAofcKo3wbq5Rm6mjJdDAbfRSeNwW5fsGuPFOe3NXa4
TmfSzJM8Fspwuj82z6rvKDsXP3qBVeDymKOM86yh4k2tf8ZBTD2Xa4PVzBWJhER/yGmbL/KrgChX
5+dHDfKeR78LVT4EFuQBcUcNffK+0C/cl219xJe90TkvG2nLmKjL4ufXpoktbY+kTaKrRgM8kt1q
UtXpbhLW0ocoUuEyaKECn920tH9JwN4J0jSHkqz/5x64j2M5ccmD62rSqURa1Onb1oVlPqAQRo3c
QSwqPSlp9qr6d+DXSJe4+b6cNHAclniK+AUjkFxvUZVo90twv9L61CgjU7edh2vwItwIMlvUhohg
wx2SWVn1DUtyZMzt/so1w625Omu7eo3uUvUaxsvpI3wErZUraGS8qH93jY9JhJ0L/XVAJM3KVP2/
5M3NJFfvZDfhCmHlBvIJhK6uv2AUAR4U2q1AScKDevY72zkeio+QyePqZlowxJ2VXeU6H6WyEUUp
Fl2Kovjqrs/0OskENDGEPh6S0j8KmRatHg/CuKiC114UR45mEedfmWsYTtCVaRD90eBqFiB/VLfK
pZtasTJwH/wjuTBxjuJZ2QmG5mVhSI1sz3htHBorqqOj/XxcE8OmPACTmo0hLMd3V7YmXs1wF7CF
fNsg8WIBTt396LwRw59FDqtZXoszaERKTyOBy8ax4kqtIW50+1Jm0VKCBXfRF23VsnYJjb1DBFNd
Cf9PjGtlZVz90pbXQocCYtwwiJhPxnZOv0zQtXroxAtNIsrKcsLGJ/HtRuwAQFaqkRhx4HMQlQDF
nnwZr6rzwX6MUuYE7QLKB7w1UGbhAQkqW5UNlm+1Nexkwie2Jge0t35XtRASoCsgwJWKk9PbQcdU
K8j1jHf9LLmGmOXKFSj1GaliNI/86WhgsoyWHkRWkBK58MllJxwo/RnH01R/FI37xSSCBsZnFXAa
Wi6+HxUoRkKKv19+EbjfzeNSuRpNNiAAoDFS0sfJeVd/bBY/DaySHhhiXNIuKtilgvL4Nb12O3xG
rqlmylUYWDJflZijWzCxDDMKpzCh3soLcGh6zIZmtbFZ7IZqKbofhr3GGe+CwrICYYAqP71UFBTe
UGy9hlryV8FLGqrr9Zt2bItO/qwWvQgV+4qU91B5aHAzGc1g/FR/6jS3iwjNsZ+ymXeQt3b/9G2S
Pxx5aZrxSACp1SLxLFICBvEsvBnQwv+hohLL8a0aJUtANmT9Lkv/MWxWFULEJa8IsZRc32edvHTD
sx1QyJv0LJcMV2S0mXP7uA7eRLZT9pEK4zpsRgdxIcRY/V+YlYXgNW0aRKiLiYOmOVbgKxttN29A
Pm1OBum6x8vxKP1ikZB9F9EMPud2Q9kdxLeR5vTbTnUI+veWPRPy7RQJGPyG6AKHHfA18c/ajTVg
O7kgG1JI6ShcDWVPdUdjmLmXqGILjM6HPXSD5e2ss1gWKGlVZKjosfNivAdWFhgiWC0ChcEeLglp
gepbgeJWCIjqtcKmZQ8bV1rPwSooczngQ4TgAzpXhx4Ux9Q77/psC3rO9bAyXvw8mXokG+CJNNDV
sgzm04kw5aKL5oAVoJn9E3Z4UAJvqyP0qASnak2nqZuqpqwh2oNg1Q6aE9rtZK4US07RrahexjPA
C1R3EzRSssX3HTAIe3gingebs0TkfwVTBfL6iJ09pI2Rjw9DmtpUaK3J0QrUbwm6ET3Z8STcpQKp
IeUd8+iiBu9AMZ0j2EbdkJgY0yR6YcvtGvF+/yuTLXH3uJfm8z3Nfis5XtafuptD2BgtROWVC+K2
lgFuHye/HGlM2CTcTRv7Wxg/XY4Dp0wqo0mQJ1KS3EOVIKzmqVENcgS9EWqEs3IH+s8vvTIYCeZu
zJacuww2Rvf3Py3CAyEMCrEFTsnK5JQ367ixCsmnWZ6JDRBAmLPyNV4r9oGBFEuRC/CFvXETvLaz
XY+MgLF/MAM9B4HPLpNOpmEtHHtq58lkXm04kqXGo8jkXcfkV0HJ2WQvvN2aARZI4AykGni2hCX5
3/DJFLOHcWKELGgzRmOY9nm/cTwJ4FmI4/Ln6xUSwFMWItXeIv5oS5X+NZ+6tGTWGxsJy75K6yu1
PM0/YeR05NY1QjCbiDcZBV0Dzp2Huo5Zf8yJpeYPsn53heBrKzmzicLhd2LKFby2gY/tNI25VnjW
hdgkwQomOG4BmPqmNC/niIYQerEVpdG++mqcsGf22lfM3o6QID2Km+Raw8zxUjNJ3s1LVH6SDO4K
IFGr41MHSj5wytXnY6nsgMSRFu1q/RqXJ/obshiRO2c5SXoP22AWSv9PB/pGb627rKz75x5N8kuj
MVJJ9ONtbxMtwumkkO3vrUu1O4vNRJb82zUdsiqwnDlvBGOQ6fqndP4hyXCAWFjyGiO4Eq3UHbV3
E8JPAmtvUUwToLl+Ra3AS/q4vKjN20nGBK8SeK5KkabKuLffywftqtDCwNTsWeWD3Xuf/mukMRmV
7Ynt+5yD3l4VMlOA6MWUHxE1XJSSUASvnARqm6CmSrniWmdLB55iukdI6hEyp7hbkdDG2XDQReCY
6SktzQu31TU6TgzZn+bWCtuG0Pr2Nt3a12zBRDCSZVkDC7ZaNl08VxZBtAjuqXka6Q6RW4e8o/GL
PDzI37/NfzMYQzDAVACc8i8ZXSXvsUvE/jxF7KSvTbqsGfKm4gX9LkTrAQHoeLjAPHba29jtmIsN
m2yIek28Az3o/DhxgKNzxd5xzvW2dzUWhtoCQZMXHKKQGTAoeDrZN6YWj4DIEEBbCDlhG+Eald+l
JqEtu/m4Rdm43AvITCyzTdgdk1B61TST8BX3e1lCl/E7UtItCFAFvSzsDhjDDk/xn0XoYFS0XCjQ
5YfRlboYys5XnEWNknpAT+2d6IRUVHfVPYWYVBm9cp+gPV/i8D2vEiKZpe2FGuk/fr5bzTcLHDuj
cL/qeImH46b/JbWvUZGHi2GkBzBOH1jNC6EoOJQ/MfvHtAiREf/M3Dqdg7dwS/1ot6/KewZcSy8o
9awLkJtv1BMg1IDtqgGuCrRBAjj6ysD4FFMz/Ho4vW622Pkd79d9OuLtc1ahPR9oKp505n7pf1pW
AcZhCaT8LudIRnEz5MuTWh/mugu8XWH/0M/uxZvTnnI6UnVgHEbAYXoIEwQ7WlJvgA8KpiDnEWjj
a/Qo5ywRwVMtngP0OUSOm96S1Iiq2FBo6iwM/at+CC//+AtPbLCd58aazyfsXwNbjksiIWzPo38P
k+jiYgZk8Y4XPT2xHAErzmxlge5pvRjVrUa8hS1ZbnsYrkQxWIQInPJZ2I4BESugPMzNMTuIyF+7
c3QJisHFWbjGdA4w4pyZ9RfvVrf9RdUzdKrNM6a0lipCoFBcp8AbNIvajohHBTsoheO5sWndHHUT
nPQB2y0hzs0nhqjwznqqf5/GkO+RCH3spKgHKFHiyHtLysLIRioODR8UDmnUOAokpSQgQUHc8FD8
k7squCuLlORRuRmdvM7o0tNMyWEq5lSnDLk6cOhZd6XIG6GqxweYqxanbY1mlN9NWTIPRl5PHjNY
qAbp/5h2mLZvRf+5vYmDvPCuOnASAAvLI4BxQtkmZwB0r/M6V2Pyqx3W4Bf+6zCxmpLxSos+0SMy
LljYDJI/MTxgjhM2I4ul2WBsPFvWfSHexaYG6plmQ/8Lqrg6Y49u5/2bzSVe/3YRYu8ByZMnk/8G
q1dJcXb4mmPTv/5Cr9EgC7X2u0H3DLYnOVNEK/+SHkPhmPnYmhA9mRuZ7Ujhm6dZLM2/xIRvDJTx
t92r1p1WlnSTG5/kxaIFPSHihST5z7JAOFGmX0Bp3hsHogdwO6oHgbt6BMjZgv+6DWPh7Smqahvs
1FWmsQYpMtltbCIHIpft0JCv8cNhp0pGW+RmkjzH/Iq0OSEcBx6Hl1rNhw9FPI0HgimkPnDLSSpX
ZevbJD+E7HCsX/NzucIS2O9dQN+7lpbgsWFwoFVSuAZjQiQhlc52EzVyARRsRjY+ucBq8VOT477/
JA5ubs/3ru1+HQg8p4Cij96x1CX/oCzu0RzQ/uO8NP76/tiqJd8nNa7bvZJWEdRo85oBQbkeN55c
/IdE7NwQKRuoSkJsZRcxKex/ztyOGz0Fptzv55OTkVzqaJwGWmlSYNcUhwdZCM4fqRa8xLPfwnEZ
I+EiE22coCjimVGsF1RdpeXk7nfTmei5sdGCMAIJSrCj7gEtnzr/voPKXrhDoo9xvSQLCP0oNHZk
S0UqY+gQK+hDNresbj/hxlayL/+CRrwlRxuxWiObLYFv8J8Gqawjir9t9O9ndv6kwwDnUBeWkGdc
1hhGN6Z61OeTq07lFiEHWM9un7grg95C/aAlt7O/tz+8V8up68TnAtLiKIrd75DIxJ3OJ5EDlL7q
yb9H54/LvaLgOPM02mSl7i7YJ/6QZbzDp0Ef+JksAB2GLshIM6qOQgGi6dLstjuU9shWa9kao0gt
34BzAqSt05jTyQx9jBqkbWmkKEgmOcOsoikTTOtbDN3XI36OS2hlbzyjsZIfrm5gHPniKjSjSSMq
OYQ6w7lh0Gwf04xj1kNS4AwlinbxG2k+34GOJilrgzgl+JU1SGkDu3OF/wgDWoqVfbuZtUQrX5N3
sBdQANOulCakbRi4Symh+4AnFVB56CrY0+KrvUCxzIeLkC7em5ChcUPFhI6cbDh4F/km2wFZuzzp
zawFpK8p5JIKr6uql7ON792o0ylol94ESRS4N0jNKmWA2wFBRWV7uXnoVOIXFMidP4i8reN9RaKJ
iNoQds60+/6/hW1R8q+sRjyTH8b9ZSaMuokaPApESeMJPO2zoTGKFsemwkr9qoosTUh1EBz0RrA/
/aH6NRQSGid77ry4srO+rAf++uTwBCuSGz7xwwlc/clXxabcoxnBVHoW7M8L/bYlk8eQg/nSxVNY
zRYH7w2fPLXyGWDm6VEKK3Pl6prjRVCqc/3Uf2c6tngLQUbiD3PIduQ+x10yRqPjcx79Qg4dv3zA
Ash5O0KiQiZhXxNw6BaYsTnih7P2aBULdXi+WMHNiBo9daWeqSFDAVluLx3TsZ0BoS8RHmiM20F3
Y0CDNp0VZDn58U37agsX36rBcNyXIJqoa6UiBtxZjbbJcLLeXsAPoSb6mielw6H3f+fOweqyAV6X
033CWoft9sxkGUb8HJG9KN4kADfDbzJS3PxT7mC6YMQtXCXdninKYQiL0MYWMOnSlwj32NR+2zBs
g8TZt6lidC1uu6jOrI55Zk4/p7/2NKRSCZiptyu1rf6kHCa05zoER8ubRV4rH0OpqX9nQokfYCfZ
43Lcv0KqgKTmDMajExnuAGvyGHw6JK4NyIB9RpBlxFjrpw2Sf952uhAEaV2fjBNEhEm2Jgta4UN4
lUEZX9ztQFjD9uSBktMQcg/qVK3bXc/XgcY5SsKOYVwAwiv2oC8bhI0P0wa+uLfXFxcvKShiQk+E
pu69v5TEtGoDXM+StpEczIE0n7UdTl7S/8tSm3thY12Ppy0zEbCGtIGREKlSnKwV7K7+MlhgVFHq
zX9GgOTiKfWTF+lKfN7kM5e8aZ5f9Xccz3VtHo4YvxOFfP0oxxYZdTGeKsAfRc4onimZVsL9INWC
YHW+06dD+6i5gy6Ui5t2balXXMI2E2jPlaKZ+pFco1/RC/5qtK9soQx68t52/ceckS/Yzw9LAVal
uy1A/e+XfrdgiZONe0x/7JiuCCaKx2+75zKgHyvg4beJnAyE9wrpZZmaIUfboN8r/OQRlgLhP+FO
2h56ljRhwuntS7xvZKJBoTl/YZ6SaWhYlbO6AxvZMGDHupDGHH4ktkomCjs9hZBLpWUslitC5QL/
YWNrgJrI+HZLK0cHXohH4X1XRhOS9eZkss8eDHP7tFR5BybYiuqZejlXHBjSpQ0D/ke+nuCQzPcj
Hghn+cRv0reoGBixBy6MKePH+/ILphU+Ja4eWdSYj3eK4KdxvSiJWnbNLeHCZpGKnafPSiPPX9zl
O9KEer6jViM5EC0iNDZIYD2ieojhmD7ob0TLzxL7OW5u/JgYnnNGaqV3Id7Q3QxDtnO1iTEZheWJ
59ddftHpxnad+20R7AGJtCzsnfxjJUAcRf8V+I3h7IVltxgBRTsdCxMTCXIyvjHlntv5tq9LTYwJ
wbH8FBE72bkmJf0oGZzoiTF0hVwRizH41B3EifDb9QrDDp8/PYCtmXMjniScZPKu87o/t62O+GZy
orx+OhxAY8wmw1Z86cIk4CsME25sci43ASIfvvSOOMDF1vcIVj+QpSBgJQwTY+xTYpJFudmcejhu
YBXHjphv9XEwotOw6CQb5FTjDap+9lVhWsbZyf9Sc4F2z6c5Fujm2UCOklvOyfQGf263cdXpPM/Z
2pu5GZ/T2eWmK6kfpxp0oULaYYPUA4pR2PqC8s/6qAqAKs/Z/jRSA9m5LdlKibZ/zdEQ9Ct0CzPh
ivFxIgq434ZZt3XtbTLrJvpEzn6zHPP/CB6yKywo54dvBewo2Iw0qoaj4ujCxDjnFC/h7TSFGZZ5
0oMBkMiDK5CrVzvW0PUWBYR2w2ii74NH6N2GoqGltucCtky+N8QMazl0Bu+QM8ITqThPPkq+QhhT
PgxsjLPDRkjUfbUgdzkYiPT3KDtWlHTRoppLPBK0lkmaOF1NYt6K5LiL3hM1eZlBi660X6E2X2+g
j2XPRPMqHeOaB1Cvhegut5oh+f16CK+Hqu+OPOiwf6TPx2sD5s5H7J9MooAFsc4EZMWDeuiwqtuh
7si46luHZclhuWH49zfXTgVNpEEPGoxLUGSc69RwOpjh5VVeTcKYZltWoZLkcPa7XTQm2buI69Fw
P7rokS33PxmEwVvaQ/Nk7a3ehxo8EPpPzxaiXvn1pZ9BAseV/4llZQK1sm4l597jVrakV4re4ZRX
Xc+4QDf+fk+R2DeMsrBQbB+L8e9KIeqoXIRLW5b62f1PGFR5Nfu1dKEJJFcMAYQYyj8hNB+Rp17v
qjvQAk7uEiYHXvt9U1jb/bBhhz0IRJCOJNaIHA2vtm1c3pX3VWek9W6/x0BWDeoY/wqG+Oy1eXLX
WAPl2Dwo6GN8SHdDdzDKjjByT0VBlKK8T2ynzAQnP0Hx1XCScbV+InM1Fcs3TbvhSQrN83DyOWxH
zlzUOMSa5UZeAawgxp0A2BuN/b5hOhO1FaoQk9WIBAtLvAecs3X6O5+o9Gd9ZMfc55xbwI5taeiN
xalxx+/45rRc3ceWgpQO9MZ7Ig9mkCOvgMH4KccvW6LyXyiTFm0ffNF2KP/lK0isIHb8EDvsTYm/
QSZrNGBs2kn2Ataz/LqcZ6Qq10qrGtTIhtw5WRZJLGl6IuCoxCXWA521druZH+67oIfnSXkU51go
KqWh92eNzwWwnVyrVw4ZbB0A7F6QDgKr4FuaxXaFWvDZELrg0DN/fxO25zZJntY4yjGIYBNtIPC/
fbH14mQxa+ldkSkAZcz6kmv6we5Ex9VjBqeagO+w24fFqNzK7DlLq4HQAeSTds9H6zN6hmJvbqFC
nLxe/Rdp59QtA7URCT5COrE4D2ZTJrNwc+juLW+b+zKg38TTLWVbuBXlS2u8Cqgc1Ij1ucV407Wo
uKam4womiyHxXNjX0lYO/qpe2eibIZUkWhhR4fMhS1VM1shxpzIRQwPkoBevJLDyvd9cLwyf5iPs
Ri74qPsokvrpDYjBxwTJohLxrZvWLTrWscPjNKu0oKUqQT/DnvhRFS4osn9F/vQu30Jaqm2eSIJj
deLSkQXNe39DZCT6n4VZ3FuxgBp2ce8FgB9cigpIZfguu9eS13CE63WZUZZ7+5UhTyJvVE4E/rcD
KlvpH/z7RlFbdEIH6dj5oO8/DeHdiZZbXi9wJ6w/1T7fvWiP4q82bdTGz3SUvz9QRbFGwSlsyCpR
ey6BSMil0TNC1lvN+m/CxwSaPiMdfvbTHrADvov5p6x0bdXM5YlWmbRYRLKAkjEzhbNrICw8GdQE
EAms4M0dFQEyqNS0HmB5MFj86d0RowZh1Xnui2lyHfcdOPbSbi5JbA/Q8uVKTSF1JCZve5A7KGZC
6/PbT+qltZxMu6A0jeVX8qHDkk0Hm8JVXvyIYV3IE2oaG4TDCPV3M8dZIgzn7VDlDhfU7Rr3Hs5k
ZTsNMozduEuGZJx/0g6txpEQT2wws8foRfPjAaVXRWzAPYq8qpCkn7hxtnwyzq+zgM/ck5a86Qre
IFBCGmtbmEF6S1ZkX+GSC2lvD8kW/vkXjRorAN6J1CnKwoknd+yUJw7qyeB8kAwhk1bzdwZdpxkW
NvYSG83pEb/XJIy757MAEZ6a1WJHwO39vsatx2UDicOXtxzGoy4E6r5a4aIYkWUU1z5M/+FqAV54
ou92jtYBeHAZm2eiyRhyVQ4QZkGlTNrH78T7JtjW7+pfZo5691Tlhg1vJd14HwKScHwl7lUelu6h
AUIZ1H7GlMV38iFQ3eyWCWCn8U/CfBTQLaknniLtkV/ffZaKWDqfz8Ut2u8EkZl12bdjHAig4cyn
PxcYHF9snyCHBODMAMFDNxYV/gYMKrk2WjAfbOXhHNWJgioP+8WhEVrn29Uq6iry0VfgC4OHvAxj
n1GZOjug5mi8sYvSm7qP80Wt0cx4uEbBBGP6JFsArcDzYX6vBPJx94w3YnoeLDAuN9m2rxY9wCMz
ZzQTK9pPexF3OundpZ+zTr6wkR0UyNbhmk90aBuJkg2tBpObnW19Dg7YbYCrACeEqEi52nVTBOnJ
vy3+qZIiyq2WvlTxFWj33n+xxpFHKigi+mg6wPycFcBXzjMtnhOIZkmTB/ciZBEMkk+GvJ6InQWr
bEd5QDXYPwUv4yX7pkRyM4v98T2xV4AkWjjVi+hSNeoF4wgyTMygZh0FsZaJhfxKO84lHB3TzmSH
PUVWmolNlqCGxDnr2JCeNWP5cQhfVTVTpfaIbboItcgisvy1ywk8bwp7SA6cAINuVMw87rekYRC6
hvgNHYWilDi+Y4D53C0eSXUSGNOFEegmeVYJE6I7vOlZ4/Gt2hnACmj8xibMZhc+MFXmiU+YPj2p
a7e4zT1R2mzJmbV35lHn0NML2p5Zz2DaoMgqMlsoIM9qAoEV/QT0d9AYTyinG6gKNg3xhvhQSIbF
l7Osk/Yb5ShSSxSgLDv6LgtrtQ12JvmqPojLkvPQHW57dcPb4YCGUmsgntnMSn3/p6l6mlBis33j
kosraqXsv8490BK8Na6tXeqRSOKoGy/LqfvGW+7CgrKWkH8NmE60r9J1zHPJWh+jfr1m4Wo2o47y
jWFiob9easa0jNxjSn0p3x9y0TOOPMiMu1+E/5PWjKs3RENW2EUuUpWC+3jvIcZzGKOzCCSjavYt
cJfJy1UZcMvl94fDGghY/fqhC1nazV4N6EOXJD50GIxBgrMuy8lxtAkfP67nZus8ver0UaYkjsar
BWAHg8rkQ5qkqRE4kRtOWwABFkFOnRgncVcWIO759YWrd6mKDZ9uGTavZzeJmcBIrjA752/gPAaQ
/cqisPBGhOVapVAqxRXCOVx2S5G+YyKY7guvPOxO5m82Y/Nz9zN+hNZhmaENjHDVFNGcY401lsmQ
a9/q9vK0rAtpqNslH9v3FzYg9p90B+VnoiQAjU/4WwyGaG7qEBaZzj/XpBS9EvkrlcWHqed1ysnj
dUOX7Y0+5b7Jaw/90GFGnjkZo2zOeyLIpMV9JYJ5QbKCTwRDepjk5w/PmJsLtogvAyPBrbnCmg/c
uWmvQjNHuUy/+b+/f9hsCfawRQu0Lc04un3CjdNWgSDEXwh6oIKBkaYjLqafQkPUUG8JEecBlv8O
E7JVYcK9ZWImWU232yedbvul085XjLiZ4YfAg8V5D3Hg/M9eQVIyXcNLfxwnX4JWFaNNVkTkpsw4
exBG62DGh8U0b8ceudapDIBzw/lxetSVuA/74Dh2eOXu7shSiKvuqrPrkyiN6wMdqlkBz034trEx
pP6uobl/uMHnMOLwFwZadAxUb0Yl4s+KOdAMOZhNTsVXZs/XsPdfDZY0j5XrhJIird8EquaCwx4y
xIzuznjfFXdBrI/s8OAHzyr1BnhhMFW5TCiKZxkZOgVtFeVKfMbdFpYpVFRW38BYjVe3JKnH6LmZ
d0s8iIwF5/JeoUPzRoD3btEwI+chE4S42VNBvlohNVbPVFb3c9btG/JfLW9I1DLFzXyzQaK3+IlR
MxHbp++AXOzcTrtduN8iq7qWJzfdAriS7BuZ/CBdCKNApaHy8lH4tPsqThRsGICIKmpXDiG5aYlp
1t9BmwzXcCr1Uu8nGIL5E0DqhI8O8NBV2NNKCHxevtPqHB4FHI768XneOE5R+D85UZ53yGIoDGBr
LCEhc5BrSRzxuiMNT5ArGmCzfgdKDUqWF7CzX7Cf9a3WUPlQClmNm1sp3Y9aKdom8KYMVELDOa+j
1AdHkLFOBEv3YxyCvY7D+fZeKhvs9FzCp5CDybSKytKkM0fgdNx3fi5Q6c+qo5HK+T1NqfMjzFaw
rJS3nGGbU9DLi1PEhyzun9NtVeyrAWDC/3bIVtf7QKWxIR8/e4g+bkvDsw9IRumBD3QY8pikvBHe
mAJAhONK3QnfShUj8NyHXq3qJIo4NFvvU8R58bcDqlxmBLOhugKrwY4QLQBepdA72Hj4UFKgDBNT
5Sa46SEaGTRR4z4+LLze8s7BwypQDpgj0k269PRa6EB5R3ZYUn6EIO71hXU8lDe2u4EtGZEXkMVV
uiOUPb4N7QoRYuZRkcddqiaWAKvZKrUyi4qbxhWWUgY+IcuEc31dKF6OW5EFBug1NCkddQ+57boW
wQyrDSUzK6JwpzAY+siA4s33V+4Ve4/JytzbAp6+THxxeP2PiFkNTYQwCu43RI6YPYx2LlMl2nlO
V8W6LEWJQasd7jg/taSlc9JJ91P7UGwSfDLhQnb46otw5jLrtQTZSqSUF8qF+FILXfzsxgzHS1Z2
yYKBWTpa8no02lcGrw4opR74m0/cROrhQS4N+VNn83/Kq2LkJXCF9shmf/uyV4Xt+zz70/VdzBVg
Dnvp6L0T1Oo13UBcaqzlw+YQGp//7D8f9PFv0IA02xNzt/Wxm16QmX2lL0+V9Z7P9jlVcn1hjhc1
IuxycoidscdUM8rZpESyNzg5h0+j6jQtO4IMbTNoOZmEWXWCMqdKtHgt+tjFkVH6er33iFX+evs6
5nDykEFsfHgXzoXnb7MEzgrbHvmSjYhhSUgCBF8KPZEJUh5ulAF4C+HgUs+S9JLkj5sdqMA1zXFR
LjQQB9+/Ev7vEuqVbXIhtxLhIQ8IHgdUywaURcGw/tjdZ/ChEoeuFtmmgsdB3o/XAJYWPPA8IO5r
NXL43pN72UytdDnWmrorvRCgFlvzqbDs19pVR2wUyNfyi+OT7uN09Q5JMPiWugETmOEHDt8JVZuc
K7XIpWeMlVwoqhZuxYmbYhV7LGiqM3X9k6yHVXpTQ6LkYaTkChVnpOI3aYPJR5jYVhrEj//QPvw3
IOk6aswQ6XwSAVCWpiJ1203AoXQCIzyxUHDE2fJFDJd5UZk0vqmJTVWwiPw6j/qPdl1je2H8JCPp
4FVc5AHtHOlX8LhKKNnGBdZRrw3Re83+J2VXzkxl+AI3s14sx1OoyXnE2yPNq2GLrQOwzKgGX7ee
Fw21oDMxebPw/L518x5Dwkt50U/1lfQMvWAzcjQM+YYSU9szP734z7nbBWnZOVou+Qhqm/U1OSMF
Bd5fQ0r1z1InvrIr6f9P4SMc1welsOhVjS/XMP9PvAMyeK7bmEEadBgkdhEcIpOUn3G7fFiRKmqb
ghiPB/m/zpUba1NiNavx4EJgsG36X+Lq8SKkaF0mNju4zaScHHlvttC0pPKiP8Oh4BY/jj2ssXkY
75LoFylZ7u+yZ+lyyjbPS+LhvlRnhUg9SSuaEs2iTEZxDO7eY84RY4MLxNdAcTyyiC7NuwhCqMbz
zDHIRPw3eeYk8/dXmLkNynx1pNZPKbfACfq/JRmb9iGuFeqBltkBkkiYtY3fE5/V3YfUYuNbKUCB
DLrXk0A1ljrA5pSWRGzzqS/A2vMLqoPIwbWwQtiVDzHBOInqUGwwxOISAlyBbytAuHbFeLsrC+kv
8Herb8hl4ffUTELksEpppdEpAt4ceqwxfkcdRZ0VPa8U1Q1XnK7o68aqkeRlaM1qHiCBOONUGQoH
c/hv/2WeLJthT1GXbentEMe/FP8ZCgy8J0+c0iJHNAY+89cLkLOHjUDLO2LK+9r2JxVLSa4g/pJg
iVAGJi2VSxVlyDzvLHGQ2Vt41isSMQRKNP+Of9QK+KFsxFfnwTqOO6G3RlM6AWIhPDgaPRGfXBH+
yDuIsAwBwU4ZRJeNmiciqWM4jKoDcWrowcO3UXRSYI8AXHx4RsHeOP0M4q0ojl8vUoY3IWW+1yO1
If6rb8BGfsFcjnlzP6+Q9AFMHMUwHlLXMRapHnGm+t0WaA+Ew+LB3cOaxkcLzK2tz4WpLOjTYW1c
vCQ5LlagqaMQJgqM5HuInzhyxqiVXPSi3FroBD0SmE5YpcVVkWPHWDrJcczszJuTyMCjs3yGKGdj
iFNr/1Jj835LCdTAvF8tUrFR9Y9QTD6JSD+oY7+FYikvAQw0C8XKwPsu76mt47YT9EK8GICCBaqo
QKCaCfnl7hvwYXFfE8Z2GGuyYiF26T8FnT/ExH+jY4ewzSntNND7W0CVSGRtTLEWpOKZ0TyNGZ8J
es84DEkPWELu8pcryhblCbwnjsbAVzcbT3qzdKQcNln52B5qYYvh+8kluwJYDhFJoWiXcqxd2+20
2rXQKRKb3NQOJiunqXzoHbUmQHZaXwUFhTuIhcdBASdympJXMn+uP9hoZmaoCjtKPcT9hjgMzIq2
Mf2D21C/GUrEBr1WWnIstXvL3Z05tGL412Zqz96tbeemkNIjtMg9dVCAua2emtQmgvlZXdYRyngj
Gm+oV9kfE0Z16ix3nsr4n1oRiBM5gHb0gnqPeTCA52ofIrj5gaOceCKCFhHKs5fQma09zSJf3DqY
FMiMvhHfqDh2TqubyyyP3dKrJimmi4p5t8vpTmNWx2VbABUvAg2gjzerB0BryUAnBkcd3+VRmMQP
e9OQnxUcQngYfSL89nE2B+XkIFakGUF69bbjS/MqJuGapYI+H4SUVQ5GlamtlWgsbGHAAZCcvdkX
16YT6vrD14nlx/opBv1U8kX1oaULIqAmaVmLg9/YD9J8U+ZQw1zzHAdXgL5FJg0BNStqeTOtJvZh
Vh45GP020TFKWr3lAM0t5uv/ckejgAtx/3N1GEVUGme5SVpWy837P4mfYQ+qcwPyZ+i82VMXAaiV
cnQyUixYwC58i8+DCwik8n88O6Ji/SGtXkaX2qHdx8JlpU5aIPTO7loLMqaD7BnnhKLjSRU3Iwn/
diaHgSfhRxZmeZzS6zCV59OEbxV95GOAjwgI6fChenDhDxgQ+6mnlAk7fwkBJWY5lotQBMVd6rcU
frFLODyKCjZFXgWZmqKLk6RWFGZeNFJZ43f1hnlR1uikPjWcHQIl0eoHJCeC74Kdwmrhm/z4Mf0O
ZNV6Z39YsEW3lgSBaseFWrOQQ+JLANkGTmaL183f/lAd28nQXmjcnTv1CjBXTAAFCm0vgIOcQCr/
dmqMyD38G7PvRnbYNCJJIOzwBS+tN5TZ2NHWMUX51qaK9ndlm+lhOjXQ+ChNfc9GJx6fbvCOsQ8l
FXyCVCU0x+oVC/pHrklD6Qt/XjeO0tVZahzAEKOnHxleb77pnNKsFthKLgbzcigCEQ6tlZ0yfQtc
9owZ/PcwXjvohyDaDnfMFWYLw4MTFmJlpGqsjOhkulHTViGshI/V5uHZfSgE/Gcl7+5v8Iidj01r
eUf+JFC7KBl25ANUmATdvT7l/q2Q7sOcdS3wz+vD/JG6DnRec+TAvBIDT9Q7ns0PWDV3xiyGNg2K
xwagzvmKoOfZhR+29yHbEaW2DUbC8kIRn6s4RbnnAQ9d8D0XCqo7JsZlozi5i9ob4ZrMwYXM7gCy
THpa7wIq99E5EgYc08zGUjTpsroxZQ0BLpBt3sBDgezFV5G653il5QZ3g9V+OlMiXFTz7VHdsj7z
O4O9ITOLOmgJ45IMRN7UEVzrzFJggsToU3wiSpqmBABUsCRqdy5B83L6N3D+Umw6lfdzNV+5lKsC
wf2/ytea0UosZLGNp2A5q9J2v/e/WUlgmucWY4zKrcTJhzdTmrB9Oh7iDhPJipxN05lQEEpS5rQ/
RGkYmY2fQ0IKA3m24sde6MMBiSkLu6SgO8zbcGwwWxh1SBKCVtr4Wtifgl4HWrz94aIbvGZd7CRF
J2xgH+P3MXzdQAWAgtRQidD26JxDRYAeDurNmYGJ2lzapMr7QD2FK8sx1mMS+QW8H4vr4CAj4gE5
K9bTThyXqPuzf/Mbc2By6ubg6IOdUtAABi31LoPW/qqpqRrGHZzvdc9K2sGCkkVsg1WIabz8a9IP
4vGRrE8eHqKD3d5UqNtdPQj6PU8dT2IxA1ICTjVk4LFN4+WtBb5y4ZHz9gQhY0H3hLf0ybgOHk2p
RUWmP3hT5aC7RJ+XYIT7cwzBw99TdpQqO0Z1RlSEQFHKGNTWTMhDo3iOf/hWbK0joGL4VulJX9pw
6Odj/iuTj8dAi6P3rDecumpHwKI+YUxVua6VmCVUMzcQ2dQ89tgVUKA4qswRYuMmn5YtkK8DUA9u
8IJez5ndf6gdQHPct/WhwnM8Z7JlOfNf1zi1goRzWN/NarPbzp5mzpbAKRxORCJdgKRANjbt57x6
TCpWZniRjzd/KNzSDnPze7bK8vut4Jp38n6JkVLnMPY8XJcrqDABI4+xyEvmt30LXDNKdFf5ZNOC
9owqd/gwH3O49QQMLV/5MN9EnHJugstK6mY7LvBNmSHeI2LwiuiTFHEZ7HOWtHzGE4oASne4a9q1
uWCrYAVyAd4HAtrjhTmWInpyF6PKnahL56tVhu4yQdZtYd4z4SdmJLcnXq7Fcy1OsL9D2wNI59Kg
/VxrgDfWOAQx72ZcuIEGb6tSsT3fBGxAfAc5C2srmur7WeKzXOx1/XA0V4h2gAWK0Gkq8hZn/Jrt
+td+wW5AG2uc5RfGb/w6+wY0r5ej5Z+9NvBymoRAZEo+j12Jp0vpHSE4DnzC2KEO60C5mZXOOZac
kj3OA9vApFhMgAYxsMUGwsICEhTsMtcmvvZeiTV8bTMJyZmt71EK81J/xelNqeCdzkU/rYv/LaMx
nD7eskM9I23jsm+5RO9K6Equz5h5QLmFuQ09UPiHhKCz0Vap1Z7Uah3sn/42FJIzSi/qLG6pqlZz
moaa36WB75E8ZYLFRdVid4X5Pe9kq4uB3+qbP3d2wb9N8fChK1R/G0BSTI/y2FntjoZs28XPgZ7g
X36HbekrqNWuAy0TtELmIPt81FJxF4VIzXqOyhVDh7LX0jevrfyaE5kvN8mDdaCKHmrO/Hu4YbEr
Vcnini+cYF1I0nOmJWDr3OxXWs20Iw8m0bm/6PY5rGmbFOleM8c4/nInqAnhk4cCI7hxATBEbd8V
xEJvbtNfkiwS58XizGTt9BUBI+JgXba99yg2YihKhk9GM9lVSzk9kMPQmiA5Yahys0PX+Fey7kMU
BJpzozTxaF/WWSjUdIQYAkvGEFNqUxSgCUfsAXXO1Y/XTOu8wQFrLVQLri8b77oUS/f+2qdxWyWL
R+cWQSG/90IEKsxgWYT2qWCOGvFLOdo46YSgyh4xHju3q3Zv4+WZ0kkvBk7q8Onu2KUDwQRCQMMZ
qH0ia2LMKSCkUoKr7y/XCBmbmO0WuRfoKFrtNTXMEOkhjJ6YRwnDOGYKLtzHPETP+sz4dKXeDoJO
0QDP4LW0ANe3HfiHb+cfaKlBke6sglYBqyzpOaNeW/9j97sLVfgj1sONiE0ciBOHSlmMafDaOAHC
5CIgX4tOAQDG35vMrR/+bke6nhsl1QxiuzexOkMoKGugRxIuW7U3eMa0k/iNWx8PlpOEvzMhtE/T
LLYjdTMXwHNLHoJYSMuU4EMPU1Yjy8OebVEWuWELW1u0sonWN8NikE0eei07iV/akWKzRVYdNXIO
6VmZrRoeOSjbbnfK2CqK1FB2gzOfuDBC9R7XT5m5IFBt7/mT0AvtQPMMX9RjxezWlwZS5nzxV65t
ZGBCyRmR8tPIgK6d5YKLIGL9PLI82KUMr8+I1UcK+n3VSHWFutb+yhme7G8RY9fHz3HS6SlqEfft
TcXpbs0m7FKoktQQJw6doF2Raub2Dwas0oe/TkRJZg0ccw3fcgq3cUsy9QgJ4MRklfRvKL+nwZDG
sTCEng5ZiOXk9hFa/5Pi/KlqWfI9MF5Up9kCWBWSUFWqq5qfCTfB/7C0FWecGsrWeoE6cAZfimGu
IqxCiPtaaU4TkYBY2OZ3VzC4M6W2F+I8GtpGcMM7FmDjdcyXx8S23ON9Se0vhWSoZYVjAyfNbyoT
FamNtO4qWD/CXgi8GT3vkrVwYOToGW4gtO0u+y+EIxGrmT5k6/AqvS7CgjNndkchcZ2NX3lgHe2L
VfiF6+XMbt7uR1Owd3NVAv08dj3XD0B2IcBlgKe8C1t4/JtlOsmExBegd2Vq9Su1y/s/+hgvksS8
nkBpqEG52My7kvdx1pDLGmudVfIlWFUafPs66MrXJjL5nh2wkBLaMTxNk3ulxmcENEH7lYvYzZjb
fNYOnSWt88HzBTacELnoQP8cxdevhonHFloA3iGbOM7p+FNfeetMOitOVgpPP6G25LZsApAw5hbJ
vuVjp6mZH81G4fvVqiElfinutgvDheOBGUG/vGGwDfej4pN39kyRSyAyvBH/RpS71X53xoOCizl+
zow1ggWQofJ3Nc2Wz/SySl/30zAiUr4q/RFDyOAXiiHHQ9pa0sNbk/smofdjTNMAPWzdrrXbx8m0
JBg+kKP0tx4rOXZzkB9JzrVxggefqIryzdwfYL2yBDq93H9efLp0lF3vGB5uGtAUzRoPn9NioHg7
lXwt6bcJsy/1Pnx9W5xTnAwtgc1bIlO4PwNbsrN4url7ec7X0GHBOR0WyXCWGPveSmnSRrmQI9Km
wZYjA+sloRc5vWVOveKEwDT4p0voCm6sVQ5boLMLMLL4cCeld3iRYjUR5mhHlgHZXBhknfUIKvI8
0km/yLsz2qPNoLM40J3YrMh3sdM3CZ1Oeqh83uq/HqlyEMyxiXliwQhfR0GZ3qu5XGfQvI4yCgAw
aCrO5A//cOUu+99q+nFoxwV4T+Tzwg5CMiF5IheqD6b+GI9OR1O+duWw5qoHEc0LoEW9dU5Z32aU
vQBUEB9W5oOdRqnA/TY8R71Ik68sDFVEa/aGFRO5JKGkqM2HoloPNjjCdJbOZcXvH5WvYAH/vKa2
gBYzz1YKIhxcBqTlCPjUsoE25S5Kat0ahtnsMIp67iONJbBns+01oAH+lkC1u500gr6q8JVEno0q
Kr6gG/eM7YgtNJDbqx8J88ogCyJKQSy8In7p3uxLDcZNJXLBG9o0Yntl++7E2FmhWfjy07sg5p6o
jMsL/UnoBNkTACikjAOpVJ+oNp55yQKXVDOR4aqCSit8kN5fd5LIC958UYITm5uS7Un5UxFZiw6q
K6ZOnFjrENNykZEU+OahNv/DlbRWyhgO0hg+WN3txXWPCB+X+CoVGSsVseYPLm1Zo3myLG2+spq6
dcxe6NlBX/CrChp4WRE7IfrTzdjyr49Z3QnsWS/nLjB8CT4hTYyx0xHf71jybnZbqvSwYmFr82eR
jtbdNoY7rIEyMjD+gwYaMUEe/w+Ho9dAe4en77pHvWxFgWK76JNDpkNdghAeT8H7kCBoc09pwp9i
ELCdKc3pZMBLtYYuQpXmXK+DtfMQqsFQrXNXXlUNGkeQaLpCo2h0K2AkVVSh6xQkVTJWstv09X+g
x7sxEswn6s7ab5FdEUF5CQSFYadP6KU9JAZIjNuL0cQHfKIwoFVGJ9Z6boi5PmZFHuMIgUzB6bbG
XCbR/LVaYPuBUSYJM7ls/kLLgOEKkCOtTbNbe7aPGgssXl5ezm4YfdIYBSUG11W1EZ56v3IaXxdI
IbAlNSMTcnmg6pvA8E2FEFqsAoiIwPUFRC2NvUxD5Lw5fsqMRo4wpvxGm+bvMoQg26xy0l9wdTZl
tlRNYVoBfGdLk+Azv2Cu4IuIUaryK8/oYOuXo5YiL7N9f1PkT8yvUvoVX7+UZ3ARahU+VOKDok3N
55SwoBXluB+KrJDCVryzdTkedk4FgHXsEKjsOZdM1kftPTC1Ad2TfCo7RK7XPXeWVCu7raODDVBY
wx7aOBj6aNLdfa4fz9oaRkZo+9m5H1fYB7XA44E5bb4H/H3c8bXvv9KrRjUuUQT7EY++dnYjC/LE
l1x6pwNeOqIxjh+pPmIq8h2uDVSFuUPILHutxQwf71Z62s1qJALX8P8bJTrWSX2aXuOSUvwYedKw
iQaYVtgftOIHaogSsbQ8+avHo0dueOa3GZkZpBerpAfpkcHAGHfZ72684i/+tito873lhmBB7AGH
oARvN65OQw9U+RFIqmOzqT6PneqZqOimaOqEoqwg7ADji4AQNl+ApT7Wrf2A3+/bJmCc8ZPbkWhe
bpZhbpFzhybaj1SnzSpBoD89aIf/maGmGG7iYOcgvVDZw26wNEGBb67EhEQLiPbkDBodIu+ZSzwz
/a6Uqd9yGO01iJVl920tTI0OupDrxQDDR/z6ww/dKl8QZPxlx4FGOLPY4LRwSb9mD4bkjO5q2MQQ
DKiTaq+InuC4pQYeKLzFp7Ubfj8Gn2yxRgredfYIoc0BOyIGe1haMCE2ILnfzuKL7BdwIbceKpwR
X02uPQj2/yekkgfhjruazQoihsSrI8Y15snNX2pj85I664lH1FfGYdv5JaPCE7Hp1bf51RJfD1c0
X9g+YqXMdf/vNkgY0nPtM556RErt/XyRR1meXRZ8udQozV+zJfEZOxLEcy06vt/RFvXiqATM9ZVd
UdIn1mbAK0QBSwDRBxfPBfW/uPnylV8BNQMPaVrtn2OKKtOQmKW+vuGiqLw/Ysy6WOtPGsxti4li
27HqfT/q+A95FeDR03069vt/vWgyRwLJk31axSFrK0o29t4QocCBX6CMLXJd/ZYyHArQJ60VbuQy
xUKN1/bGoApL6LR246QFh6qAJaw3uBCIMg7i8lqE7O9L4dhEnnul429dv3upkXEDAheN/2NM8BhO
MvPF/5agZdTCU9B4ecEF/lbTLLohbk5Q7OXjr17ncED8m1BotdVxbkuGkw2BOn1XNMHb1nIbDek4
2Zohiov1LME+77FZ20IuJFf901vmkusKlsl/f2UI2Up8Hgt8ygfudkM+7l/fWKII1+a1GW6lOLZL
cyHJEEWFLGd7JRac+6iJ77ZOF+CfFOsrr7SDLJYiTl72sCMOJ2/EEu79QwX5Kyfc+MoQTS42DZoW
2rwyluKmzjeHllgm9NazNsJXc2kOHUR1JlMNJboCR1DaumGQh/ZPt3CbYPDkjX3QIx5oqIY+U3ZL
aHRzHbqvy97teY9ryQ0osOJJqdh88O11SENZ5mz7vlHvmieWTiubobVb7HMXujDeu6e+5oEZBSWS
oYdy9EWrCW74K/lFJadg/cNRPPWykwFTUxN1dlJhIk1nLOqQZ4UGwlp/64OigNDt4/MI1OjO5pxJ
j7ulwkr4OlB9FSNeHGv4azOdmED1buPxGH9RJxZG/B+vtSivJBygF62xXWGO4Vh71XG6dMAnk0qE
bSxukoR8sxqTQyoIHamv811/ufz8e1knzPUJScidsh3cVWW8PE67l5DISwkIKyeaP70SnrQPf2O8
bTzNDSUWMVzoQ4n2I/tMbaIr/7M6pFhFWAJqCCsykkDGhhN0O+HsDsJ5zIGdlJxwCVCyFmPhODdh
GhJ2XpLI3hn64Xph1y/bA4QdCpkp8ZTRaxFbPxvCoeL7UVaUjbkUBavmUNxSDvV9BqfZRyf46XnB
Ff7hPFAUf7JM04CbSOgjYRLib2NMTNnzL9Jaw0+Jar/OHHDCtyh1NWwK7V0WW7CsLq5dpxjdQdLQ
6spdtRbtloEzba4Jc/gXaYw/GIGF3/w/se0U/2+A6WFfpBFP2PFgmi1nCYquexCycNdFWhOGERV2
LpO4cAH7tzTB3YsLxxsqwDqn/E+ccrSqmnt1RCFHr6fYblnQTtYFn/qtvyaxyCkqh5TR1GLxysaM
Wd7B5H7uHbWVt+05rObFpwP8omNHg2P9E9IwZESyj3iMaA1zJPXF5ub/req6JhhavfzpqKNI1uXj
xo4EOhRyAHRFhpgs4JJYdeOMD7o3Y0s7mzLG2LBMfO+zy0YCZMIqdeq47I3mAnTZ4tUxU74m+E72
/9wo17DXKGAldR72QBt2n0DujOYEu2JZ2T/ZRfG+PhJ/jutzqebAZ5OnMh8vgRHPE5ovOcKEXx4C
LIRak2fXGbwoRxHZNeqyQT42EQ0mR7GUUukRyWgoxz0lsYr6WD+hSoQtgCjz3kvItA/0diGszqiV
JLI2xbEbvgTlBAG2pPeBgDOK6NwOjcWavtiKO2fPQo+rqYyTGwGgQYbv93vKIe/hnnrq6EcfShg4
Ux+n7uWzqOxbCW12w8l2jHU3zaUK620cy64Xa753XIN9vdolO6dFcHtLiXbh6/cC+mLwCrzYiV3E
W9x+eeg4UXshfq9C1cmgFrQWU7HD+7Pcb8PLdHNCXzvOBuH1dG+5m4rVXGuPjuZoIkiSQH81PQzC
F3WYCPhR5/ZoErz/URGOxOcPPbh7b+F2OnAXKQsCogKKbAYnQRRNWuf1MIT9XrwtTIHZ6/1XuJIu
tliNCdOps5ddm9SlqaCtND1L1oCXH9oV5Puncw4+zCIpZXAwPTGkTPQoO17BxSj1A4Ll/sVVgN1V
hkfXR44O6XzChHbnVTwofiB5jXXwu64KzJlfbpfdAjfbzi+JcB6HJLNi+j/bwjJbeY+PMUDmuF6A
f1yg8brL2Un3ywvrflxoVTWAeTpGagygVNU47lD+SkNk8/krNC1tG016C0o2U5UxVTHKmUlbbE0y
kCN6IQ3WOXCvIobDlxX9PiiEVx3oIapKX89GTJbESykyrsitWkmPesF2D1kRaWvKIALZAdKGI69q
cmK8ea9/XnhsgtzAmPTmQmffMJtNk7MM+/yRczlLJfFpIFpeNNHX6E5aKpgXFUcEDN4SRyQWuawC
ns8B+Vp0Q6mG/DZw6wUZJReDe+qIfuwXNm2x5OxCzzBG4qdUVUbO7/A/D0enrlngb9szNahqbXpn
cwNYYfzWW9613qdIo6wJIytzv2vglhRrGLc+hX5iJJjOooUn/E1wL3HF5xY7Q2H9AtyqvZLBwIzS
gW1+e7mEKcpo9be9EEi0gLVWGvEbGiYf+YbwuRmMzS4baxWcNqPXhTMmx/dGdZGZpPH/QLSqFKKb
XX/C2JT+nmK/yfXe536F8DDjp6KWsU9ZBj/lp/ZYPuFaSluMoA27cmnbUg9YXYLIlZhTZDxmicV7
X5fj8e8BwUeQigMNhKhtm19KIoNtv2bDITguxhupTFwRwc9caZzpj26PC1Sio64HOrSOenWF5oMo
jPsEDEg3IEKqOacX6wTADWrnN+rUiR3RNZAuhv5g99LRxaIMQf89flXyZcP+qqfvrF3E9xczEV53
ml9XsR+JCxC3T9xUEshqkFNAf6soRrCZbKQaKeXih+nMnFXspZWMuSD4mhHfo/cW5quCjhGTX8Al
3kEK+VVojL0FO21xttbbYXsQOAn2vrWLf5CsZMoxwomXyKgpg+oGJMLe00tzwDgppBFEbGQ+Y7pM
yOMQugmUvQXfI4WUrlafqgVaC31K6Rk8uGH+SlQ/lHWMKuz4M0/fbNdzTbRfwlRJ1diKNwMWV0vU
WAtDlbTC5k2cKlpJ+3mONMd4yEQu2H29rZRaFJTQB7fHOmon9maWu5qnvzk7TvUlMZ2jVZw1x4Xp
BmIBnMTD+qrOMHpDPySTMw7LgUZkriRelU22/XNtw0V8FeankOW8Q122Vs+l6z+pwr9ncgnw0B6U
Kr5JLldRLIUomtXQvh8GPsHrupnY/1Dt0veMo1qf6mZY/ElDVjwojt03dhaC8gxpV2RtJrkGja09
gkVABnT/ZUAiIBCSVdlEV0EDZMIWCPU9Mp/L9v+Jx2BQN7YN8k+VW7YK8lAC2j0mrRn0ytqpUQuw
NNHChJm9knEkfK22ElCYulg05y7TBp/4zt3kgO6UalpLNP18U0rz55/aKvH7Gc4rbbl2I1g0RpLC
n4N0Y1rt3Ha6ONcYi4a2xVFM69eaHrzGgG4SUJKGCsR3yPWKRSKwb56Q/HGmakDZ/XrGfRU2nlSb
ayURglJgoBdU5KLbuksj2r0SLXnlgzMaMjkXfoHmeKKt367vPjGHw0bfAzIPmKiXYVTXQJRgBqXy
435OQHqFNU2cW8kH/V/7MyaFVCpBiQLYDbDWh8aUmm9b9V3WAwSfMVvKyLX9DACdW4Omu8nKxDsf
bl0ErY5OgHx1YwR2Jf+yi4VMkZFSqq0WcyF8nknma+1XDVqushrrnptqcCEGMqc0GrYGox2T5IYI
hgTyY/tLwF3LG5PEmHy1c8NMWcdrZ+3xyjq88tJMK3L1nK5pTqrTWEtMGFPYBFS8Yc6WQmqTQT0A
NI6Mdz6AdPEHtwzujnbqSsrCz5BKooFk1QadsShdwVI+31YGJwdKUXeneLPvqalW5DNMw7Hfv0i+
wxS7IA0ncdu8AHolfUwBI3aSDDLNsMCXlxF8FbB7JeUud/cxBvPOWp+/EPCkJazQwURp/hcBhm7f
bJAvvRvEhF0mli0Yl++j28u2ix0RwhraU+i/5xkJW34TLxAa+2GvHMiRS00THWQZPwCsibIVnZWM
Y1Yd5D8hz1tVtP+ebWHP+S7ENithRigamDQ3TZmKag5pKlLZIEtxUrnUTa9GgO/XJAelK6m3iDV9
QMVkb9Fl5ACAg9s7NGVdOLDB9ROmlLT05CySSLkDstYpGqdADnEiNAhtnJRsQiK8uebboM6ftPz/
d3c7lzDDgitO9XOMVENpVZOuQvlbXsMaGZF05ki02HLHEPPA5XBE6bNe7fAVu4ErZgsk83EQYibq
B1QpFDqK9+VDOkNJDn15o7GQmrEqeZS86VDmYahqIuQjfCWGUAAUCoqosIsr7ls5Ydi3f+ssh5sA
kqM5PaZfRleXJNQcmrvGFBqzxHKh0fBpt+UawwW883CvNqZoG2fi7zL1BA8gjp+k65p4p88KP+Yi
YyrsgCHpgMQhN4q7i2lwHrdD9PLX7QyKST0eFWBQwhGCqx9Y+0ZUBbTg1IUQccjfnewFdWQ3IMwe
MZcq79Eb8tC2vihjb3yHON4klYLw+FA7OZKQ36YvpbaBEP7wp71hXzAcgxjQQRKB0VgfqYZX/nIn
5+78IW7lBYqSHNzhmPMozwtNA1MC7E5x7r3ed79Yn3DN0qMcDcFBJCFedC6oud1v54N1fL3uKJ4p
IlJsbD0JD7OVNm6kN2t57cC4MnPzGltUzBCvviEtJnkWZ77MN2G6ShlyTfmMTJpvL5pjXDn/wyq3
hP+F/q6r61WY/kpYIxRS+nNxhJzYAh+5ZhyRe56J2Dm3S5HxxDPM5dQFWrq9icQV1Gqsw2ukop9t
WZLCDYd7vHhzZZpB5b/s21r6KQdsH+ac6gKdRcWEXOQYcnS9DAKBQJPh/0IrjQAE2HCjlZ+aI356
3MDVgvjlfWXSO2+Ww3AT3QjQ6ZAfcspChSSdH2TqhtWlKRm/7g2kGyEogFTRp+iMwNrnQlQkmQbc
ORUMnc0sDkoemNsI1/Py34RbCQ2kkl66Yq/M20PJy+8X3TG6MOOWWzTRy88O7x1V7hPJt4eXweiM
8CDlUTtXBrEXhfHmGLvYkpskd1w8aotwwi8uQ+nFX4VdP1H7sW6OLk/6qZXUOPYvLYzMeQV7xpQH
mCoRA13/cPpRMFZQL+Uzpn+rDxJpp//oUunL1OD3U0z4cSubBE3m8aU+yOO53shs2V8Davy5AScD
45yuJN808UD7HatmRMjTyvQ3gvMioHyQe31YcmWfaEDDRAWRTD6ze596zQ6Opxa2RMK5OQxSosri
+RfLfapVsTg6h9WYq1wmD/SkTR1DiLcHTNbuxTZpTaD5X1nUkKCd16o19od863nq/2xqQUkWBoYW
S9JUag1TLRBfs76VX/GsNecQKdPEF5pmPSZErUXTAop9kT6eKixI7H/HHUh7v2oDTb77ToWDv2s2
zgfSQartTLNmTD4cFUWRrz7lmzPlzJk4U8K/iLKl8SBu/mrtquoCNv0ogGEbEEHG16/dDih/weSS
Lhx3KIgE8rJX/QtI7nFFek0ybCGxL61SJG/qKCQlgQMjMfm/n4xJ4QF/eCDBXPO5yHxgWx4s4UkF
oyL+P4L2yjC8W9/xqPXVmJVdoIlv8ZJ0N7JSswXwFIr1UYnor/X9VQgSiQ7erjUFHBrhFwGV933f
eZiB5yo/aWJxqvBQ8R6COuIR4QVEbMpkjSyYjVwXAGD+0uNeT4Swkm0BN+NDyg72rafuvkzHts22
BSZbCYWn0suCo96XArWZWRnq6WmMtzO9m6Fv7A2iNLJ8mM/ShKsWfMSE89ZZK+emQfL7SZf3I1Rb
ITo94sYIXCCpELrZLVtqZutHuGpU2UUqJWpWFpWHSUXGejuZ/MiSMIWH4GPAdpbAwxudkjLLLMo1
MJGhY7n2xc8d0s1dn5bS1aSSlD2+7vjPJtrmbFmb8IxXOpKd2fTOiLoJcBQ6Y5WvsfAq7aP+uN5W
qC0akMM4TdB3gu4/RFD2Zgi9bwRrHi2l0ZQ1qrKnVbzYsocTUbIqns1J5K433qDeq4cBsBiFMONb
EuGPD2oNpGKAe1Q+NzuBrNmqBOGewWHSJra5YdsGC2wVDIooijd6rmwvi6y4fqUeqwxht/t+3gGT
0/ux0w2hCsVT+Pm9UniAKFcIc12ATO1P967l1Mtek8Xot1bVlm2O7uuvgzYxVaGfVEtBoPCiDGNH
goaHIC8j7xu/17yBuJjZoNaxLeNXqj45Mqqm7CiF/Sd32Yvw1FaykEoceHmuzfrlZ9eC5cZaGjAc
gvniUSruV4x6qfqK7jnWnMfYvSazaV7lqxO/+1qI7eeb4cv785312DMy/hLYOOWjIwC8owuZlkJ+
Yi89sNDG4cESLLfuOgCwifILRuRJaT8njOtXCqcnpIayM5bSHebCsTjT9jMKazFgNs2C0CcM3wBF
l9c3TjVvRCHnRhYGr1oLVl+lQKK+cC832sXqqxnResDXOSjvk75E0QQfdGWCf+6s+aJyyDFu6+kB
mLUN15tKjI/L6lyHWSSiBu49kFOb5IvgzxkCaJSK4pywpASBBVdolNe06tVZvEQJD8DbcnU6HpG8
dmV8EtofNwElhBfJrM8XaoRyAOOZ4BQ/EPiDPWRas1kOkoFe+LNctuIXo58321UnBZUq6Vgs5li4
rgQaHEmOxfWp54lwB3hjmWmB9ht5XXlwoOeX4R4VXSFv8lZABPb9/6ZDa59+m37rXtRpKsPojvvV
ha+Tu2ypq9m1AQClR16FWNesHmhTt83iZV7284S7dUnIGyxoBiTrg24HxDKLWadvfXt0/eJfUyFw
pe8HW33Cs8XTie2j9J7iUTUT/z/htM39U+QrE45Hlf688ip8ZufiA+TieVrmJbum7ZB9R5Bvy0zW
ulUMKyYMafDUo3UbySIfUdVtpv8obxZT4Ch4b72tQkkWyY4smwhtvoQDsa0qfAcyMY0H1CGKGzPD
77ij9joGnHuDWCw/6j1jm+jTpOgSajKB1bzztJZv/Xpu9uEjV3aTK/9235ux14jat2emJp9186ZS
53jWHRpIRvnmLfv6aL5I4kv+quPbLzwg848w6f/OwHYVa2fX3Aj1dpYAxPeVeEMF8TaH6Jd9A+gw
ouJppZ8ruQiJ4J5VY1+Zh+xxQ4RUkWKt50tLIz7ZLON/KXlOGK6OevfUUkZEICSU0Kw5NjnbrjDd
oOYRBxA9iy24EVNHRK+10YDHHTO+y0txXo5gSv1ZXNxRbR58CnxipAVX3e2wwKD3qglDBfc1hSz2
QKXXb26YBsCgjGzeGeiERA3ojNEefFyKMgYkLjhKng5LFU+0iUBYwwQ20UjfAJ2xjq7rsr3WMyuB
pOTpWagnrwp+ViSGzRU6M4CfZRkzUgIld5AIETAXAcbO1TyQG+pL7Tj2CUCBLT52iF8CqHtDRi6D
Zc93bDA/mgyQUEqpynmZBEjFbhTOUaG0b1duhv/SIzuE4NegrCMhNfMAPDKdBmPmZBxDVBnJZ+9A
YsbK7EgbLZBYobDuBTGJivGEBiD4T5X9t3kOxQv+Kul04UR1qUPcSNKTkxEaFOlFAJUaYvWHzmxj
cZaNINqZwSiuqguzBXxqw5xUSqtmBq5GkTguy9LdNbwlxV2TAKHsKfmjZ4BDxslumZs0mg0miCBY
ZlrpWJXqOhqO0wfxIVcads1f7El/+B+UjL4h2c2CZL4qNOb3aamOPn6jM5aCNgvKuRNwUpSdEZXO
hVWiUc8ebP3fWzf/6OU6mgNpKqUA4nfx8j3KlLvEZH0hnFDd2nSPS+tDfcZ2gO3Rl9in28StE7Qh
wthcK2d3cA2Pmweqwnt/GipxVXggwz4IZIkji3z6QClZk+aoMrRtQKX3QNvQ8eQaTn8gvTwN/Xma
gHMt58QimnB33iBtchfrRsvV4MONkW/dXw3HNXGavan8vsAO+YJ4jwwIQTJKymOHvFSONPWTXrUb
xtbGJomYpJQS9K0OheDzPMoPUfw65jHld1ya6AiLY08VOscNyZTf7E0YYIiLuHmyOe/XcOkkclzJ
8QAmWLQnvdmSPNTIPKbtNaKSntaMII7f199FsOsLmJZCUxHoWGBb5B16Sj9VFpugGoeYcz8X2qWJ
bIZMD7fvP9FTRp05x+JVsJUk6zgI77kCyXGbki8Fprjnzy9eae+BQEIHt18wLGayfDN5lrxSx1Ri
p5q9y41tT+v8U+ATuwwnvi40k+RbaPfFDrIGbLglm1euyFc3kxKrbY2Yv1RgZ6l2GDbwTzhNVh41
+tWRzg+ZBxgxhrtJlG+U6XLz4FHgCtAHOfCUluPxF+v3AQnz389g8FzMsszu8QeT5Siitm/lE2PK
lETI4xdT/MGvefoMxrlG24z9nKMwZtTmAFwuda/wvztutV5qDXECqWzMWB93AEmoar+t458woIY4
h9gZzZ41PJ+W106twvkGIemba50J11ho0g7JDK4Llqn0eaxegA7hTLVUki4hn9bCh1ve+mT6vKcQ
6wSa6bDqDzQ8P3/y8VEJlSTrfeRXzL7b+AbLr60ignlDqBR6VsMVYMc7f4dMpS4FTLD1Xe3vXCEx
6rLiNR6QWXqkPi/ymlxAZwqL5kNI7l5yaMLkDXjDqOans04QDOms6rYN4WrhK0de9dpD3LDp8Q3L
8/s1YZam2PJlB55na5DCwGFBETThIuV/Rsj2OlvADinp8hwGALY1TWWLZeID7TYC8JokGoLnsudV
aA6lx/2eJQgOWacLRaPo5JpeWBsFjgoUoRuYaClvDc8p8NJXQ3gn6l7nS+uAMKahhddJcNxPy+WY
io5dA0XGro+IH8hg8tVyiKM2sOKoWcdigV/enTLpKmLIw7a4J0M6ulsK6Ym0yZb8wU2AykEJbJPg
C/k8LcJmc5Q7uw6zJam75sPH3Oj85FVyi/+TP3sDv73lhtm1OhErUUNAVCDvQP8IJZQsGsfj8OhJ
046gsr3aC5tX7jl2udT7Cw0bGTWWXwSWbbsHckJ6Wdu/G5D4jTd8YQHuxte8NAehvMj8rmmxFHjf
B4BBUhSvt9MVi7p9760pGOzcG4X42akd6PSSoIqA8Bw2fENW00A3CJr5TrcLxWAVoFNKkam1D2qZ
8kV+O/fyX0O5r/MUHqxst7tgpSAtIFzAw4i2/WQ6rUPA3qmxH+vCldlLOgxB+2pqjEBkw8aacx9h
6fYHYh97A3LjvIrflzlNOlzNY2dsIYLiTMQ8v4dwV+/2gO81JUt8GTyJVMpWgM4xRXHhzQQK+ydJ
MwOZkMsHcOGdLxU8TuY6ioRaCoX3uU3z7/40oj/oDwznYXN5S14opjv+bgNDNhAN02d5CZSkP6sy
Y1Eit67qhfvVGpxQaLZ7rYFu8elwWL4ZLDbQCwrZ5++MeyzK2vgYcHsXQNUxOzQQAkXnxxEO1GHf
tb0JDJc8nSBWtPRNTsZqJXo4Q0iC0lsfRY95SDxRHZpggeWrRFiqBUpGsVRjDBOO8BHvyxp4Bxp+
f7GtENZkbaMwps5Cpna2gB6KBje9U6uLJ0+D0msWBnaayhEXVx6eOuqbYZpZq6BzODsUOp+nqvxa
0dBe4+pHNTqFmXl9zm3DcO2wBkWEOKZIO0OUx+shVXWTbyoUg0JmcROlvi43Ny0SSk2DU4Mm4Rtm
ImcQAl6JgNWkzbBx8kf+MRWoIHby+WRH7XrGqBmGnRJlwJRktbb0hS1LwyHM65jnW2CZJXPs0Fzi
HjXGo1wuz50aUeHHHuPc0Nv4/RkcBKqW6WTzbthsSYj1reEpJQ5OlYbJ029NFnLETi/SKo57waZm
B/9vusIaU89Y/b3ODxPLF76bQUN0SH/Vgxwiw52/aBpm/IvHXcDibIRo8lrurgsuuP7lCWk+6Mq2
wISp69L74dJIde61CQckjL9MlIU3/KmvmPwym54NUscf9rNIsBnP+cTFgqDWMr71kyaKljx8a8tq
4XjKPiTbh8hQsTYLMiV/WI8z7V1SdYKZA8Vu5oWzI1pGebJlR0rHJ4Jtg8k3DoSeCV2FlJP3wcHI
S0biWsN0cutIYOIE1wRMVVZ8vEhby+3ydzyUK6rbacUGfPXMF4rhaXqCBPQ0EWBkRzIFGsw2qJNs
Um+V0/LytupILJPDTSe7QtvK7AwwPS0zjLi3Z9Ipv0mRHN7qnRbkqpkTyl9tWCJp1JK/Q2kFeLpj
wY8VADIB1fjtUKnUFonN98au2GclkJ18mMI6jA9n+ogUg6mvqIEvsGkdv2uMcpNW1CL1yDmx8xOu
V+YWmPgZWkFtLTJR5LFnBDjvDVtrEZjhQm0PL0f4/Qgx/aqutOUXPkPxJSvcAB7wx4CrDZOh1KaO
J/xebnC0OUsjH5xZLddm6cL+wJ1M9AUIe9npTDe0+AvUwWmW/8FqQSyjbjUE55iggf+F4VIJq1yW
hfYrkt8JCUsJx8TNncO8oKoTy93JrhiVamQl2FwghSJ4AehnLgjSeq/jbIUKR2CVjl4lx+hmhd5c
DUVBnKi3PE8f844aP6d9EsxvKBVfaB1JWS4ilEsgtbHv9EIlQtis32tdq/sROeyoVDEQB/8laeWs
NrfDhyTM+jikd8/5rh0pbMz5Axj95kIxNkY7yMFOb6N5hcp+bfvS+PYnU5Uk8GaUL36fKoY1KLeF
LHkeCtKAkgyViX/eIFX2a2H774r4zaQOpGv49W9QsVM5I1zETt6R7ZXEqFD3rbcpQ0n+W3pNjxTj
I7yxzOLZGf6fMejVuCktXTMIsuDNaIR5K4glhgOg98TGZZ1cMpOh0uFS2fI4bDF/Xfsmb+9sEvY7
UthbW4i8bm61BM/sdw382EJ7mBrHqSfvZ9kUM34igGgcsxxIFbUfMyUKwldOBNdJwxlALFIeQh9V
B27vxa9tiCbGwqLr3a7+EsBaRtYFiy/pJJF0+TFWMZgPAZfAWvchKncnnK+x8E5+oCClyvtpJBUm
j3piqbd9v2oj0tNIG2+7Yr26pKAL2ZXgz6ELfmU0PWSKJpHiPSVdbYVJtZeLtvmUFNnNruP5gZwn
EvsKPr+CUJxUhigoWuqQhk7Ry/GBWv3wiRVa28zjwtG6zD6kbRpMLkgB0HAJBxA/+VwxvI6oFWe2
svDxEj54ww4hXJUM7YKWItbDH4dMz2/9pnkf908XbIKMw1w3OaYTEBtK6C9VMz+d6vUwHCHqbCyu
pyenMElGN+fMuux8scnBOZcVZXp2bbNsEkbp859uTsnAyz7lm2anUOXwGxT22NIATISye8xRER4h
xlQCW8gH+FmF+JIqgflgypSjbytb1Ua8auZUpp/o2F60X4PK3+RxIGBorsu2PdCpWrVfcDIqAxsn
pgkG4eTP5RE462RQhzAABBFZJrvLHryRBcK0RBoa0MGura6pW/Ee7VTZk99OQgrmbjV8sRsz2O4P
+hL2dVKheLr8VvyqFXJJp5rxclPMddM9XhqdU4IqdKThHqGAaLPyXq/eLa9P0P5JIcVNwSUxZcYm
crb97N7S4Tb2USr7R16GDiQB6+A+DC/qv9yYImkE6AYlpjAY17cNT+ijxW3WlFQ9Ba8+MxOrkx3D
380qLkofIIvC3snWF/r4nfydk05Gj2OB+zf7F6rzvxEGtiKSZ/6Q5UoxmDVq2N9tub5NzRu1I7bR
P1hVS2N99jn/V3GXUa0L/wqRr/z29wwo/GjTaqc0SiupZOFO3aNG2jneFJZZjoxYZ3Ac2drfMDar
VQQcOhUVmCvSxy01oQKqQNvDeegeZaJUUTDq2+Uh3LWFtD+/+WCqeHAnRvkzd8xFqVqPIX4XCB49
3SnSrGT/lK0fp+Axmtenp2VbvAh4Z3yYjmEHVFhj7xnZ4oE1tCZ+6BJDC9o/tnXWXBnwuMRdPlK/
3y8xyqkKagfoApnGrqHPOVt8sfg0VxvoHIO09OEWKgCAJPxnVbYGDZjJELO6EKHyzT1llXM5PLBL
rDvRQj9KzbsVMK5ERXmF4EUDX/w+KLm4138xc821TMG/oKJvSZMGHoKWSIUdb1ebtluIo2OZT8KP
wlOAgy/XBFZvfQCXkGOAmJ6B0rcB8zwbY/8s9i1hUlySY78jH9m686y1eq0Fvq8lbMr490TB2JxM
YQ06Ll6rvjHLTQNi3wpkAcE7HMhUjnOz1IgzlMO8O6TCMCyxaP0p97mjqQ/f+/syS5ubBw8DCv4f
zzMxnPFea9sOr+i3qbxWxp0bBzQTtWc7RzmzfT5lZRFHZBYUBDs/OgYKosQ56ViAX9uQdMuN/KZ1
5FdYsJ5b1FdR6+mVP46Mbtm8R8ME+Y/6ZY2OEJX4T+BDxWJ3AVjVeiU1YHr8FuSajnaEy7VIxdxK
m3SRyxk/NW7WW1pRkt1XdA8yBXrHte8zg1U9elzosufG2RcvWPKZMmaaSP63OdqmdNCaC7+qKsRv
v5UBwNagoVcGvXuko4c8Hs+yTg5NbsW0OOkb3oe4IP6G+fMhZOXzGWPr1s91UvDInqqLPLQwZ4am
nIvPyo7gJgACTW0xRphOsuVWo1ZA+HzHByG5rOP/m2E+fTIfSJICPCBqcUVNjwIEE6qcAho0/Rxe
0YfCtgTR/sR/jT9kATbJiHM5KPSkaoU/q8HmfFwft9KXkUypNNCXN5uKlRIGBnSpo7W0VYrq3K1Y
tbgTrQnOnC8W+BhydyoIOFfmQzQArzYNlaLxdP6IyXthzis1DihBHbsvruw4utZwih5Bx8uEVHhA
kQ+IwFKJIaZ2MJ5hvlZ/b7YTz9QlPY0wR1wJBOg6u3oki4qbr+MGQZp7hIaV0FIZWiK1baMJ0HB4
WsNtiYHgojMvspj7RM9wUxS0Ji+yu9fh3ZZ5u7qW+vZRR7OrMN7AfJi8SgGr9fkTolDC3xDrIs3G
/eps0+md6OWJixrOtsGogyk65ES+dzWKJ7utkXBgcqHPWq1kDQXFV8VOukH8JbT8jqQ8s7PxSLDM
7/9RE8YseLtmEzx28opsKVGmROFxVx81BTRGMP7mpkjC/vLMxgx95qvMS/57rB1T7bQ3/UI2gf3+
JlkGmwqhHGRb0gdxEMWk/0UHri6fDbk033N6XrLJ8rmprOHx9oIPNLuXL5Fw4hBR9xJm6c1E5CtV
LMCHNLxAdoIbyZa+FejOA+WF6hHYk2dgOscZzoUY1+ld1flnj867fwx3UXfCoPKKCorkKr5h/lsY
xh9y4JIjzu7n+UGyoL+9AzySLckqVfPt1MrbtbojaxMj0DFdV9hPNHwmsfNH6I72AAmi82RJ1+wA
YHxhZK34lfzqYu9p/faqeeVGIPAC82n1nDTm/m9fimNtB2eZ1IJWoQiknDm4Z37Qub/eY5iBZ1M2
F6yDjTWobEWw/HP38vlYRqVJEN5+lV9LWwWpm0wh38KI3x4FcsMbU1/cJcSAYdd5QepTss2HEQSb
1Ac9ANtSxnSCsX+jSCvAPEZWoFr2hryI4iWBkbRCNVn4KkSaZKj1Ar0ILZYp35PGnCFJV2yr8AO2
h98nq7mw6hLnXmsWdtSChLZPb30j5HroZJYd/qqSYdURTGLDocStztX+U5k7rSz024FaIaVUSiSU
bsyJM365+6PXLs0UjBvkRnsKjNSfVQry1BO24vynV0/wuS6O3jJQMtj16//k4XOjNRL0C7CPWg9d
eosWLjeDpXJiq+W1SLnf1H6gt6aE4Qu5/vgyeYf2wDywlCJeHmJRjNj4Vo5+FG3xIWfKrmAAWuhy
VOhmkPwSF1As4Y4vJArz7zzmm46DMZfV+ip444QwBvTSQyXoRjPj9Gl7VOSMxFLB6uD+XwjGX8Ly
6ceOcjRXbhPpT5pitBkaUkUIXDbUDDPTGk7BmMuMHVo2B65Qyvfwc6Pz5fbHUT1wK1cvNnXDmGVR
Cxi5G3YRhPNiyV8xf/B0EjVPUhU8sPycDFMqw1G75HyCqBewLXNWU66HRiIf9a6Kd/b/uyi1KXFc
JKpte0Esx4RrJoF1zi7ktFYEkYWpGfdwnjAjmXEdyO9F9eTNx/lIAGrHONyNhqi6sur95NERTRN7
2pRSEM6ntJNKK8ljHZi3SJUDiCfiPCcANNvjqHRl2QUGwMcPd8LNOFnrKkNFXu5g4jJJeVsnbYkW
VWPTP3mLg2zZV2+Z0GNxo6OSzoN0LXZLKal4kHOMsrbj6sja9EgGwPsB0p9Cyja8ZdIIvxGNS+2M
bLnxf7dO4QeVIArIRNTA0v83U6udmrionIe91l5jIR5wexbQRcVtWL+EEpFifYbeTBuzBRid2nzu
uB/qs5jZB2u2HnPEqrlIpVDP5WaD6GAV5ZAJgDXQ3ftvauBGfCjKWs4AUTg+yYER1Sm0Iwvno0m3
jBa/sqG/GMAReamOVttcfnhow6/eRR3HaTBAHhh6lndO92N95WY6vH18L2ZyPEjlK+f2si025mMP
i4OC58Vr29KRuXz3TvujJ5uno6CxMiCj+fDznoVTA0wKDlob3RpKV1gss4hb3Z+5R75Anu8l+GuJ
P6CP5uFX0KyDBa+WN7nzXbm2Iy3WaqDIQplm0c19yP2iFlL26SULdphULuz9/2VGh2Y21Vi7WBSQ
qIK/7WFFA+apv7D+4WZneN1hOvQ6uYIX14KwXkTnnxuFRpJJjuvQ89O34y1tyOG/aQX/Ens/YzBC
sptxHZtitbJ129K4R1IDX49qgYyQzU/R6D4d99q62eINe5uegtn+AsBPTu1eIk+xMsM0bTsraemr
HvhlgQPXuxxXj0+P/9vTsC3HKUgzGDRU5AqoLyn/LUVUeQYplr7yIIR08PXpnimB+K4P0YweTlXl
woVY9tTOnKxiME3gu4Gr2IR9a/F/wGkIwEK6HVxsSPKZ/AwG0aQbhh15UdKGfgsuKwUY84V5b60n
iP3QijHd/LnGFt1+PJNj8X9oHAK69neKuosOZICWMtw2lGyF1WCJwStsipr2MZhAdrbPKJ0OYkJq
eUPnHKugNOxMImv11NLti9mNSBUW4m0BQbSWFG0v0bHn6J2TtP/JdqRUY1QhXOc77CXDVSUs7f3j
9KACKDIhGzHU6j5w14HYm3KOPKSUme3GvtbbnbdtQNTUEU7JfGR2Gzl4V80nB6sICXUVRFwPnWUu
Rb8TNhhU9esGnzLMiKI1XyMLUKNdt7WxVf71HBqH/syFWvSPlLkRTYDQoy2JlXGAWfNDiixCSA6p
ljYPE3oE3xwjttCxdjZojJ2yJzuJhKPcC8nJLy9Eo6Ml6xtlHJr7zRlfn8nxARa38AXXaqJVgKE/
2m9QaREQc09aRp4m/uP/ZsvqGvoOemz77iKa24TNOObyYS8I/6X4KsF6Akp20gWz1nezVCdYuK3w
1Vcz3g4eTaOhwRURuQizMROb2KPt8Qg5tuocCBW/8Di3Xvw98pMfqemJjsxlZnaH0uYh8oEWOII+
Nl95dzR010uN8NiWdPUt2wgahAAe7O4cra6RBd7qAzG55QQ3rGuAb3E2WM/aQwlk9oO9FAz9tbi4
EKDKrbyNNIUTfyLo6yImsx/ztsgZ67BROVJ29a4fKL0s6bVqPzDbrKG1vP6p7kywms+EQW9r0Y5F
VLQTZScqv6TNEpRQqFA92ZlevDptccG/XI7d7pReIcBdkYaD6FZamHaw4imsMS8oVBFznxxtZ7sE
9EDiSo2qnTaAXICkjvqEUDE0e8RehtZcat9GC7sgNZvzCM7fXbxgP8xBWvRSqgBeYW3kRFaH4cPp
rw9w5cE1IKHeAhi6O6iDoFmuJxsw4s51EwldoVt+2+tdn71tENFIj+cEr1xJrSWgaS3eDgsL0Vvp
IFNI/fbNJxokoG6qiEP6Gb5u1JpCvmWs4SHzt0jNbJ1he9wxIGFPIFcOJG09/zbkfaiRSnXMkKSv
CTa7cXuiRckwTjUvcoQQg4knSXKKzYVsM420q/7sZVtCIAH32PFx6KpPKIKttxSewXVhAfk6C2IQ
OvzBMMkEHymnAiq38Exj+d/PGd9CH/dOiCzzLiEhpxzVeRA5ZJsvb7TL+W9/dT8fxNv04yScyHmo
8wBpp8QIQVQntSYBcvntUyfnVPPSVLfUMmpQHLB4XHtFPpb/E4QgV5M68oKTrsVrQfVDJcID5LaF
KcfcN0Xr2glrhT27HXhaSH63rP23NyxMUnaiY2vj9G6qj/lb3eqdKjUmdOfEJqfWo8hK9Kbm8+jO
Pe0LrPhdm1+XwxF5LtH/+VI5bLlX/3kbFICJRQDRwH/cLfCV5ElcXyG0nZc5q3hrB0kqJEbvcV10
mJlGWmqd8nbxz5fGN0K8bw4HeYUSDW2fVDQPfYlVYb7IFFrIfst7vzScAQdWvf7WnuPEFOFs/gFc
khvnwksv92JPXzuyKkIKf9vgGaW3KoJ0EZXs7uS4FaCsJ+bf/+avJOO5z7nGKgjv3SdT/ueGPkHr
7QnzAECq9P0m17aB0g6hBNVNH1PHqB+QLeC0F1Ezm0125pmKEvxnhEN3KA1+T3vhpkml2abtkcVe
RNiC2DZ7/3EBA7zs6D5djKvggBPU4WiKw9NcKrHPrJ51PFcnmNBlUR3ntQ+AvhIUbWtEypzWIOtW
FhGXgho6y6EIvXtBVVG1GXL8WOFKUZ/6xHuBmtyC05V81YPkG/M2pa62tCojjwngWMXoFKrGevsk
KmTWPyAHhUwF0tjCbKmP+m67Dk9qfGPeAHMbNGXxrBi7T3Obshon9iiwRZF/HI4X8YYJfXgcQb7n
ioI4FDhBLdVTyg+rNT4ocb1AegD5k+NcHHO/wQkbarHlvwcGvL0Uqcb7pmdYa7D+8FqqawRy8wYy
z/eybnWRN6PpGQYFtWXUeKK/8NBBYOpkX4WFK44qBrQVAAg4liQNYytQ1j8a3eubWLASuEps8ZnX
bkgnTQMm6myyxvcrnVdnhCn8zo/Mb00kff9mDlvf2qFU/BXTvJU+kRIPb6UjGKNggx6sPfm6TVdV
M4rT+oekcS14+9V7/+JCGQj7uPf/EbIR+mlbavI/4vsPgT3sVpQxLA2VFXjpZptb5y2dV9hnqX0d
B254ICDctYJt9xUMDwbOAWwiKDy3MBsinVGNoljYo10+TBdn6UFmGGXA77ag+9Fj24mU28aJ78vr
YJBCIs7q3frcLLh0eT/iZjbMfuythPLwHCQ9wQOoSVhpkxhsPi9iQF5QCg5rVX1O7h0wEMhV2JdH
QOEbehLkmfT6csyzZBcm3dTmH9C1a9Ls3dFr2KQg/RwU5jCPIqU/A4XVxaYagYYPvqajC1yfgUlC
d13LAFCl5zDoNcFFpWBDs+ra6r/u1e7bc9NRaHoq+GgOg5X4zxn6CSbb5+883MC9JBu1i4cOsi1/
SJKGRr+e0Ypc+956GwD8WEvex4KBS07H2t1tagbbXMGEC2rsjRQygxECUijnpEDn1XnCrCcYQpYM
l99t4cM7McN4QLMy+TIevGzkWGYklSwYOFy2vtre0oMy8qaaOI3Q0aMnm3B465E4G8WEQwSLWuZS
1lsQCZA7HhCDKqW9V1t6RHV4NU1Uu7aOqwwyWk6Q0rUHzCj4zUieCNgh71Hc7U2SCRm51AOVufKC
GwAwWM5P32kQUpGXjVe/PBZNWqWsvxMIqGk5+FRZxn2xVl18YSAjidvrQBIjgHCXIPQ2zLpAKrRZ
qd48QBVgWY5NYenwkin550eGFXZ+EqLlV9AhHyxs7sC/iLn9PR/SMuGspcl+uUTS0zbvo22rCRqB
uiXHYucqWh8fE6z0Nn3sq/IHZ9h8PwEYbtCCY1EcfkUCq4keUF/x2oVMJd20tLu07qf6pagvyPQE
s8Bmayrp6G9vondPU8UV4V8IZ1r4tnvW3XT0AjY/BDEN/gO9PEF3JttgrjB4Bc7uLHbH1VRPZw91
fayCzYY/WTtSGQXY+3LilKvxRonkKw+Pakt+n6r0ER8aZSz/wNMErjFzNX6d/hIuxY3XTm7K4ofi
CdFETaITWbL20ZxR6lpt9kvtdX8Pb//wNwRpn/kbErmbtczWMV8J6WQ74lfOtIXlpbM/6qPO3Ddb
bNUaNQODDFSGh+yevS1be9qt+skoDvPVSiFxj8QKwI8ENpC2QM9DUJY9l57CtrdFJch5MKa4/OkT
52dGuJPPkPzyEfT1gc2z6paH0R5UNSnuHcuuhYGvgR0vmjXZNZ0nnEM3g3EVRmR9kjUuvHp8kn6L
ovFwRW/8goQT4sI5l0KG53yXBdOmkOIBXXOhczL87UePkvy94w/BJqX7L5DKmynwQpA4h0hJjUqs
zGoIEx4YhzoHiDgM8dYTf4ZwUMYqpKHYIYBX0FYuf7ChRztk7GRgVfIkbHc26WjuAx1z1RDLDAXu
1BoxVtYvGZcScBh8PiVMcsTEgi92H3JpgBmaMp+q8UGpqJZygyEodWGPxQQhX19cuXoAtBpcXTG8
Ysw6aWDPzaaP6048i2jdqy6VYgG+8YpcsiYCZ0Y9//HwL3y9xoKaUMGoJnOBW4Z1d4ZoTco+YJ0P
O9BpbwJX4O3O+e5Mnnm1dBZOfjRfmrAMA88j/8ei++6TtwEKgZTHsBCi74gRjB6HnHOnU1CLMT9Q
G5/db9WMdaF5CLa2ZANSFpJ1v9MkaFbJBMPZEJeDPjkcvrLq97F61IiESTcBgcB1DaY9ilxtNS3B
BnjMM8+5+mEXuwquX4f24dZpIEcj4RMTL1x0NOWI+ie9IFNk67wmM05uaQ0WV/SMHk0ALXUsX3co
VBJgHP/PkMZNwOHW+SXyvYPHbYj0Uk/K6460/O0i1NhGCKBcgPZunFMm8AOljDq+nP4+4BPSeNEV
uQvJPu8p76/nj83XGY20kcuNKA6cNKBv3q1zc/fabSKo/eeRAXk9YoZnBkmIHm+KuNt0ZacjsKTU
AqhkXba+alSJW2aLgSPz3kcGJcV/a4qa2d3AtKrUwcIEViKmjbF8TfQDhguKLlgOGeyuXfTbYqCD
PH6IIJbnveLDsD+DzrEX0RFOBEIJhc3AqiOyBiQvnWKBZsZaow1IxqlLcFfSR21Vgiv75Ugk0a8q
cjXQwSAJxpPsLGMdTv/zhFs8sJkZ9xtjSNWXZdrgMGRGJ/ZoLjWAziLw8PGeDGrysjAp1YU2THAm
rbLn3XZA4Cxnb5yPIoueYbT+pbeoBiS6ELTPxjDCdN4r/+g2h7poZmtvi9MwBTGrBrgbZpcIts1C
84A68tcoEr1fRoxFATxgNkFwQEpL1nhoZX/TIjBeLsZmbxogp9JdVltrd8fkstHGh2XS7TNl3iQm
1AWllNlftjjW9UA7kGc0FPThqafuvVfG1fRPBNKVboWbj869bN8wsQpRhmt4fPGCGEZkrRlA1r3A
s+xmoXlzPE+J1RlOr4/f+Zi+uqU7nOtqxYJX9M9YKKUlcmjBF9Wr3TJEGpYdsgZU7XP/uzy4VgkU
vkh51X6umMEfDisxv3c3FHvanQd9d6NEMReYzZgvPzVfSqTNC92Qu6s9cA+69mLIAa1kF3r0RDkf
wokNtgnnO2YjAMtaGshsE9OJSL6ZYcoTEEBOuFBuk+63GaQ6I6r3+8YhTan4SvSEEbKhs+ITsDue
4eCNjZUwhaQZ5JSD3GSXqpUtxSMlQvOMVTcyiPBCgxzU1dLDVcEjQQ9Hpsi37eYKXkx8EagiredI
tkYIn3rMzmAbd5ba6m+d+iMZEyI1z5Ya63i5QBwu76Xu8wZzNh7f0W+gE+Y3bnGhaOwfh6OkIAKi
XuOfTgYl0dXRbDmluBI2Wy8aZiQlGYtCYcm1uMo7/vPpUq2tE48Yf9oBMub99YF24LbQFtPnYQsr
EXy9A5P/1D1gaesGxKgoX3YHR9IXjL1HSwdtd3NVWBGnwqgmoa+vuuIygMeoEYNyrDdlI/j5QoZu
I+OuI71ezo68Xtz65LaFyvFdBuYoMgwGj0BR4hy6Nwu5Hxmiv1gMYFagp5sOJ6kr1YJKNeiCATjs
S2z2w+Iy+OAz/HrM0hrBq7ycuXr1HkmM3wSkG7WazH97lWLGmxhbPaqqeanN6IMoLmywHzvDRnHw
qr2Lv0ewexh5u9wwCMbHV1kX5pYpUs+7jqy3kQE/OyKiUDzABjuoisFWNTcV8g8vz8ko2em6rCSp
jV2SJNMbZcha0lE8O1GHRC+cJgr4UZ+ZMAsIVF6dFEbmUU/NBuLwtjrcPMHfTLkkbk7Bqdx30jRm
2v5WSUqof8x4dW7EAbQbN+36FxGTjop3M7VzTs9XlKF+OSthwTotOA3kTk1PPR/85v/MUnugl93s
ML5eaDZnwuhMk8xMp+5aOp53Oo2//1TS0C7qGkLi10BSn3kWymsYZU947GIPyeduXFtsF49Vikmt
drFf+ucWdXDUEvbGu7GObFD/AinaVQxfDgdPziQkA7NMuu6GJ+M5cGwTF8wSE7HuheNhj4whxt0W
sd2tpiMs5x7ZdvEO7cKTqrQyScdjaPVabKCrjtMslYeQ1P1rXOJpG8EZGelp38MitKna8tukSZoP
bOigvEgImmOBFTn3Efe7sN7ii5W+gr7pfIdmGdVnrlxSxeEr8P1GyME8m9WPfdymHswTUAftiL9N
YOlaPqAXA635opeGwAdsD0+IY5BB0Fp9xYwSyt/jXaspfbdcU/WyhuAGSof0k0tUOYqpRl5fR/GO
uUyRbaCkjr170BleV8t1l5SB/Fp2LiDxXKsNVHyI4mkDV/3e0mlQZcoGsUt1lxqz+GnFwZWMiJIv
e9+bWmspETVPJCUjUzh9+7PGNTGv8zlml8Jx9N+owbCBXUUsGT9z3+Je0X94rLJPuun43bhaQdBL
JQCGAjyUFf6m5+hpBRHszSC26zV13Xs6Uqde8G4nQmYDIu/RcRWkL938Ru8EvKO3Bd4x91Sqdg4a
YmIAHEBq+7/hRJb229Bu+RKyWwJh+qo68Hkr5mslnYTHLceI7L8KViEnAfk1yFE2A+It5Vp/nM6M
fQoie1moyHDt4eTZfazPHkzfT7AogaXKQTyA44nC7YR22cmF2OIL3hY7UkH/o36dpUp1KxuNTd1O
7mzTtjN8byuwzUjqJioTIK0K8/FeExYjE2AJ9Mag11UPUCZssVhKz8ykcFGWqI85y4eOXx/LJJlS
spdqRJFo2m12N2l+CBgY/iSh/rsYbFDAbVR8qCp5XF74EJwUpLMMSwAr+UzQTdSq2UKFBouY/hm3
SnWay92HASsoMF3vRsME3V4Ruti1wYknjLRF2rsgMOmJXmZiQifOycrqF4iQf2YXH+5wjzEnsPlT
vDBj5xvD1kStcTcD+J8BWQmPEQrTRraPmUnJtt/1yXm1SJNk4rkzD2IwfwX5WtKWnOocQ+QSnWvW
P6xJFHPqYMHwz40faw0ztlV89L7iZLrq6OtvmxnDEwlz4Mk/HSdlyay+4etuKowpN7/QN18QUVG9
KC2yADRfRMMBxd+U0ILFn5z9nqnVuQ3NRoov5hHzmLiJ8eTa3YzNZ1SMbLW+4f4jFKCEfeLxkgbi
Mhnrthav/mtdEjYPj68txVRk/+8qyKJq7MdSBw++f9LPA3yPhkfCeyJiGPUE3d8QiXqWPp2NJyET
9NnQkYcphup/vM3zXWXiCxA8Jp/7VkWvcBsdJUPjhO9jG34sX5UU+zSSZkmKQALSfsBUvgZuXqjp
rltDA0Cxl9SGFO+pRewEgPo0MhAKpcNRelTWGNYcO+m8eVUfzI5PjaZH1TzCQcuVpIZvHKTye2PQ
dI+O85Lk0dlaq9SN7Zn7zME7kNLOaOvDpD80MUsO0UPgyZJyk+C9BhTPtd9HWu8HDm5uJ7mI218k
+Gx5CAnxw8OZ5nhnN9Vpy7LMIimO0p1LJEKgFTxAQSJgN9cZq/kyqbdfygxln+ZHQ9rIMQpY35z1
TwTlDHAtuwiLhr6cGBuV5mi7OWZfTdSAH/v47rhNLANIRwjz+/WTwFypg8fZ4OWtDplVs7JRc+2w
C8rUrvWdJH4xTxeCDgpE0l57xl3TlUT797U6NiB4MwU+GdZ0sQr/B2dY0QIZ02uMM6K2qCDiamUQ
bc4gXg282an2KzXZTGJlxu19ohrGdPWU8k8mkW963wis+hU6PVcHk72luy39yma8sItYZOkk8IAl
DhZDqEnCkRt8Kzgtx7hHOKsa06vJTJJrjkzDMhvuAZYCjWMtbuasoRYWMcJUO4tB69CzpzTfhO2q
RcQ4vS157uEM34x6F+sdsv6t8nSmbG+yZRhQ9mOW28sqGCk4WxyR7ap9lvRgWvU5IkPL+sxZxmpY
xdgOuuW9eyNuLb8ria78CYNF6zZuvJdjs0x1N/tnWnUm6wBEzBX2zwnOUjSBZBdMLAZOQv2WKk2m
7Nsv5SwFjppUAZCIeSSexKfmtgx09/LBeCdGzhIrVnasC6MnHXlCxkxIe3RXkaQesk/DT+BMyP1k
TDkDhtirl9MG+QHalS9U4JJNC7QLqRIcOi+YVzwd7+f56EsUqXcf1fh8kncXSYNLywK/O2VWdTA4
WINxIAKmJB6oGgLGT7KCgMxGFRCOGo8xkxcStuYGp/zI1t2eG+vGR5VxcjuStahrLSoF8eTjG4xy
JOIbtqkV0U1F9vY3xMQhDLJgOM2KZ+EwcAQMgkL37C6n6Rr3xemtpZi+CIWecbjM43R3emVsXfkh
kEwVYr8155iNGttYNI8YNapsHniMk3tcddqNTL/JrzzMEO2UMTr42zacsYCjLA1ELoRYKQRjac69
FJJZLgdRMwu9/zXrla4ENIFJtwuJFVtCBa1xKatc2P60i5rQMap5/ua025Evd8yX3oGDAlkONwhq
KX7jCe3XCcfIX3XonLHqQjE3snl91p6doCP220sp+4RGhzWyHfvfq695Ghgk01Qhs/i3otFbu30H
hrNDC2h9BRUCXA4QWGLVBQ7ZLatYKU+tAZ6IEuetjuoaD1iDzi3RqX4r2MSIHlRc/PGTMN2nyKvp
pdlcnBM4oG+t0cXttCTPFu/9GUe7LbZYVWwLrMUCAEaJJe2xpnLD6Vf63QBEmRuwUYa5K5vql+wP
iFBjcmaES0Z75tWBVgN89BGWknbLtidMsC+cpwo5+HlrIf0RdpQM4phIahMIenl1ihxvcUW6tnN5
k+S248TN1FisN/Z9NSQqZ3zy2LHwgVLA5GJjf1SGBUcDhqu4in/wM8WeGg1np0DuRQV/z+sfwaMA
O+svCIWN9XUAbSeQGYiqXhjvmvfYdRjw+nPtaFl5jjpAEGdJ3lIULF4L3KL8cRbIZB6VAwULiSBj
qZ9LwdzUckACT3WDQXOU0jTDPJ08nCMLY9CQ9fMp99SreZLBWiBb5MPnb1bPJipWxbbV4TZOP1Wr
wzLoYf811XoND5mSnKNSXgAWa/KFg32agXtlRs56877xUTJ2HpQ+3BYaOWhuYtYtMaHlARFMRLs7
QCZ9M440seGuxjJh1b3N83W4As9GeCsDLQify3TWPeGOb83qBlXGRl0O/u9d/Np+oeEsUfwVU5vk
PZMP6sh2g5JvvZ+UeD1u/t62Wai4Qn8oUzEDU6Mb6CO3z8KRZka+oC9PoYKHnwCRertbZuemXMQm
vWsS7V57/vQaanWVY8RIVXJRvPegMSHXnv2f/eBzsMrp6F3/yKU/6su4E+l8WUg8sX+moFUcuHHr
BodjW+Qe1buxLcP779tUFDHEphdSVBMkJ42bhoAhCKnlv+pwg4iLIVNk4B+HkPWd4nphjmwTVgt/
nKK62F9td6oSLTzCAI+70+zF3et+76NCwbpAZEmDZ2+gVT1DtRIjpZhmm8rFozvfTCdiqT5bnbjX
ScSLpR0RAJrZql4kBZGOE/ueceOaNmkOmaRWGmTauz4j1QK4DEVuXEQbpDSqAZxbndPMGS+ycdm7
aLmyqtDO02UKMXHwtB1ieOdRmPnmMYarKKjCxCW11YA3NL+4dGKmqQhH478SfoWCahENSJiFB7Bt
E9tRlDjW0ihe2JIQUK2YoQMj8mlT7zZDQnZKDnbymhmFx2DEuUF2qLbDHII0lA1ZIV6HF2QWI7Xq
LcqsJMYSg8NaLOJT5eiwEujw/Pv0QjYt3evq228R9GwObhgTcSrhyT/VuvI5uRuv3Jbi/FecGj4S
pVXbPKHoaYykbibQ60EuIVz1zkvrdRh0/ijLLaNbF+P+7KgJdLRI68LxD9FskvzagEX86NUJsCQM
RZfKTMcmwCdXEZXbFugnT9wBgowhOfVc+fL4SKLAYXVOXNDRRV/5Lh1R7R8sCn/VKh2BdLnq3cWK
eYomQWRGaOrWF7tY5E8noz3omVD5RvYwclsc1gXHEs11fpvLsvM2eqCEdd/HL7mZr0FG32EG5pBt
Nko8Kq1O3Ywg7DtVFFEUrB5CkdptDb8iQnGFUZZfCK5VB1oSBBc6Fux2LOh5iNRRJE/HuSiUr5uW
2HLpAyoLSu1tehe8tbnx5KidkOeIAjd0kArvo4k7jpzUvQoPPlj6RXpVe84bn9eNlg9ADUqTyOsM
XnkdXB5DZ/DlTj+76l5pwbRtiyXEtT/lGQxfZ/vP0APw0dBfOz3z7dz/Jel7cHatQYTYZeIwN0aZ
EESXDQLoOMweiGiuGunJhEJKFezpuRmGbm9OKQghDi/iaFQefhDaBaiJQ8rvfq6AAoFCSE+gqgUa
t7B/9az6Y/FNMiEOGxPBK2DYj9DbYOaCBNM26q8xDq1hfDn0kutA1qGVlkTiwgSjofvV3HUnrFMo
HAqotntAuG3TRZ1e20G9AhDKaenQpxYYB3hOpfgzdQPPEPGhL5BTPxML4nxpcJJEI3UZOyUY8FD2
GCGNc2Vhvw/iJRZb5dxzhr41N7jfP3Lhyj7BDJ9H6SoHWtvLfJxLREW+eWM4aLmrb/reqo/3WaCs
2f+jiGudNrDZKykrRImi/3VxX8TvcKobVd7uuFFoeOgIeerVv/YHdr+om/1YzvYy5kqP2LwI3y2I
06Y3rqeBWb1lIKPMW+/xt2FlORUOBNrbi52jYY16wAQvAqjzHiUQtd3HMS/CXyKrV47H41idc95d
1RCrR1XrPmRkyefkHzEvzLp2Z4ypQwLlZw5YTRZFdWxLRnJcDNIGYJjdXZXg9JDcjHrD11RaNuWA
9NneCG8rThyp1eLejGBPAZ6DnOohSO7Am2/6nwOJWOM3/IvrmNQQeqIsECKd4+OFsdCkDAfLwB42
rL8t9CiT0oRoztthSPIP2a7zRWU2JR33MK8IssrMMKoh4q8WTuYth0rfSoVcz0+5gIfJduAOSB4y
rzEjWyrLxsCYUlUzajlk083s14UPjPphqIApLx10ZEQNWTOc2gNgW2ZKr8y8Yjc7SSy6LouLf/7S
K+ZGqNtaJF5j5M3Txv0m3mDk/P2hFywtAjojDOgb9Ub2LC9RMhPpvjspxTZiGNyfHaApmJ1I/MFO
h5ZB2quQXC4WP/MaUtSJ/5Bu4JGoDnoOZdFGJ6vYxU88jne7ext1h8ZIrdeo3yRwWpPKFeW7i+CD
jrvPEJFsfKBud0b4RlO4At2RybVdewRwufGX4MW5uJq7ux71VSlgHwQ1QTHwNDpwoLV6SebIYHbV
htDuexCjXqkAEk7i8LHt4yT/eV5wpDaDk0tIzkpejBUrEW3HQWHN6f7ASFD5aUVQSPfbjwx310Jv
CbHxemVtnRjfCJqt3+Z49n0z51VOo5e15kmKZdJRC6fo+DqcMnN8x9EKhK/lCtDVbF3gGtD11IJn
+qIol3RvGZkoLOVsEj0fKdevqHSYn1x1Q/PDbn/oI0VeYHDHX2mbPDcn2Lj3TUg9gNIY+rHyV1Xs
KLoJ3J81bp74ZhtI+cUsrRx+cwDdYdi5IC45vW04YLtSYpkoJIINhfjqa4UInSPOzU/HsmDXQvTa
3rBNLBDePsMOzIwaaQ/aGvINTuWJm/+p4KtbQtRVsNrYrID/oF2cu1JqgBQdLSL1pwVeoTGcs9Gk
yCdsSuJnBG3Yh7QOhMFfH77ApGXfnOZmE/ucY46Xb8jByoRjyXrCYo8uXnePjNXSsbQR3ZD/8pAh
U79v2HRIj3zaoHKYm8+uyYrbuon3EZa1dvqm6Al/hAPEmWe/aaMRawfMnCyj9xz/zDvBSD6y1xbe
YxoQCLOte8eySTiqfkdG3/AiFito+i9IpR3jjd0O2+GfnhJ8ZFz7SQalVDF+B3te9Dcpx2UknLDc
hM+R/8yVCXfOzLiHY571alww7xfRgWfFvCA5l/fKo8SkTgBjbcsPPI1aEuXf0+ZJlImMb9VAlokh
BVDiqdKuafj8xIf59fX5ASt7uasrJjmDZ40vjsjUz6pjAYo/4bECIJQ6/+BJxWj41fGUF71S3F0t
ohjTEQdiGTa9NpG0bYcyPjUp7C1Z9+1hy5PMM/lDR6766xWRu/KLyi8AyPklMM8SqKME3uhsLiBS
l6rviWlpd9PBA+f/xea4IWcvCV1n4YF/fwTcOwid5q7H+8gZQFcgARZ7w6q0IgD4DGIZefg5klqZ
X96kMmvUXmEkUk3r60YS6aYDW6iFHlCMULnYIi8SswW8ngkQlaW8qrnwod8O7y6VCCo2RFI+M0xk
IB+8MCZ1fQthvSE4Tml4QoT41yHD+vjOUMiAi0VUr28SuMa7Pb9DSbBhRv8L6TIMnwWrUrM1z5tw
kkHfLn45jyZadhGqFZ+nX9Cn4m2yZZJl/4AkP9Z8ZTdLjJaTI850GYvSK35/St4CibOYE2lH+fxw
/V+gIy7fDmxyXT86bnArAomShgskoxm1yvYqMWpN+YvMjJMbF3j/XOgBuIkXQwxsHRwFmheUWWfW
T9HAl11ES7YMF9Hu41L2p21cZmWWEbednE4GMsWd/NhVufJinMFwPesZmYeQvEJE52B6aG5UeBkQ
jMhSd1hHwMJw4U0zs4Vp0SohAt0IGa9D+yXFmOAAQdhhTQTe5EJRzShIo6dDI7HMMOOFWN9pNW5h
FbKH9c4l2RsjUxbnxvnRLtN4rY7QBhaSAeg/2z52USIUOD2pss9ZZ5PWww+uwkn/doLkqq85ogQf
AI4OP478/GQPLO/viXoV3NCTjSHW2XMibOQRb0zW+SLKiqItjDC6tWH4MwCSkxfX+xt6W+S8Sq2d
5y+zylFHPNxTqrmoTostm/1ZyhYBtCfns5zyACiFXfi+EFgC8aPM0Y6996hk4lUVCfBwPq/GmAcr
InmhoIrhbzL1aYMLvOMVzd4hRee6G897GsaT1ZJtpsopeMOUOGTgXL5WafEDKhTlfG2nrGev0XTz
6WSXZLTOcL1WAU4ZoRAjZKW9WrZsSNuRVrM8NQTD3RfbmYAfQYL0M/OwUeYBac/ZTHFtzWpIxax3
qkMPv9PaRc491La2leoFVXFcjCWPvHW5i4PSxpf3kizv3QmqC0kDSh3FOgVyLVJj63PxEPmX9vf9
JmA1/ZuNm/MwhZcBwNYj00ehpr8h95D94JDRNCH7qkQ6jP8GR1wtx678r5brLufnO6R7t/oDWcpx
EHIXoeOPWIBJSbhUrNPGzcMHRz7h3ygBk1eO7kdWw60toWAHhevtk/XKegjrgSCQOw7kMbEloDW4
vDitNDRFRZw0d4GtNez0Lket+IdH083Bk1zzVw/DDCzR29wZjRsBzbGdVEXDoiyQ8C740ZDzrub0
TYDcMo1FLQnUmQL0txlenQKlp2ISjUqtrfx7APZVZFzus/yvzE7pHcN2Ao3p+PvbEJLxNWoarQ1b
e8BiDi0dqh9SSntMZ4/p8j3OXFcqPAjrZkzYjMHsup4cgXUFUtXpSKaFMono+u6RJGgssQDhZoxv
5gegMarK3sGb283RDP2+2A2dJHbDoVjqRBFWbeqZ6+vvjtuG0lK7qCeZqakwRm3bVZoKvUxgCJGp
Vvy72Al+fkdR26VGRpoWkCSHY5Gumnsu0YGFA7ICUgX9IsTWqqtIXuqva0qMtwdHV2/DaAdGZ26O
2YRma6cW+mNNCl6iipj5prdzJsFKSBFn4m+z6bJ2pHwXkd9CLLC/KV5qtEB0X3J9JXtduTkKBdB/
0is7XVtyVuKDDN8aFLzthQmsu3OLp8W5+CNF59UouQpxLmfovoYSU0Mo6eBk7vI8CIq7mrsUVVzH
kVrlpmQq7taykDLt9c6FCOUX8i1r4MgUnmJZC3UwQ4q0oBZ5rSuBMjRZpcYA059v/Hza1ZpZg3zH
eqsZZbawrzY8T7e8heSUbhGb8rQxP5Iu/eBiqbSYyxe+RcXz8PU9sm8m16PKbxR2n1bjUEuKQs8s
njZrHAdBzStUq/+eiFafouxktiTUrQI9BCtVKJ04W5ToaNI3MdC94RTEllDAE9ZCWy8C+Y2Ux2kL
sjjXXtTcRWNLCe66SBwcyZwLSFOfLU/2sJloQlrrpBs5/qLQUFu5JMfT7tVCZUIhDNPeCA4ynsGm
NMSEH56fZqLL9x6dSMwKkrxd4syLgDJHdBzfqBA7i8/fG3csEGyfYwPHeTeVKbEZeWwib26YOb3a
+YzhVhaoN0S6Uo2fl9lAa6ggmqy5Xl/O701nz1d+fw3TlyRI7ckivqeQdd/FVhFbFydA723oK/ng
5m3uhjrTccNLuXSoUBqKnO18mH9GAk3O7kX3LVDZw7gOB2GeRLwsZ51J1EPvXoZ7uEOfRWtZEdNL
hPV69pBaHVfl6FUmhZ3yBYM6i7fsoddtNmXyy1cs9kic01ipqM/1BuyuzK+j10dMGEwC2bfpSyQy
wk8JYVVajgw0nxGZqotEPaACBsB+uJh5XeXdi27dhxlnMisUqJPLVd6/MHM4pFbfC1P0BpFybwH8
g6xFK6Gb/jH6K+PU1gJuKi+nCUsZ47cqGb6PQyW3cPCTVkW3GbvVwXk45ELFVCz7KxlGquDuEnn6
DonIgnV6rTXOsvOiqFUP3oghkPQzw7qlubkLw8bBjRcqiRP7wfLjLs/6FQQsOThFYy6nBpj1V+dr
6cFjFcPegWTrn1Z8CaHKuQD7xOsPiVniyAH7OuYJUtH9f7flGhfNY61fHPrOO8zpcE23mFiVHqhC
RhIhfutv3h1NoKKGIfsJn2I6sic7oQL3eh3072l4q+Ws/SNODhGN0mYKMSmgnOXiTcrJOWwtNPFf
J5NdIDwRWQVygunECmv2FU3pU19J1epeC7ziL+RezSK0dryaTaV3CpTzAvtkEIKuPL4KRynLOR9O
ptXBQxeytnOyE0430t0+w+ADgH31cZ61mgQtKZNtrqkLVFMQLkdCCcy1YMtvFdltSeuGz0eNrFRO
4cjZoaBmKwPTfqRXR/nzDDnY+CZDvxJAphWbw/HXjj+ApjOXi/+Z7p7PV3viasHrD9tGMAvpbfrk
jeh3DTEgtIn5WD7Fz0UScZBe25/ZNvZDGqerzz45wb/M5+6/VJbcaap6ROoYgM1xlNG9DXtEbOUM
P7vIwO7tPktf1Fk9nTBaDlV2jqO/m0pxXKFzTd+S2gzixKCNPg+G0qXKqvESDEenYXAhKNZuQi4Z
9QsNyGp0mepI+ZVy2oEYwBoTj4ANUYbs11xHJedGbAHCbGyVaYM0M7zAzQueOFlusC2QUQ3fIQNl
9BMxJRBp+TpJ8ISodZNJ4eiZ+wq50Ll85TvTzivv7QHFkIFuMGbtDf9/3WJdJ9Hv/qgjQRougq4E
NSkwwNXZp0f/lHRzYVRvSGEOIBlHcOn85KO/66WhaAEIlC7e5kYmvgFogOjKyXyY93Ll6LM/d+aB
bFPnvNX3rIgcu35fip44iyz7zIKjszaM6KsYjRvqoX94ZKE+h5SdAUUGaXkvTlPHFdHjPctaXfA5
uKayPPtsT2QkFZd/ywU8SNleufrv7PqGdfWPe2IcT+DMCmHWbSEwFUoVIRWojZLKtLGkJGBobcvt
GMve58UWIS7w2sTUxX5hHrQYv4XTsS1mkqziJ01RwUjvMNnH1OkS1N/Pf/DYbLulM+SdBa5uL/Q+
j7pi3QmhdZBgv65uGN60wc73QoAOgffpDC7VodjmtIWDe8hx2xMMSJrCjW2Ggd3Fr4BVyeEYK61+
KwRUfqoAWkXJu9OfmRDI+ycCZNivGBXK+nOSASIrQ8dE0vRT2TgpH/Rf6RXQhLuZSRnu79PMAd/D
wXo3PlV5+wWUZw+EiXVpM/S71UuaVerrtFfjxk5n1JH1V2Vks6Cbbl+U/bze3zEw9+yYa4cj4SfW
PJI5Dozx7OqbmdgN0Svcs6vXBbSzE6PY8VDfIOOSIsd5Nb0vchCNcWI6HotX+le8vVIMmYLm8Duw
fUBYRe3ait5Xp6G793RPbVBM0ZyJ5leGrJfyWV2I29ltskYPpjBy+3kE9ECZ05soHYbMmSYq6CAI
nZ0qiZiotE8yhp0XLa/+I4pXvjzg4wpI8C81ffvrayxIGtAz71guSx7b0I7cB33LMCi2LQJ9SsGL
tgF2VfyXismNCu+I8ep3QZXb0unVQtkfukua6FCRz9S4keuge7aNP7aRF3YgiwMp3AlrrTQIyebP
zc6/Zpn9cbVvOpkCMHKo9+RgCeS9XpTMTxys+Uoq6nZfbenq0D8gJWkCOjP9OWxxDQePZ9MTDtfR
eEsYEfjgZK+rn0D1EhUaWWkwrVsGU8PQ7cWjglwoYJaFY+w0Nzv05K3MAJBCVLfrxm4Xx1BNS+pm
2FXW+S+9nb59i0Ujyl350fSuahu2WshU6wXqtiY83WHEnByXeRm1roPmyVrDRctwVX7ISaAsIS7s
O8ziNjIcdOE4OAETc7P6FIAxrhZ56RB52kVjfeUfi/HxYqAX74w1NpQNUNmiyLmtMdz58+hxUgLI
I7EIisMbfDo+BvGY+uRmtpEXkB2L+fXG7V4evR4gxNj5K80/mZzZbruJFobnW0W6TXC9DhxPmHG9
OuCAy0joXV9xHvp72qD280lml/TuiR2ulYOYW9hasY9+oTy3QbDFaF+6gZQp3umboQgMUdMAdY4w
XiKqXXK8emPevFYBPQKz8IyCxEs0MAUV/O9eZ5QFNLdH1QorjCPjvwBzHpcgMgrot8FhNKcbUl9A
NgflgKC0ngOsFPM7Aea9d1ulaubpuoOtRksis8mqXL6xJBALNvUEukg5HHlK4Q68f/N2JsXEM2/f
QnXdOE9KMamuWNf47wQjLFQ18EGjsfK+LulXISsk8uWhDpNrNAXkoPUcQaOMYs3sw+gotV9yfTfg
d4QmJDve0htcd8DFqcozsqKbcBq0OLcg3ylcD+VD+y0oOwoPSmsJ8WYfnm+W4i9rhF3dfvS1c9YU
9Up8ptHN+X/CMQfTNRF7NTvuF0j9gzblGg8cwcAdEopvQjbx9q09EDIt9uyUSNLTptx9p3ejqgpd
JR8LnK+Krr4qlswYaCRvjSVKYyrcyMVhnIXhO2N/GxU1gaoW01GxJ39ni3S4XVoA+4z1SlcEa9FR
ks2mB5quNfqob5K2HD+XDLKYkzbMC25/xiTsNuAiq7wJglZocjL5Oo+BIfia0kTBqkW8CNU2MEC/
M3KpxtkXV0M9mAFXnq/5IewPwNq6mf0RNUpQVgkJaswuEpfdSpHpXWqjMpBeiMXXiVAuN0PTT1+P
xNjJKZCaBpn0Nlk0/i7LMGJLeqwB0BZ8S4Lq6H5KbqWx/3kacNsprMmOf+twSq26y7uQsaqqA/pI
mUXOG6VcPoUaHw6iPEQRTybkbyH/Uu+NcFiC+OJwpB+Xuu9qtPCnKI3ObAuMZ/BFLfhBg3d0AQ1O
joicrEAwYbUDStm4C0iE7j/o4srNW2FiSHJ+UF26CE+SszzsY03MrHym5+KEYrYxp/RQ9t/tWkPq
hqBElze0+CnGeXL+e5y9p08BmgC4A6pl1oKFNS5cLjJ8DsHUaPTtp8tmFRdL/IjgXbr/RfgbwbuR
dBfxMPL7vRHWQfPW1bmrlaoE6oxZd2PAoI/aJS3Td4q4DN9WAa95ErzMFB7JC6r9TLKiuBt7txxK
GeXM37SyrDWphCSqMUNo1awwqpJa4kXM0P6+aFCVTLkNB65IJbffuefHDZpXoH3GunO15YqtkiFs
2Rm9wePYGrsb2CgpqU2nIPgzAgaE2wpIF05WL+aaIYU8HuCgUee8d7tjW4YGVd7Mv6mEJLUGwyJH
VALuF7edQqY2T705RwwFWewfJXaZo5I16u9pTVHdAKiHu6XcBOHYcLyIHsScxMSvTBsyP930WFLO
wZO6TNHUtZvgW9JdeGMvQqRo4UMqlVNctrAYFA+w1bYA6lCdcgGVnG9lrhY2uog6Qc2TrsN7dg1I
uozbrC5brZetBJOJZpOz8YC8syjz/KPMAvmu3U3eImxCKX3/eX6fg9jkX9z2JxiAxug40C6sRtJg
vR8FUqSD7VkWO+yA+Awroo/Zo/Et4JzedTPeD+A4NH14Tx0UB7N8wNwKrokOAWmwI3kOLyCoBdZe
gc5ijmbdjruNMhZ4N7+PXGulzOaaGLwPKtsa1tWJ67rlLM//I3GhvCTCRWjmX5UsDS3kyiowBwjE
24mZ1jDNHhiEEqU1sNE670f15Zga4/T1Puysf5x8KeU3cJG/nxLkMGi5MegZLParQJoLLLmpiMsR
QxkbsMhBjPItYblvofzYVYaaCiT6Ij+X+XsE1ll29fe3fbQQPysxD9AouOPdLEn1spqcRGe35E9A
xQQrFa6O2xxX1PddDGjPKiSKSGJISzNlFDYN6YoM2qMYedt8JHH8R/4ZSqQa5o6JrvdsMN8gQi3X
JXwybZQ/AaXSxrFyXOSBrFoEpoPIghUMHss9lfO9xAxUAdf7PyjZTVzyFAqg0uKUeRwJ4pmBwrVZ
p8WtWtyHaHFO23g5EeQI83S6yxGy2kcpi073gTe9f8hkk70ZrtyX1GXZAuoq8bKU7cuTNxQECbIg
/bQ36V9trnj945nEsKdkAXM1xvwCDcZgoITL/dtO5uJgPp8EIvoQjTb4nAwRRqZSRFN+C2eoHArL
RTVfuOo4JCDHzbQsZFTtRHlY9DV3PPcWnHO32Vf3HbRrQP+3wEiQKXBm3bko9z/jqTNgvwEkApOv
0VMgcUFx4Eot2JgdnjCKxpni+AjplhD4JbL1DMgmLxe0flfTJEvnp6G/WqEgeuw+ZB3+5BClG4bt
fk7NBe8edDdOZeShDt0n/ogYGgJXHe5gcaGDzfdhMkNV/d/ptjCFtuHgZZXWWL7/1TKRSgzyt6Nl
3Ks94Pw0gzfC8FjNSplmGreVv+AP9QAaFsvP69tf0+8qxXGhMG8heavzXrW7V2KrClSsK7g0sVu7
fT7rwhlbt6hZAMXxK7Tv/9Zq3DI/7wNk+m/j8uTjOuhykaQJ3JRgkbgwvSii6GenLscZzW169J5a
mx0d1lYKb1DKWulQL3j39sSJS6mU0k0BFL2BW9ltevwQavGVaRLzqYjrscnvFlvnJQcwPzI6k01N
dTQeimESm2wiiwzGJNL5SkgdtNUT1OH/nlU0IzbpNpaGu9jnGkZ2ThxiOMRaQbfAvGzh7aqP6Za+
3sIUXLP7IJA0yvIZ+mWUSFn9CG4MDlop3xM5xy0L6GDsFaKSm2MRK57U5fv9JL2ZrTtP2YDcgv5a
JpQMR/otl7BwErYkO26VRAmuUt5ti5C6onJJjXMRX0bGSZBF4BJDJF/DSGKvj9y1NlqA+H48RFDQ
7gg8hD5AoqJWYexbyHNyvbUAi7GRGXIobjbCOfw0ZnYOtL9IAw2Idxxib8IOB2XGfPcy7i4veaat
sM2xXavap/iGNnmPOrVvQxcQjChS9ZzTCZfBSsTLDxlKW7P8H3sTr4Dib8gpiimKvXc+WMtQPfaR
dinfMO/tlsYc00cnjrmZ7eVwtjWwYT8KqokvZ/AIMRAL67Hf++geXepwfLmhO982gaZ4QdTFOkKq
0akwJ6Ck1jQ3oHco97hcKTZmTKLFidJkb0gBDXDCuqPupPcHI4o6eCZI7c2ayIr+NvJ2zgtcFIa9
vlhZE+7C03K129nW+jTQy4j8VtxVa6zEH1sC6Z/BxcLt268/34OYpSVdIXqFKHKmL6aC72CFu1+N
NuLlHsgUz6nENhmvgiEzGNl+PxQ0YjK41vM2kgr/zRRgMnB/55XdIvWU4aNQ7YYiE5P/6KUoZinG
lfU9lsxxTjQqMsz/SnJV3CvwnfZkMuqo9hfhezJcU9x6BFbqNW0XkIbDK6g3R9W9BJUBAsDBpFD1
cIW81zjuKs2JluxXlzSZY4+ULvGOMhrc6V2DgtUz4Mb/GlqtSaiO6l/dkQOhj1TRxKzcbI76Ebi0
aV1KnLVy8mbI1nOvenTqNJO8VfUnnxAh7PP85B+nxh11cIfULNvOgLWl+39UDqDLBK7reNBMXavW
2S+i1RboQvbqkPrkt/45QmnQRUrhlUgIDq/mG3aAIrVU7PZ4fK0w0rtOUaJyq6pREYAeFSt6hg4v
KoAaG0GZ8cglvWIJ00wCbm+16Bne/bFZh403LOzdfowZXL6dID2AAfFQ7V7D1p6wNB/dVWM8isK6
FnVl8dSzLHc02YlfP0lIJ1thosIjHcCcUgZof8fpvwxUp5fJlHupFmQGUxscoFWWcJ4bY+V/9qZR
t+55p6yv/7kT40BGRpYNZkwvGNagnbaxZUVFw/CSNmLEZTDGDfM1qqtv+lP/0X/EtoztgFb2Qt6Z
vrcke51A0XmoM9ehq3SWeBVOtn+78bmj2lrqijBi4NJhZdmahTNvKbOzCa5usfpBoJCsOrEfqEOj
cCL49JiHsxB0PknGkF1E9TjZp0uFKef7yCLhaUjmsMernXDTgsDUwltYm/dviTvCxU/gC3OPT5ur
gra3VUx8RR+1DmP9IjU4JRnSpD9SEqgNEzIq04raqYQZmSdllFf4ICflO+vWC4zL0hLSAr8vpMto
GW3s618RtIezkg7rIPkEBVksyFVpUfnKFG262cIXaw1f9mF1B0caYPFLP4zOkdosF3M5qu1x4YIM
GfIrZdgXm3N/HsYhxAt2Q1cpL9XFhkPeeEXSW1xlZbm3+XA+/DDRxoOq/ARTpk8dp613XZz5OwtV
TDz1ibZU1Qcvl7AeUJHXjs+FZ5UERf82iZBGLJ17ft9ZoMYz5zy1c11vdFh1ITrrZ4xI7K8i6+OP
fiOiiYkqwza16wnskglip+u2JSktudrAilkn6/5fsW1BKztW3Nqu+ZXAHEeeU6/BX1KRiEMg57fH
rASW0yHWO3SPZI0sIgVNmJafOTk2/a22lwzjOBPaHldozrPQ5KABIwNh4jyUHvL4Ede/xp4o49Bk
zEhPbFv70Xo9E4ft0Vedi4XvS9AokydogYUKinPxzSMd2mASqGiP960+RDjdxZEQeFZlsa10oMHS
Kh2wOp1/FhfyPozMlNZNk+Mi/2CFvtwiTstibA0KDwWCGE457FAK3qa+q0iOvJGwmmCqQ5JjAtPm
l6QKjGesESQCq+kBXbGnvdZB0XYjzUBHAgnAQfVbO4J9cFBQG4O+IrzgXRXDXv7qnZA4CEfwrmMf
EciZQ4QwK+VIgSmN6dsWGzmBuLTS7TJAw1uF4HTXCVEntdgOGe+/E3VD5Byi5M/YEXR33Vv7w3Lm
gn/yAZVC69QX7UuBGkSZAV4klft8/VD19H+vUYNXY/LNuAw5s/fLwQf2owgxnZyXR4UEsABVVKM8
QW+77RkkJtYIyEkpZRcpyDAL+nhbtmNNrWPV8F1wytULwf5j6AHp71Ue6rK+NmPvMWyqWtyqvc7u
j6Crjm99nP7MaUIhRQWOd2uW8p40N49zfDiols9+7up0zBRkN5C/JjesEEA/aDh9cNeh38zdQkek
zjnmV07qF9DXT+4eQ/Kfk6PGh9BG1amT6sUaaWh8P+S5TQynTdnsWwAnyyGCU/1velRnh9CwPrvR
1WQ6lEt2ZiH8yGJn0IYThhFrakMqS2ThTksiVbv/BwX9Myjm3HWQ2jLUodfcf11AFC5iky8uvYdl
UxI9xryQrwQZVY3md3gSgFM9LN67SSz+hs7shTiufrHcEYL6c3Hw3Xs1jlpG1Iy7GdYkNdt+eYcl
gD4x9QdtXOECw5C6/luRPwfAN3yrHhwBJhmsIh4kCuumyMsI0rlR92YZB7tj5oYh34xsgXOxQ3g2
ilwXc0DAfaq2W/w5BdlxOFGlvmmaZdblzWge2sTPX46ca3OW+jYwFRbK60YuFo4whRZzM9nesvBQ
Pa4Vsqy/dHo7wdcsj1kQqVRdmEQcZk3h9gWL5Nrtkd6Xh8PgYL11bSJCJYfOwd3A6FC1aCCkrJXV
qC0/i5lslVlKp3iASYU4/nGTYRE0HHQ4EubJ6V5ffPwee/QJ3yTNVfnCbTV+DxsAqbJMq6AVa1JY
6zHFsq3U2Peulb8YNa3zK/ZWmR+MGyzIXdiZhQDyD6PmB1v0F9vM0N3H1j9V96aTv5iihOp4SDS6
AOfki0AiNufOPnV6gzX5Q+HiPjUpN0HiYheIBF8T7Bq3D5blBt1szWRBIpsTQzZBN60rlBMi3SDJ
VKIHGhHQDXGWeXSboSFAYD5fRg+seP6NcLhf6DR3nhDkk93qqf6IjXfnokbC/aVzk+4dM/z4jgZI
rrC6kwT7kPm018KqDDpDCTrnmFee1xyUVunDhJhoV7atAiaFgUGMy2pzaX2WMQJcdPyj7zBP9VU+
XZaMvQ31fGugPxg7HWaFjsdzjngzkGK68l4g35iVnBz1uy8ZffhYsh+Q9mikogU2RAtKftII7qt/
cQHCEJfCjgn/JN2Yx7+fseECp1OH0D50sLbSSRp2PMt/mp4cY1eiM/HSsI6bV2F9H5McbEMHFVt+
2EDzqANzAB1Uoro3JuT85kyOa6snOB2SXFogh41Pe4VUgOHPnE1dA4KLvuhiApG3tsSLripA52Ui
TfDTGVBOYktTvxJ3hVo4FmbmyNTH3sTpQ9tcJr/unoLrzdPyaIhhzO/XVjptP1u461wF+ew1kZY3
mbJXPKljA1HVNb8jcAdnzTeR7NR0Bjdz7BrFvww3SBYgld7M9HinL0Ouc3NnV3I4E8SRQrOHMQLW
UrKGzji9qdo3ft+NczsSRqxeIKua1j3VFThs0WFpcKp+KQy5ex0CnaUufyvmDeWJPljnDPVBA4f0
uiDAaNl65XEQelorVh0gQelS90+06wMaOahmPZDk2bQxUwzqniXfTuMszVDR19GQmA6SOQJ4anis
qZ/VGHu52OIqCvNY9yZfmzPPX8DV2mPg3XpEjD+5AFvf2ZlTpjGpzJBIy8HscF0ShT2+mOD7d727
YCU3UWtDmhp8V8zT+g26a1XW8Ah4NOmZC349J5uCAx+iYN7BG3rVZ4DGd6YCPyzf/dzQACiXTx19
TpwUJV1BPCdeu50tNaliTVLHcqSbLVXJQXEJ3iKvOgODz6sG4DrhljPIKJegvrsQP1FjSf8p0ls4
aK8Xm6I4CU11no7Ac7w1dOiGk1xevq2wcQuqRUczSq1pqR46/adI0KMi5cFZaMFmaWCMhYr46Ztz
KCiXXIjAK9YH3xZ6yKWqOsJlhv0Byx3eAAiTqbG2RLqlHgV14i8n8KOsJCJaOU4AjEZa3IK1GpHc
iKXTlJnuaYn8D1BuMxrNJBGBjjNW4NEhC/32TuEwV6haz8xPb2E4n9CuJq8CsQ6TEddySr2aNryH
/51JBvjVCHqoXntr60/2Z9RB4yX21IaHV+8SsJAt5CNn4Fs4Oy2bRsS/h/rruNQcgJJR4e8u5jDh
Jm+jBNSbI2LEf/VxL0Gz3O626gz+8h+fg0v2bwjBd6ONcKq02hCT5Co4xf6Ctbfiu0aHlf9rN/Z+
VOUDG82rp73yxVZjR5Sy3NHgiyGLJRrvV2mvR6xruX0bsJzVTrPyioMzQASf9hgRfINDfbrUlSCG
LXBqKwyYADqq+yV5GVgIZc/ENRMVnoyzk94ITCMd9UqNCJtBdWQg3i55FpvLkgPmgNmm8WCdoh7K
mXFdTjHWgpPFQFLl1fztmWFIYX17V3RbNcJO2EDhDV0bNWYpWjF8lXLNOW64ag+yxyi+z7imfBHf
wtZPtMeb5RD1sIGZvxCWj8+9Wpa3n0MrTFb6ud2sD4hQSua8GmoAMJ0QhjcLqu6Zk5ZYDaFtLVOC
pj+yorpdtC1PkOg4HcvJ/3hyBjGQcKhRl6R1CvFQxnamKpZQZizE/TeV/bUBhKsDN1ZOvaj+/nRR
dTAIt6zZ0momkHAx8/RqPH4HQH6cmgM+32B34ZRCXpjF3cUKooQdmjUvJ5RXwT7gxBPbOHpIggIT
vIo03toBA+qXsdaInLUGTz8hyzfrcwk1Az0At5vGqQdmSVze3PYjBYBcaxA3vzCO3WFgt/IN5JUj
3YQfhyWB+kUlIGnr3kCbBGtUWim3tfYVBuyh5jj/mGGhp1dhx6ebdE7lpJihUnnBrJG30JgVktri
ZJYSfukhCK27weky/jaqgSTD1RdCB+aWkeGMtzWoHJLfITQI4zgYJfZtJ4uPWwUBAd67fd2C+MUY
O8sQ0d8H3bVGhxYJVFv86TN3wU8v20IRX91WFGDoNRcaHs7QlWDHYU1DSrcSLm4QFw1h6ljyQZEO
TRoAunRDBM5CWvCy7lzTm+eAS5wDGVMuR3Lm2wBUPZV69ekiafJb0tG6JhJzj0X8gZyY89wsm+Wv
zSlaWsEhmIgnNAFE3OueblGUBNw93G7/+TgJgkqwr+vbK6esUaerV+37fCxxSk9SNDW+Jnf0umkZ
m1qTU2mVvR/VcdF39aKowOrjVuEN6uxTpFVMrMVYZvGYYQf/TthmFnH/0uQldaenHakIqCFVFBlQ
KisdCbH2b0HCZH1eQydU6jCpFBOVKRuiM6hzdop7BJGqNX7YsLU/LTUuNVOoQEGY1BTPMEZbbr1Q
UCDluVY7QHQ202lT6sui0c4deuPW5VQCPsUy7Q2BNhbQHU6U6svBLSxJUwKIAmK+5VwYG6XoX7bg
fFLZ0dZC8TI0AgIsBkKz6Oe7xP5lNi+7aaW3uT0XV7SLKDgET8z37LyQNu2UcyWItpzo29BSzvQA
jVUQ0Woti5yzJLR4R4RabAnsnlRIAhqGX90w6i/6F6P1FllobkM8v3dfyg6PNJOT/aDM2aYvX4wB
GuL+MHsYaoC90UYiFrBfmaJFhemKmqeGWIQXCoodZ/Qp/IllyEHaTtO+PLxjFdk7bdTmG41xo35e
e8gWALQWVSOIKlpXr6sngvh86kiwnc3xXeaVWlXT/ICO29AoIIvHmkneQjjgTIu/HM+G9C/Ppcy5
4s17nRVI74KYGbJSa/ZXuatshihZ15Pcctyn3PUEuCY/T4qoOdWenxS7q7m4UNbSN6xe6FE3L4te
hrFXzptgA5T715Ten1pbF+TeSmvLCBKF278bqrvCvSS2eZbuhMpa8Bx8TiqK1KmISJ9aRqeB3s1Q
EVww3KYiKcMF7xGrcsYLXL1BAqVLQDWWpaBpGT61USb4McrS+v47/R56LYphD04tED+87x1sIoYv
h4fNlwbR4Li3CDe2uJtF72BXjqFDuG/t1RuakaZUGBqShiLOs1eOkyjkvUsi96Glfrt0Gpk6eNhI
zHynPeUsbuTgmf/3ZbT7axxjK55ngNP7eWcXBUIbRjOm669/iSIs+FX9+yC33o2Ihd2n0tu9aZ59
bwwbFSdTOd3+NtBACGhv2D4RKi62/iVtMRctJZ2gwW8tHGBD08zTovCrYuyUHwJpPRtAO3IpX60r
HNhwnnGOSAKMtrNdDLXA+mJkQecoZy6nfifkPXYJWTTOG833Z4AVNSrE7P09HdlINj03MT5qRHMY
wbXL0OY6GaJCI+zQMEud8RAswH0717xtZ1ICynOI+DLuedhS3oEmnoj+Bfp5fHEqxYNDiHxor5zF
WflmYAiPcsxlIbXapWHpxikNH4z9HRBXf9tqTt1nbzU0ki71QHuid58lyi4PWgcNDSkPdKRWoVuv
5bCEOoSJNHcRMvD109DaLxh/X+1mxAgeaA1YCZpXuU0HEfshN7aINPWZGh8KuO14gHKkNrEQg9DI
MLDPtaOycGkdv+/Oatl6yVH+a68gs1s138qUJ8P/pDTnqx5oRKBEvHb4onl/8qnfG2QEBopNAxoh
3376jy9+lzzxPf1o1EOs9QyK1qGbbY2wj0Fv3XzZvwEZPigW8B5d68Ltn3o93tU8f4rQgzEwZ/6/
ZR+jlziOp8LX9DzIWJdaIs+56RBe9Vy2AulzXSXI5FZdoJ+sj+Rvx4JKdMrFeSu7Z/4+2vUfjLI4
uV6Rq8UdXEfk02R48OyveRICHIS6uc5pZsjAuypT2n/jKJxZjAF1ycOv1sEGxpZ0ldeE7MQgnrZi
lBdRVQoAHh4znQe+78StNtOi7uiFqIV53o/gr5YeW14XKy2Csvs+zbBDs7IwdVmHdTShng7VGVB4
nxmi6m+42CAAsajgoinA46EVjHfeAusTs1N9S0QuNwYlx/5zPiUimQortXgMvRy//xB7c5rHNq5G
cu4ZTmj3dgrJ0uu2d57ERSVCho78hWq9tTlqOYKrc0C8jtASKMmzdndUI2jKu+3hhVFUm8oJmfxR
G7HGBamkUooozZpJ2O+lzVKVIPnw9TXzrcxyQ8KdLajIUQlbEGHyDhKXyXKsjm59/JWDbaXsalsi
FJ+xZROFSrEIWUw0FWBp6ZmefRm/OBY8eYE5LJZiuoDbtp7BwXhQ2/rAVLfUouTi36fbHa9QV9hU
xb87nw8CuwtAYg5gGiMnHdT/GIXuDtrfveFnksfGb4zrpgjgnnlr6E9QkuG/segUChcQnM4S7D1O
PA5AAilxceyDGcQHToAiBn3ZD4ZH1S5BLD7r/unu22Rp5TDDETHIbMwyhgLNNn9QrYGW9/JH9qRU
380uvx787YaUtovlqbko8y5Xo7Kj35e1rWc1e8P5fIAIn9WTswF8R5F2ngIIWz2UvbRNRytIBfEM
fV29tU5xizIkrHh+4EMe2fpnN0XjaXyNDoDZl0GZR7bqtxu2ocydwVG1TcVJUJ6lqrTxTlJP5WX4
ktwmVHbzG3yvepCGv1Iuax2QmR8YWIxx4Fz9I7Pz1L61Fr+GXOAGLf+3aiMgDivtlmDXGNbsTt1P
ieIhXWfwfaJMVcQ8X0VDHNZBwN1O1AQEi08OuIkP47bHdyIbvvdyWR5jGvLdPtOJaK1BaiuQenmg
P7dSXxPcSaHNn4GSrVp//A+2alfeTrXTEPmJKWK+Ujix5QSZg4RsFTxcOo2BJlRMsy9oXky2Hh5H
WmsTXR2Kxg29fQdVFIux1XDg1JkwFem5A2BpC0IHl1QO4DZJNKUsxPijiFPm6h3rtcxATYXs7ERq
Yj0cSqK7y/WMjWVqiWBX8Te6Qvi3jGDikqmH6AWi58wVtA5tLnGuSvQw0umAEHk4Yss4ga57QUjb
GfeH4wC+n8LgjNb1pmP3SGD8cPJ0HM/iDSRXAsCWK4hob4mALdb8dEN1BBuhDMXf9Ivc4pYprlXb
ssShSHWYBQTCXnUnJqXzJphp9DCTdcXyXi4sjjewKA+L0sDNM10MxgVTUrovC9TmvLLa9wF/5R4W
RkJrquiAMB82pZpwbom966bFRR6Ys9o7Qd0WQ6K2Wb4NkzY0Llmir+dW4fxs5q+UCaFck2HHZrnJ
PnvYj/AEEC3PY4xbLMl9CYRTK2t54h60q0CiEi4pUGVcEoj4bhj84tkEtQawn5zaVhDogu6Ux7+L
nVflt4kDwqE4ih2yBKuuyGlaaO6kt4a6lv9LYZmxAhKXyDVbyo0w9++QP7cwD1+1bQ2Ji/8ghRly
93tEK5DRYKxwRZhdQ9uAe4iGNDMZT2KeHnonyw5Cst7rPphIQcRvwCtQD+coxHhk3DDSU8nViQpt
ROXnjMnsuQ36stQVft8rHAodC6t2O1PwuytjMZ09xTFaIK2+fGYYqxkdFNbX1fq+D/3QpXWp1rJZ
z9eTaJlyg1+ryD0WHcx3uMBNBrKHyUVewLS6Nu0ubfzKFOz7vF6upOc0ujXaKPFgMqozFbZfxAQ7
oc/NQ5PNsrt6y/5S98LwyotbEEeIxCgiL/mlydwTDsbo3MdTODjWSEmFCCLtrUnNqy14HzdsB3ja
yBAW4ncDXPYZpFOuI/wWqehUsk989zLBKVX8oDMt7LrmSnsnkjDb8l5lyW9Wiwpy7HR84sMCVtox
lkekJJSwvr5K60rtspHi1IFfbNsm+uAGtqwYMZadHNNjYMknfx1LMv2udzlrealg8JiEjroaorhy
/21cPYHVFHrkU7jhjHOKXEk/zgnFkvwGexu/KRZaMnAiRPpo3p3m97fflHlJMFm2ixRhSd+8v2fh
CBLj5IUNbiMdnXC1GFZEEbsWy2WYLqugIfeSLMreaWV+o9Cz8/TKUJq7PbSWj2ToA4hDnFJ46XZC
AgkyQu80X5DgCoA1oygJjXmgtx05Qr5C0fKiwpD+WBTl8r6ajstcL4nrz5xkCuz6qzmKQuOl8bXA
IHyPuNR9y09bw+pHLkszRxm6nGdjgIudad4NOGb9Kyf75ie58k2/ZzwVCvdVK82JOAJauMzSKiI4
bE/aFXdEoT1cirBIi59HLLsWjsC0n1MjttKZPrhXj1hK+vdvdPNBR5/q1uS8xpWIkLsKzl/eB6+3
FCmxWlgAJMl6tyIcwv33HNSCGwN7sLi7HRrHjcsPEULkiS+78KKKr+gHlw7L0G70wz+p423UQAIq
qR76YeWyEhU6TFgRkXfmx01iZfG8y17iPM84dqhqVTAR2uJIV8bQNsf9vSfC6WWinN6c/ztyjow/
2ZwG1rFgG2WqJSYJc3LbLGW62Uv8wiZyF/PHzrqtSPCkZVgn37fRq1rbg6pS3CeCPMjllvkhXwNb
7E/23qMpg7gG8YTkFB+boj8BBlW05n7D/FkxDgQ3vxOJG59nfWFsGEk9mztO9E6Of2B5fA6m/VWR
eGFp1TguVUSHLmweEOQW2nun9zIwISAiqFbgrCkkD51TqhZkppf/zwrY9pzCtCkf+5iUlZNIo8bP
ozSCeiKBYyF1aeAjp5SNwk9ovmvU+X52O/PbNAY8YOJygAq+Knnyk2tYvrc3O3mfdE4SJsQaqWK8
Fx5x+uNt689lzmockwvudXbXMO8dONIL5J3Xn4NNcUCTK0gwnLU7BQkOs45PGm8B4C5S0gpFbnma
vwBKXUr+50SEmsPYy80i/ZJJUruIls0cFWGD5bV+a97b6VpHIbvZ/rowrOfdcjHCVCP5XBLkSBEO
tSWYF7I7W4kXq0QcFafV6bHTCOK+eLM/t1HxRzLALRU9BTHtVLF44KlRoknsVGO7QXo7+qmn5/WN
xMshNT7ayLmCYEVFQE0EZxBr3Qh5BXdZZr0clIhiRwVkGK2AIamsHQPuEN3HVk2yzlfEN2r/6EGp
dfxmOYZdeRiVDQnvRMr3SucC15wEHtK8GrArmzHdru0HTsyUNlzfUWh1cNIJVf7q3Rtmv6WvfFm6
El48RdPz2sgKNJTLjZflvKDELley8PfwRC9oWscLNNXx3YSiWQD0AIVJ81soNhv+uepsq0fch/3+
qTKHHmKcYiOFNdx5+Ac6umYhrt2dQH6SPgzSw2kEqTY2OzKlgxVSLzzjO3YOVZV5uf2F337ZcpXz
yeE7CpdqNglMuuqNACYfy3ARVPCafqC4NAQSYb/SfPpg2Tpnc5W/1DB89EoehVHO/pEzfcmnjivJ
pg+Ajy5eDBjMJPMY47QJpGxasQ170x5+lZALheGz++BKDOgrUTrozqiWiCgqsB0yqV2n6m/mTQ6i
KZlC8npVwCl/Fp3yTcWZRSGCPq8JtTwmxDTrP3xn2C4t4K5JFBb4emebgNFxVzA1W7JbIf1hjMXi
zuks2LI11L/jtnlIPnfUCap1jYxCJcL6LJLaKBHZHIEJJJKARdpDarA7kZAYZ13tJgMb5km4lnj5
LOIOMld5D8yqtBgmj132LRoogxUoKRugwUOFjWXVFWmG89OhTofG3F9rXQF0qFth2RWe2JpodZjU
pPcfDNnunokaeoag+zS0f3X3QA9qU/nSdKg0pCzEKYu5/JRPyyxaiNbx3He5x7tqtLDAhUcS8gyM
JNTj9JDF+C68lYJyG574bj8zpq6jYkm84UWULXfeVy88uk36XeEQCHuOGc6Btr7HDtQJ/yXURkmA
M8S1az3j7ruoAYtnTp/cnAGmpDZpOSi4qllqASo8wuIzTlYgZHJHSFXU9C//BQ4JHirxxmC0tMuz
JGuARcSrz2xFHMQ2PnXbgKCHw42lquH60nGvMw3qJYhBZKfD1U9RQ8uB9hVlq9RN/tZiR9rU9m0Z
Dw7p1eSisywTbTmD+wpdBj+s+WwJ6idprT4xPHG0xXfGcDHqOPQfODVxPu+vbj1qGoIgfRqPQrY7
qfPBgVf4c4pAF2F4T1h/V+pCmjTwu0icn0gtmK+lzrjgF3iKUUeL+WTnc9eLbSC8JGJ6Dg6/CPwE
f9NTerWsC37/dW7ToD7pTp1EDp5cYcHNSYCHMV3XKdWEFBc4RbMrm2nt5i4Cu4xTZkacVAZkgCW2
G9Pq+UOPRlqvngeIL70uDG/YQNKrIswY4OEYe4un3G7DuCqX1YmMDMSKA0d2C0YQRPyLmraSt3af
pw/Wwj7YTsROArD1hP1M+e1sirhNsHsHix0WHNN8QQmjOwH69l8UvutlCzmxIaUjCjAjJA7nAKux
Lv5AB0/fYtnEJ/m2pbFUM9Vvlp/TIBEJ0FGIfSEjVN+7yHkK62HQP7TraPEYnfNhzJWeblZ+rdW2
h0fPL/4SkZRxFJPfEEmjI6yLlqiYSWgvzjaHrALkmqqWYjL2908jVKI6ZW10ZfNHpb3tYkIcdRzu
+BUmcr9dCNppFlBD6FlEJoHB3zqap6kMt1DgjtZECsVe6XJ9vXKDFoH8uhx2Z1eb0u4qpV8adVQK
al2Ij05qiD5CXEm2A4T6UPcOqKDNBqyx+j3jQ132G/TbgrEsXowG+n5XBe1BHIpkO0jvE65STi4e
DzjTBSwBjJvyxZIzvxsESDmr3PIu2zeFYIhV2EbFss75mFpugyREYWzM+Tw6ckFgO9eiDTVVXLhJ
eLujhtwE0KJ82ntlO501b5uvUM9OEgJYPeVNhDuiH/reU9ZHpgR6QtDyAH3aAcncvs9wox9hK2py
iiRl06HLuC02skr/cLWvB2KKs3K2BKO6W/kJwUq58zYYku8UbUSgEJLnBt0CGfwfmflIlvRMWRc4
oUd2XOWlDTlV/3f8URI7hjqG839TUyEYQT7EOuUWA91FY2dAyXqs+w3KwBYGjQ5BGDe9kBJ0DrDM
BMJkn6rkFTev590XLfQB5FeE6Lw0EQ16qeN9XSVUicmqe6mey56qeZ9FvAHqYH6N6XVSmUHyjCnI
9LxC0TmSMYfI+EygAcqB3ScPmUz0FAiE4FjHhIVPz6vpFP+jXVZX1Fn5ckwcawj1LsMmNg7dJpbw
KEb3s2cIxaae7mznNdb7P68NnDEEb1bwPmc9XZ5cvOVquaH71UrAO2ych4vcxxftNG94TmMqZbx4
GhI7o02dR2S2f4ep4UdZWMT2E3njNrlBKM9iNyxccV24t79yMrVpDGoMiTInLVCBwhWAK9vt1p7o
O0rcWpNLyoNQ5lLfBc5JPXBk2/qABABziLBp3U5WqI24o+vvocTDfRza8yKuPP3rcSB3pRp/lqGb
nAtXHJM8AvjsqdT+Z1NMeKeIYBdlEIXCzzfT4LAqow5NBNVbH5wT5Uw30sR433AmP/v5C08a1nPh
/tBRyiGCWh6smEUQuxoiCap20fD8YajHdzDMwiRJVIQ1GiupjyocT3tyKYt4L4ZUgWuHI0QBWeJM
f4KKR/me6Nr1jPlHtXHPZcLDRdls3uZBsMWTfwjNG478KmRig4KEuWd3r9kvU7vRbAJ+pPbc9Nhp
nOzmmHlHbMs0xXfyXDChznqg3DcEJbSb6K/XN1irEZe0kWTUFN8wDbTLvB03Pn/SUd97M2i0+LfE
u8jPK81lORyQv05+wTbtJplZWWL4loLkwlfy4wcra3sSxkVU7gFNaI8VL8DyBtX9wkH7jC3Ne1OH
wBIqL9qiXrD/4Yn8WqoZdeCcCVI2nvStW4/t4J2UU8TWc6+/i/cxgd5IemQVcEECodEBpUhn3iq6
TTSy0ALunpWmlL+2hjkXXSGumpdH/AX9VmY0xuCMj1njuZ/3RuS4/iZUCJ8BJ3afHiTApFC6z+1F
nnZjesMdKKEimE58QYfe79XWhA9Sqjt0XP16DSyC3SGEDjXsqzAYLzNom8vEO6Iip/aiY05k9t91
lC6dfosyF5i5NJxWn8fkwQWwznjGTUCd0EzwtgHRaTLKK6Q+10l1DO0AV8yKJqjTUBHmTwwtVCHK
KbE2m2kutO8jSlKRnnLMOBqVggYyhF2uiX5gmtp9mpeTMf2buJwC49sJ36KPdG9vpRWSljxF7Ag/
2e+D5kVOAWpiRlD1Ee5YEOybzknoB3fe0cudVMtjh/9loAbKeEfFpqtTrxAVwVQ5mqBwEYOB0tCK
pHoSFZS7CKBuJk1Kz7ZDVwyWyXkYjgO1Vxt7yuQEPT8LgyXstm0rvQOrXgFiVya74fxyGm7+P/IW
7A1pgwhzuSG7omXzYQBNzNAwt3Rt2M0/Ve6pZEWUoyTdh5WG4N2frwqhmWPXTvR2q8KxUV641A7v
KAubzv5A+aGZJuvpxFX2P43MSsTdBanviWzZN0q1ToRj4wNU6DsTSdTPxJ1jeJh3platiFx9zbtF
AnLH8MIEmuBluEisJxTwmDXiHPDFBksLWNGrji8jf6P5Ar8/41vZdMK/omFQ1irbKXhaiPe9ja74
mwU0HPdRwLdFvN5i1rAWJjHSYGbyfLmtWvbsEUqgQ6QkSvGfAN6EDU+c4aAmbk31tS9noFGA+6gc
1EXT+YVAoRODhAc7qEyurXhXFMWf33qrycGTgkMKEC7ju1VaKlQll/TdPWHXyTeznPLmmDpUouVl
s8uINdz/jmvGOcnLlUaeNkkqyA6EcYtEdU9fx3jV0SbCqzpO0hNLnzHBWOEVfj27qi/loRk8Sdcd
SGhJtqWnLrosWhAq+qkpoB743BcPDtWiNDmBEtDGdtwDjdP6PlJl/RPAOdin5+WlVT8Jxthq/lVf
wRsIAF3rxLu8RmpQaDdumruQEf1DLSXcm76Zo3CbrfGWelfGrg41CUNdQdkln9teAXV+OoRrBF3l
0K03+ZlqFQ+3m9NSHgoRGn5RLy+gMjdevV6xZDYELTUZvkm06VVCZkKpPlo7iHx6e5GZ0qtWmPwk
aXRmVNvA5OMl2rDZQ0v0fhIiYk5da/4A2Ozt7YL8QhXReZidatACyMSN9bVgS4kRg8dHSWGJGrUx
JLp7p99Qqv+YM8z7AvTTVQw887mMXrCBxQICr1fQgbTvJIO/6yEFKwGaNpN+ycC8xYpgA98M6pNM
DIXuTNWigIyWcwP9wiCT0DsxW5ffZf01kkzUGnjopur+tAY0Kbuy61D5Wjo44IwOY75rXo1nJm0M
hKjCb/9q1ZRSHMs0zDFFl4h/HVhMqVVxVPI+18tmkQZ0p6e43lJHFMDnWI9CgrvgL/5qJRL1inNb
M7BfFleNArfOo7yA1j1owz7BLjI+SjzPevHLpF3GfLg4s4CZ5ULvx6ISZsg4J0v/KhAy+GqkNRc6
xbb4EUhpjb30m5TLhzyMybcWbcaIB/ppsbVRcKDr/HbcLEW7ev5dMTk6R5KDZ0vJrLzECL5TwOfU
iG864OhTrp/r+OFCZmsmpUGImhZweHbsPz2ODuFdQEgKQig5kk/gxFBx18c15uaZaBcI7/6h6gFR
gmS7dyZWpwT6EWSf4/penxt8wcuQlFLQLyWEs5qn/tubbq47C7H5mycmfi+WXKQ0YoKKFUM4CEcv
zXyYpoFUJpNtTur17F7iK3IOEn4vfBe0d82bxKz7OhNduS7E2YQI7fDvZn2zzzNuRUcvjVTidokg
x2Bfn5+CORnJpr7+MulhQhMQD7adXMvFsMccarv9IIDIkif8UvOTPzCaFIjZfKLzGimePIivm3kW
pZvPOqNmXDtf9ljIpLQKmYs/T3qbKVr53GLLuf/FQwxz1mBV8hsJJHVOu16H9mvRZ7LszxD6F7bS
CRoVhQ2SXpGqUtb67vI0+PaLlrFdRHepQPuCjmSqXbF0AbCLWIv2afOQYeVKXmByT0Bh25/2DDNn
w5Rr6V94MY7Sadqse+gdneIIOe8vsKAYgSXghtKuFa9ytdmIAZcbygJBPcwooR1QYuMjQ7DJnj3l
M/56OACR2a1PgdubTubJL51YHJLLelvRCujeterp9UOuKBC0xh/hTlBT/rc6CIIxYKfy3EOCMgmc
YhB+FF4JT5hihnOPojtHrQBa0uRHUOVNX0FpXlsu3AiiJs2TCtSIVVQFvffbP2pqkPrrzzjl/HMp
bKtiQkOHXRViU8rdWO0xEq5BFmLWGHNmLixsWxjxjbfkX4rENBnzDljcNcowi44BlD47JVsCeC48
1DsxAn1an0bjiyeQx+Kb9mXV4OfXSSF80yirR4C0mrdYLt8um/2Q2mOC+YyNTc3owdZj0GR5MJ9L
eAatAGU+1j48KYKKKeqkJcDLdWX7QjYH7ALWW2HmPaf+7CoDClk3k4vL1LQKo24iczBUQILXCqCC
U4opGm8XuGuV0VjM6XrnOND3+WcBPwuORbbFLdmznYiu9e5THVX1Bp9ZXPApvfwvV+iuWZcvz2oe
rNJB4Q/Vr2AOEwl0UOnz1BDUYYKGECz5+f7LTP8V27/LqsQOcWFXXvip8rftMx5K6JfL1KW91E4h
7v7VKGzlyI83VXv7QRL2+tVwc1d+pUbqkn2aPRpDragUzQOv82kPwPrYZ+vcWM1XYqn24Oo7Tryw
GOLNSMuJ2qCdZq8mfTYT/3qt3fKvcD9kFRDjyyZSlYIV1UqJLyZvi2ZfZvwNYiQAVf1pCoaVjXMX
lyEAw6Orb7G9UU9BRkFldZ5bwvOy5fu4rjhJtIKG59JjTrYPWE6eDBoVmMB5ub094n7Psa6fDC3Y
Qgbpi+avITOlugFIyr/f0sjTDRkpIfYqf32Y9EB3fDDObVkBd90YhWbXRC/fweu/4JyQ0k0fMRI9
0UGeR4CseQHH9mdW6Pqm+ovs2JiSbKRX/WPm2SYeKoX1dUJ4kcVOcsYRVx9JPzRKQ0lFTDM1OsMB
oGXAVeryCP1EAuS8cJ4SLkwSbImQr4xl4K8QiVHR2hwO8KKryaTma97wX2N5n5oE6m5OfAcVbpLg
sddrBr79PyhWiTTHUQV0MnNrmCCmdf97JViNtLMiuS10omxB0tRfCDEeu4ldPFUegR8rNHOgqi9y
2vXBt+w9qVW/sYzbbxelIj2RhlyK7r/VS38J+wpdHqE5a+NWQuLmgiRYAnQuudiLuDeAVWxCwZmk
pNoCSQlMnEptPXECTvm0DsqEJ981eZgSS2wMad5EOheUjUMfyfdI9/uMKxzz2FAG7hKytc62BN+z
DjUbOdkALd8LW6vhVfVGPgLXLDdmh95RGBBlkocZGb1NoCGQSHbBbebqz9h3/0vEk8prGwIS+CCV
fXr3kCKQGcI/CSrII2Pj8sFr8qpXRjvQ0qQFsNuUkk3egEyIYr788LAQptxPdSX5czyBVcqJ7zVR
jhOuet4TPiW95QqRgrpFlPSQ1a4gvUn+7SUn2oVcpS7x7OClJllAL0pyfxaxE/VI54zhcCEIQigk
FVSk6MgKv7JHeWKv5Er4XX7NCZD71iMnxvau3QckcxtwU1dMRFZadp3iRZvq3bYX/oX8WjCLj3xk
EIaXSSJt9gQ5b5Wco14cUCUfYR8rQscugZi0fwGIjaW2avn+70MgKaz6N1WupKQakQB7L6HPinAI
pS99H//p3HgshQCo6w9+8GaHGhVZmzG4g8zXw4KwU2H2Bhy5eOoGS2g7mBQEWcEjK75xO7BRBhRl
ZiRzjwnMSM+i07N1TIPEUbmV1c7UzOnkn3rgsO++ZO2+ejfdMpl/JtZ4yruit7p73xGW34wh9oyw
yiSPek3ADpYGYtnNDucRG5RMHZlPkGGIvKj94SGG8jEdPordgdOj4NfriautscRDg6QUssYEe3Wv
S6fjVSZBrbwr7x2vNCEyQo4ZqA2swnRNHIAIbiM3SVI5Ii4qCSUS7pmipdAwKy2PjGjLIw/pRqlX
/NltD6xZe55S2MicWXuZKX6NdWkCy7H/hJO+yfcE8BPzkL0IUgcrqn3jLr/OTXp6CGQ++KaPBhrO
4AzLDNg+sZ4OodgiKLjfldhpe3wipWJEwLId+V/UTqECVp4p8AlDn57PH10gZmkBv1tqqfrFrDOF
/qfr4pWn2nE38y/pAgX0u52E122JUtFwUz1qMHtniBwIe7TXO8yVWIjC1ieseOlwuR/b9MNwZFkM
L6Ex1VGpuqwAXr4+oRu+uPrg0/C569S15DsCpM+DN7MUPGQUWO3rrYaUZ7HJxYiXypK26/6DT9m7
ssYWVaH2VFTUHOx548+0m96s5lQRUl9r2SyEli5kmN4KvgRxVxSj+hRFcaArDzMkAMRmTy3tLX9a
cjULgD1IIZiMhSEfavF26RrzsUu1n1kanepmV5uRCZeZaT2YQAJkg/mND0G/SIpVWoUh7s5Muhkj
SUD7FW0cUcHPejAiMTZ+NZItRfGDEAValKsFx5wdd/jpcQewaCNyEmog9OZ/h7OEKhke3xMG/YI6
cGWz+CG014TVC+631GnHpJJCIp4zlpoZW2CXiq7WpZU6Llt7d27e+kAOGzoZ02AKWL+xYXQga66w
FkR3XnxTQ8CF82WBhrRFUWwlq+jaBUJ9Wn1LXtGPCWDuvTiO0L7qRyOEFaIkV20GYTSUJSKoYjFq
FpKIeEqEGFgPFw65DNj7AJbT2u7lkiopBzNKo+nm2fpBrIOSrRuzqH8RLGefL72z3PA+Q1c5EDVq
d+8RCFUpPGeCFbuNwjTUZNutt8HvAWn249dB9akIEywcNsh+/p2q6IFk/hm2G1CmCDfhFduHpUnJ
cJ2NBRjiay/03Jz6qemiA0y0pI4We28OK+/ZWO6/qsgzEQQdaX9eOYCESmPPp5eQuff/YrZSEUAC
b+yqWOh87mF05CSfD80mG7fABCuwXeofrrPHbSx1AQ9YnoX9zYveIbfoH9InuYdcn2NHmhLzxNCr
YZjkEjoCbScjfUaF4N20NEfVuRI2o9lYBZymWsczvBiyDqzEb9MWBs5TDHc2pefbEAl0IQl/z1Qg
V/lf6uB00XEi+/ndDkVbkSidXcNuab7JQYqXWhqdgwhTt2GGLCeY6TrE3kZO9JhAm4E16qMb8Yat
bNag3cr3hU4lIos1NvlUa+4BjBkj3PExfEdMnefsDgcdmbGgvIm9GgfSMP40J55IGR8FXV8cFph1
cPeCbULir75UQcrj8St1QLNkO1nx+Dcb5FfiIrFKfjd9WoNjtVTqD1wYzGGPfzPwoD1hLjyReQw9
VwXdz87dmuPCz1ccoBYAUU9iEI76/3v3APJpGkgKBWLFdpR0UPcEGfVKibYqCaDmePHupTCKmSZw
8ITKXTpCB+G+IgFA5j6GuO5i7byYOKAcmApV/mlnlNp32PcVU2ly9fvM5zWv84ru7sZc+C54w2cu
8z7FYIgI/YkyX2mCbcCW+JDtf/b0yY08iGPZaIzaukW5/OFUBIraG+aVyjGLCJLp6srBZj8tIuYd
Ix0PtsNTBRNT+nTcIQ+ys4UPGdrq+9BhJS38Qmumks2y/51ro9tjc7SqA3sgMvPMCjk45LoatLp1
F9WfYPsuxUJZPDpsjuCC5rjp33Mf157ak/52rh+b6OxbpKf7KMbZxp/8nXSg5zScZmOXCQJ6Y4gN
STvnqL6Yl7Q5+hVmzBDSr/8/8c51mrOaqRLlPzCdV5g/46YT1LIXgqMn0/QfhPGaP59Eo7TEINxj
0TzhZlR7vYQYAX21W4p+itDd6pfn70p/6+rTytdJX2pY0wNtDGPGtuX5MujsCI+1H58zbYczyVI3
P5vlmi9lOQsGBDXboNo+kWaHP9k9ETtKBZ4fV1MrON4OY75gzoYiSJCKfXz/CzZWUdU2Go8/8CXo
advyGaKYndULpVifyei+yZYf2hnS0O2Tq9ZfIT2gy96efnr8WgL0hPNtSFFKw1oRDpD0RrMNXzpH
CVcybDgK0Eadx818rei4wUsVkopRbJAwpBhERQyXvun4KS0JHRRgTUSUkH9e+ml0uCvL+SMPqFvZ
tlVVm25NUU7bnzZhqDvkjZVJeg2HojxZa6fO7PD4ECxWiHsuI8pLrilF7JiVU8IG9Lz5TEXFWGcN
7PLFhQUq+hjdZUXFbutOeWmXvnDWy3U3PeFINWgJju9SqOHrTDh7B7Bwll5yE0D0vylK55wkn1cX
cZUZDliEO0eJt8Ow9zGmrloaEXHaIidUiKv1xs5U0ztc058JKwNkZPs5nM3qtrpq6ca0mvnnYL9a
ulKu8eXz1fK2V7qYP//qNuQ087vUsoFh+wKZXqiw6G5cX4Kp35oCf4pEEncGv84+iu0oXzXmFsc0
BY30HMLrhhDWoMKX6OPTp0TbjmJSDrk89nf9JkqisY58TqqGSJhRgELJ/5Jc9BAlzxWP02y+HFZz
2pjNHA+HmGt5ZIIgpREl0rGThYJp+9xKDVF/nQ/GKk2/3RBqhCtKAaqiheimSPa794jUweI1lP8p
LuEPz8Y8oEGU28MfYrWHZ7Q320ILzzoGdjQVtSkBNO8eGnvauhCdVTehWvOC++Snt4zlT1zYNliA
+On5Ct44cTc6lqsQGuZGTjZsy3LFT8hY+Go51PQRZA1OLr9AYFlcvziLvXPX623k+ewlZ4qWNUhY
QeBTp0UsyiMWNjyomQjT05GY8wrsTr8fARkARorvppLtnCkQe1jq8/xdCUo7iGjWNQjdRHl0yKqO
wLoNcQ1wXz+4qiL2FsUXCskSQVL00c/regNbLlolKGHrjrXzfAg6d0lQMlzenRRSpXl6ll4wOgEh
RuvNQzph2AE9dLmlsGHpcvkV4s80mQOwDG+crijoQmc6k/HwoU5WSJ8Eq6Qwfr0qaGLsPf7fRMEV
7qUYuVwCoSQVpB3nF2invgCp7jp/jE9dqyOMfmX6DZUg3sHPF/qr6uAv6mdhoPBMg2rwdImdKQw6
xScPORyQrS6cH0VuyzbKTGzH4S5i4eMYzXu18FgmQUfZ3P7q1OXdL+Om7S6fgtkGr0Qy3imC3O0A
+d90koEOtpMz0iCjmIe6LP84XQi2kS9uP889woixCowci3c1BeGwISp2T8x+63sZlswDyTJf4g/E
4Ho/8d8dF/PAazWCO48aFYwn5BpMKSQakBItJOxvBrYRjSgCa/Yr30sdUf8TPraQMBIor0shOaOz
u3Y9M9o1VNRdyFAf8RhT3N6tvygzKl53MZkmFlR161ZXiTVDYKPm8371JLTjdlbLWUxB7l+eZAQ5
LEWupJwEiJgvRr7DBZFpmTE8adc1SfMvvIKnNyPC//eJwV+TNx1V+hLI0v5uNjLc1wZCEAu2K9aI
D8MQP6G/7qAXLOgxju4pfmMOYl3r2MlArEQXOFtX5SFo9q/1NO52Uxp3uf2rfhkww+3n6MN3KC8O
UFpjvFKkdREd5U41rZ33plNiEcleLQAajuKJeSBtYTtpapd+ub/gdojfEp4OLDabcr6nlhyl3N67
AclBFgukrzjM2nQl2QZczw22kjYhbuv1uvD20DsFsYR/jkKJWGB1hTWi/2a5Y9TF/xRRXr3dSdY+
ukdKlSNSaXjW4aWeoGN5UVn7yWT5XKC4zS6S78wlM45eyPEinqT1J/gbAErhMpYXaBjd2upFgeQb
eqrVshkIFcEYghqEYdbP10471TjhCUCDFK3NIYkY6RkP3Wf6ivsfRgsCdX7oP7mgUuXNGUHpnYbR
BJTJXgji4AYc63uyX77lV1EJ/Mk2NMDEMP3WSE1tG1cetKyd8NY1o/LPO2RBsEG3qTGqBF1U3yqC
+AYaKM0JFDgVnPU6O5McO4++Zx0TwuKOkKkwKlsfcndtnu93zLmhIR85vU0r2qprAFZNhO8zgWqw
N0fskRXPbw5RRICVgKOer1B7JU8EJ4uFndABoQP0Btzv4BsQZfasIj5/tjHouVMf4pMzj6U23RoR
DQHf6xC7UMZdvZwylfGdNmaomzfUB38cduMpuOXHAahBzFiDYah+Zx0YvvP0sWiRffPlUfBQeiEJ
HlWciyMCEznTE1w2gckcum9AgT74enH98sTMvJKDNQiiMR0JNE8bJUuuuhlYnVVQ8pQS+FXQ42Cx
19AreUz8JdERutg6cfxU9HCc4Utd+WTeg8Gf/tQMTGxSe+bXsRB4qvMMoO29jYX7HrzmkgEqISW3
kUjiexXyFLRZsaKfYJbHF4XS2KpICjcvF2gJua6bCxoRbGc1gYKi7AuJvICIbby9MNG9nmurpOzB
asDmUtHV825FJHesE3D5SuXypywq0AArT9gMrK5Al9hfKh5el9oQSfOMlCJ+W10rAM0Y/VI/XaTx
eckgxL7PjvvhNGUZtode6MIraXo0z+KIX2w7z102Uz5/vEUc1KisdZ+T+nXO/03GXtaAWQV95Tj5
QgmUujx8M/oJWndZlqpc1ojQlZtwYfyNdUr9nR20G1isVtcKuxlC+ukOn6/jqA+QwbAfm+/aN1tB
SjYXtNlIwG7Y2n5a57NWbMGAGiL36bIpyl2Qs72jqV0lL12aSdPA1mMqOgFKjQwFtC+pTHQaDmAW
UIUoSavolXuNKGAAmIcNOng3MhKSpeu/6b9oT0trz/oXp5sS3gFuVE9cqpL14qFXCcDyaKbCYffP
vkJIQsayXseHUGLkjAvU5D2vZZFbzszkNalI0MU41FKnLXKcVaB8WiKud1UIWOidSV4fuiXCqBQU
Aaj3M+Lytc+66ks9imRLkmYbCrK+KPsJQA23UBdVSUP0/8Zuie/x4UbOc/b7wr//t7dsIFhHsWqW
hTNIU3U2oqO726IrM5nGxCSyW0D+EUxilyzhawnYsiDbAH0cyybvFTV1KGk5lzZsHStDpMZgbyZJ
NjJy8H2HaBqNamdYnE/+atmUXb8KK2ZB3QSQji5WU9H+8e1TOojjCyNOeae9K0Q2Z0tr/iuktMi7
sctLMCL+WgZVXCPDcbpVIHrqTHuERW/LqBgh+siuvFSjCYtT7GydJOVhsey07I5gTeB+bv93f1Fv
u/e2r8kpzqVyodbrYl/7fn8ofRC7ROCVBdeSETMCpZx+naxTallT+TGTOmvKrsEKg/pzuJGGfJ6X
YtXl7hdYJ7kLjqj0IecHijmf7RsWl24ZC28kpk4tjtSqmta+yTN/IXH86iVxREVghPow1WI6JP+/
Q1Mjh+FWyRn778duevTl1HQDrsOd4zsz80JicPlsIG3KlAxcDoQ5hu9rmO375EMuLcMpPtwfn/zq
95VKK0VKFzfvoHYR/ctQWyT3WQXfFkoLxIQJTnXO/A25iUt0HZNpBGmdkGaogE+x0WvsLEjMKwPu
biAbLiHZRo1mVOlyUqolnDV46UOpNmfY1hgcOOHBUNckcPyqDb2GWwD0TKUEr9d4nq8781arugp1
8ZKkrLBQCpSPxOgtiia/neF6KFhl/NLF/3xJe5/pa7GIOKmgWI00bKv1AhjrWnhw7h677kWaHoLp
S8tO71CyiLMAx/SQOMtXCPLCoZp9menP13g0KpYNJIDzz0EM6FRpfhrT3qiHXK/ssjQpq44Sfi23
yXY7jeBTSym8MpvQcZZ/5nBVWr1cMvjSOh9gIhgGyTiLmrO67L9n+CEyCT3HJ8AfAgr7Yf97Lnb1
9C5dRub0VvnevA41k1cnUIQJmV1JIsxA/89cuLM3QiPp+Px5J+9wEMp68Jax4h9T0Blybi5YJlRQ
ljQC2b7g3gqpqEVPHY6mOl139P3GJl5lZsvWAUI+WrcbM9Ulpk3fMzQ3v8gJautdPXe9k2Kk44qx
9Jvn7RgPsjbOPT5xhkEWM3eEuLvV6d5GhkoBKJVzr0nkB2S4bx34qOhc/2R+kZNGd4JRr47fc8Ge
wvEVnR8CApEwppJZXN/4S1nM24fvmASER87YVFm0UmEKCvHeVUazt9YHfYxAu1IcNQPIp5MTEIHn
wv3MHnoHpFi0h1a4ZfdBRPX0FrOhGMXeXbBF0ae0QIIE5cE6S0o9AgRfprIwuiXtTJTeDnmn/Gw9
U5DXr0tuZyhm0cXzR61UmE2Vt/1VWQEV02pOMOGBzOXGrUJKpkoxDROwb4gmAlv3HwaR2D06OZjv
MhzArqHMRKnqUopXk0KKaCqrjqfsQTsakvyuiPwP06fIg3iJ5bBjAegnXAaZVhCmscE+oHbS2Aa2
8NEH6kglTQ41hD6mzRzxMpY6daQBwkNdNRT30wPB5eVCeToP1ksb82/2fvmskCe2FLngUNHtk9Mw
mRCrhjrEtd62V86rDn1cWJEF1GQzqq1Mu9R5PWM0TVdH25XmjTIgYhPC4eSXO6i5bvljMadkcpXJ
fM0/snROQMwNeJKSM9FoqBYq9/I4WZCTXyMAMbD1HSVhqhKHJt7+jwnbwYnNGle/AJl7r3pO8hj5
jHYM2IXV+nCim3tp0ZEpLg8wdkGez1LaFFRdye4LQDfREL4NXS3umhW6jksUinSOUm52VlHaMx84
w3cuiEJIXDBHK5f5VN2R5Wh1P1AG6ewY+FEcB1BMZiyQqqOXlZ4u6oSRbMVAmMq7uftQcuMB2B6B
ikO4Uli2Mna1GVU1k9cEGUXQSz1UC7/1nNUXQsxPBCXNyRQbOZPKyw1C/N1Lzn9DE1uqYQGfpZoS
Ha6SwCLn+fulPA8zQpU1UdmvQY08T4PkoZ7KiRSj78+4uvpDwyn+3sp0Nph+JufoUGVXf/UPktGb
p+68WtvfqUkiywe1QqUJjmPLc/HDFgN9F18/KYWfQTCnI/rcwQRQ9f3hcR1/pzLEWGkbUPxG4Tqd
q0lwJIUDqoQ8VO+PjhLRFsnV/xQf6gNy/QnKcLUlQM80vaLhQYzGDLUluSSpgPG9H6yj/ag0ZSsf
6Xg5UUeq2K0LqPb0B8EONxlUIBrsjLdXda3jXwJZ0kz6H5zooF1sZjJmRNl4M8EQ4pt3CpTyRgqG
w+CiPRQ7VIG42ow3ZM4tEeLe8MAc3+1XIIwdv8v+sXo1NVvKUAn+5E5ZAlum/Q5Lpj/JA5Ei6TK5
c+0Fu2sbFzle08vDTV7hMRtMgw8eGM9vfQ/HZ/w/lRA0ymt0d6buvwz6kx5J+RZgOwLC8T5oh68O
ArHnwFU+AOAjGdawZWgODIQEZ+O22zSqOD8pjkkw1nFGmFYTE6rjQlqv1b6oKJP0c7T/HLgSGKRp
k4ecY0tzLmO0OCw3hesIpxaJ9NREtbCntm7Gx/t1EYWQiZpyVu0+7H0eVSGQCW306DSeoNnyUcZp
fhYgJlUAIVisz5FUIZ1uX1ghPuMZOHDrljdt8jCXsbDKv8X/nbSv6T5wtnNjL8fltjjHY6vApQUy
LS3DvNS5HMMOLuMXgg66ZmTjDRJppWCCtbjfRIOggOSZXG7WG8tfrSKQOu4ObKiSgpGEOX77p2tW
DKA319NsVRnmw7O+yr+0Cxtij9ExtSKruaYTCimlBvhiY3bViOdhM17rJaBRMefu6AFe/pYaVjXD
rry+Nzm87VaGnRhHze2dRh0DJyicvoDk3QgkvCa2gXiztv/Bvt6SL/G+E45TRhJ8GfrWr+i/wU+w
Om1uBenIt3Wrxzx87u701IrimpvF7egCJ8y85TnPQc5ZvBX/cQGnDjLWnHvwAJKh8/BUyrH7HJbB
PcNA7DeROk53aP1OM0182fKa2nknEve+CEj1zQtRVvOoC/dK65RLGppndxAVrpFoEV/HtbztU9Wn
/dLNiGYw/Fq67hVTlfBqp946322jseIe8uyxmQKr/PMZjOV6bCMlGolq5pOjRtQ3zuf/xnxaLl+L
dZqQQng4ztb1jprniYBMxvkG+1aBf00BVr3yRKdoH7Jf1vVr+trUKVpFTrvx6c5/S4xxuJ19gQ1z
1ks3J+9AsWgE3DIn1UYCx6qF35Wo/F4n+ecbUidqEXZfphm+p5M9C0oF46GojI86gPAh0qLMEIbN
SU9tZ4v14aBmoSCpZ0vel5WybvfTDyM963/AV9RV19wDrxCemFuUJMHEr/ft53qjjyn25lfw1eJc
B2A1fKzC62QJ/bzCG5C/czswG5jR+46MmIK5N9G7AzqWC1sZ8tYMcyzq+2eAzq8DtPPhqYFV0Ukp
6pjFLSfoj1FZCgu/LkjGsPqF8+/z4j58nBeZ5MeaYTl/I5Q5kntx/7zX3tvjqjgs6RHT/GMS8Hwm
YGKAHIHu2QDIuEc+2Bm54g3/KabEz+yZZ5KhAhzwd0dOCl379RvXASuL1o8Wn86iKBXftcgrVLRx
w6E36geUOqFmCaB0k3IcYrKPycWi+It2oXE+I+/0akZyhLaCKD9mABjC4AhaGhZKPASnuy42jUHl
Ntdt9156LlFQz+vD5yjrYvW980JqumYZvbNgckvJ7NcSVphzo46I24q66x0u3SjPUMTilAK9jwcm
1ZAIkXNnfifHmiXi8HUIqSYr2XLIC63XZ0KsLjh7NkYtDNsSTvjyE3AgjtAVhaoe5Bprw4mClw1Z
Jbw0JlehPw1uljxqjbpMGaGcqzHa3A0eyK5B4r8DVb2Vxo36jNRhh6uEx4wjjtbtCBQ80T+1Qmgo
IXh6VVpsUK1hhujvqzXH1Qn/LxSFJ1N9pFbzmArVa5uR7LrXP9e6sXFrxM3pFrVmhw2kagDSPMcy
pvPKHoToBaHLIcJUHeofdv+NdIoIUt8LEf46g18Krh+0qqI/hTvZVxdyxnUqKSHxXdPf1egdYnqH
klERBUFztMW94lIy0RX+7VIk8cGTj2GjxD4KqnTD4vV9hugBiTp+vMsxB2LjrX9ADoYR2NAJipUE
WZ3SJDR8QFAf+A9wkO5J5m0JF5kLIvKIc3WI+G28mDos8M2Si1GrMC/TbksTWN7pzT7wXtQir9dF
2OBqNH4X0z5MjMtPdj84PmUttF5H+1djzNs810js9fPzap9Wgl7V5dvWPAe+rgY4rWoA1ctEUNcy
5aQ3csBkhMkVgz9hOcb/IocKpGp8QWvaN7Qzyn+6lmv+AbtgvsX7FcnQUcrZ5T8WLbfw3DHNaw6o
Hz4q2z0mpIXSzmMxSW2y70VIsorFLobrLLbagSvKgzaakBYUe5ePLWJT+3veHjv4kEL1bpCakcmK
Db8t10agOs5L5O5P/namvfNSLH0qwLnzLaIdk/hyvBRZ/ElBShpQe+4iM7uOfGFaH8qlKzt3a+C6
myEZw6vdhSF+Qz5uf+hw1gB6eGfpCIIDGebMXiD4ugcDOC8myl+vwD03o37StNmu2QRkHnjQ9y7O
syBC1Qd+nugXYJvwEEWlSkYj3twEMrORB8uMKW6R593j4eNAyHk5JoijiaLfQdQYPiyw+OH8hIcZ
GfkUkaWhn3dCl9fD+Jd6F+nwEnHouMRDyg7H5ASB0QDq5EafHY4BjbBr1yn1GU897t5XnHNfHdq1
XxRsZ7uS08/2Ikf9U83dbGB8tCMzQUeofhL0251XMbIhHYiWfQfHlo5gdYsl+yXUm0BK7j/+lM1x
NqXyNo71LWNHLyHO1jWpff+LVOMDi112XY5grxbZaJSc83CopLDgfOdvUKv1TK5/UPlbK29FgP3i
lSOXHebFntL1+SRnZGkeACe0EzOM1vJSxPBGPBNuedfWApxBPrc1Mfo0x6/uXIPpCJ51zIY0SGx1
sJVmOpswoMyvOwI3fs2kecQPw0JlUcGkTnsZC6bBLeK/A7rBUBlxH4GWIKTlB7xHAM2rchorlUz4
ucu8Y6BqcjH587/+Vs1NpHxx8iy60c7kkOBHMlovYdNwFKTE53llvDAt97zTw1KY54gfHGa127/y
gW6yCmX6yzwikKcbuQUU4CId/Vmr4tC6/3I3K0sqOqzXHw6TaQHxEbgHIszKNtITaR+I8SckyPjR
3yLkVBECE8/I7nm996YNxwiVGucSj0cwYhYrCXb6hOn6khErQqe2IIYG4e1nDAwOzHXlcVOtqjzW
49u0z1SNDIJaIMz+I2T/7AfAIUzQ8eecaDKj0BJWUkiu3LVAIO9YEdPj3FBUXaIBhl+RZEu5egdh
hub6tZy/GDo034BChGLZlj00FYuwgBy2vCnzN6QPHsjnB651V24XkvGRf66pilfYI/AM7coPPMWN
lyv8bf2vDPRAB3gDZhY2eSBcMJ3L0i+hNyCDsf3tvgY5CQL2uQ2Zh85sffNDhvQ2lT/MpMn9xuXv
tqHa+CmZK1KmBDwwiWNNstI5E9kmHSd+frYRZVdfGkPjaOD9dKI3xsbx83BVTSD3eGRzkVKpnjcp
Rsja/+jCsOPVGvt5sVLQ3NKjxAyLuSLS4zMsNRV+gG/LNKt/+f9KudjWcAhUKznascGIp7PxhQdw
rgiZPp1lL0H4eWvKwCXMxl33SJJ2BOqfl5QO9ArCFh6NxlWImh8CfAKKvTCBy4G/Dg7fD6Rm7piN
wy5+yZG2L+MzEWcYkKnhRpjvttgQaRcxEveouIiiVcxINrrjd5RwQJwKh9NSjT3hRCOysfufnSHl
yZ1weH8sFdPXkJUwetVaomxvi3KE5D/+QzfMQtisWqsjor5o+4p7gKxr72OZ45va62KV1oDX5MiO
vKqzugxuYtVQ9qlmatboXYqEKWB32Wz+reoxMk1FXuGDVaE1hWExEpQai4pV9mJG6RyWQ97XODaQ
H7J4Hu2ST2t3vta4h8ZE4wdAdcidkwfjs5XD1qYvswuNi/H7+vQHeKoe0md9Peum3bw9fu8//D3r
uxCVn1fVfUx5rvhoOrCFywg/Lfge8/yLLOrpQnonknlCEimuia9iwkq2mOQm2D/wHSqbl+9kXoOp
DJnCYAsPqfSptsxL0osvKTRYNBDWDPL4nLRqhM/RFC31Qv+JTRYOGN5VgnunhthEaBOSDRODQmrs
SiMMB9C2rnViYXlNIoLehZnbCZjcSgKWv/qZYtckmK1F4jiyVdu6vcJQuBAkGkUQL0SWJKwIIBRF
RnwxbGTfCCJm8FJ5+fLTQlx8f2mJWkbiscCo0/ii5K1rWQnQEy93pIZg0JaBp6csXIJ2TbLX0g1K
BJozG3ESHnO5hVza0khNsVhXnDZmP2DiB61jmzZFl8FZcsLkTu50/5tlOViboWeAh8fFpaSezYl9
TT2qbHw+7gsU6F+xNEl89c8V/T3/NE1OklQ2RNZTReg6ZZecZ9iAQi3GXpBRDq7KL0T4M7rOmUmg
XnzKJY5wmSZtTdmgmhlT7CAAG89kTmEUMfvxHeJVvCTfgUBZccLfv48X4uBAflgRlTK5isZjGXnn
p/VdJLKJx4+kjKnyoMVXHL5WwUsoJ31QTCuieQpbIlNYBYBBnoP9iF8qqeMJ3BFoacIxu2cpiPrw
FCAZ17HHM8evk06m44I8xj4Z5XAHjZntil+eUPor3wxCVfkuuaODFKQ8+bUw+EAN3WpLbnApJqbA
rEQGWEKyoL4Xay8J7E3y+lRcqe0Ev3QuqHxuPnbraNyFpRYtvqobynfRQvEv37kPprq2WCYtDtvI
xC6cIcrkDeRpjNF20Yy//zpjU6r4IUOH2cHPYYlveHlzokQtBGcM/Kw+kPg/jPIJgh3dfoTpeeIX
8C6yQHqdo7aoStb4Fmbj8vqqXXLsNtnTxUE0RWoWFxEi9bCd0KEHLhqkYSGqpa/wWavkpDyrmWeT
19I/jYfyqNCjQqvXjES5tDRW8jkpFG/nQmwxh3MRXPm0hw5uisortd7xhOwh86QCeKuPFd//AJP4
tZ/q4EGJ/ZhxCMBUKu3I2fukaXuZttXiNTxBzXksdegub8/9d1lG0KCz/k9i5Bpwf3uuIDVuHRSc
HG2+FK7E7noVJDFs2mxmXBQF8KRlM5RXAFoW3t+oApyucialoTCDfVTj1WwA7FwlmWrHhM55mLiC
I4TcTHw50iqUz117+SYMGNDVWFVZU4E4RANGnDBgkVb9BA/PBqD0RYKf5RAH4jp0xJTAQe3PxIrL
YKir847jtnxIdMjfmqZJwGp5fwNwGDjGZy0g0HZAtkUYXE7CGxBk6Xqd3W/wd0Rt7CzPVIa0WJ2A
IYQstqGbDu5TVldYTHMEvrjA5dJMe7y6P8obcVQ5sd737Kt9IpOeijQiogD7Sw5GbP3AUSHD8Sef
bC3wm4WSGB0YLyV17syF1i/sUsWVT28ehRMd2tqP8J8VwOKiY+0ojcE79FU2Pq3z5hmYuaBNg+9X
mEVTz6wr/GrNEuW4Ij6VbCrpEoP1bdKRAIvEpPh2BcoYR51LTQJczKBcawArAnfgxgfAb/yPqL+x
Cw4LJFBx5J5s1PwL0gkcet8D7AC0vWYSk+zfLVkvoyABThtp5by+1rqsXRflXjw7XTdhT8/AeYYe
qTfl3M40WTuZptI/9nOkHFeyhtODzEPkU7r8UXEbwpGYpRVxxBoDzgY5g4xy5jKenyke8RBNeym7
dOsOGZX2+MGwUMqUkVrz07r/d+KgBACdtdA65BG/922lkEHAlMJnxaeM60qb85R8okwL6L2UwG1V
ekR4fLZiYhQjtCtu6Jm39T3M5rqa0bg1Fgm5AH09pdC3paW0AjB2EDBD6iuNKuWkX2Ifra5hpIZK
86zR0/xWDbRm8mSV1yki3ha4B7S6KdMDpmB+HiP3keZfyuDXlhEbzHGeiAn5en9TUblzyUSWDRCr
8TmO4+SBYXeYPYpIeAlVNUu+cezcbd27OIncFB3uebbNGLweGgNVkRwsz8+Px1OLc8UcAoeqzX5h
AfZx604vbJd1zZ/+cNP6fE25sQbz+9be/JvxwFcV1fy+C8WGDlBofkWpHGdByA5bWK3bzqhtI2T7
VQ4/Queyrp6hHHsyewPjPNri4KvOR5U9l/gdMuqz4S7ZGkp13PPrSDioi9x5baBW5arZUQiWXfDm
ipshmzMYfHP491HGYB6mbnOlNdWs0OEkfWNqN1Zyd6gK6eatJ6ZKazc7YBdV1+FCIHYuSKWgvqGy
jS+pZE5ZiiXTrYxmj0V354Nsyp1oB9VdOQ+yrO3ctYYov3oF0IoV8ViUoXO0G1m136aMnAWMUL2Y
dkbYAccawW7fSTe2iiKvWiFvPpl/4KwU9BdccUUFy+MquIfLZwfD0Nlwb4WEpse0F/rCAc5Ypjf/
YmXiXRhsmjvp/is6wtXVTVz4VVT4W65ymZfc1X9lJr4mZmJRBz2bIbXV1+ml9YCOxSKgaVeLIVFc
M+GXunLrzdd2mzwqoltFdsUFJVGHLwPhmwcfBD8Zv5IZxz72wo40JrZCC8YZkoQinWwzrVYR0Ou3
64kC9nVxNvSHHYOK9js4InsWPKG6bqdIDNN12WMk3F6k3qFJB1+I8WW+tGVbencFgx2jEq0cLRlp
hqIKazbzJSSRkAJvnwF6kyooBRvLEFd44KHs0Bd/j/m/FMfs8upWVpgtZLryOcrW03ncolKvjQeA
m6+crNDerRjtCsNZ7xbrOxMdNQm73SJh0jqEaEmz0AeEFfDuzvRpWi0PTV1LNM3x/QRLHPv6RlkY
Yan3xwfI6kQu/LbeQdmVEAAZG1qz1cAN/+pkJt6cV/p+gWcsSCejiltBVlpakBK1BX9Vlj3vHmeP
0ckCiK81CyVBIlkC7AVQt55sezMIAfkaXCU4OzlOerbBxjzh+ZEl5xyiyXQXtA2GdXu88+xl7wWh
zOmW/lxrFxmUv/7N9jsSJPt22sHxsA2njASQO/NPWZg0YPa+5dUxqQRxftkWkod7OqfQFHcpvpa6
gvk/WHXVXkz31/Wakrwa2Zb70JXRZrcufz+PIgo7AEHhufus6iZiI91Lz/ZV7h3NqCBNQAUwiBTt
gBOnnxMNY6RLdrNYqipVuf8kgZOviXZ6BveYvEMQHFN5izLSbnJgwIXETMEEEKD5BtF2G5O5s1a7
szzQVaK1DDFLOav35ACZc0CIkQF2VA9w+n+Y9lKvyB3SQRrSGCGqlhPRnEDE35wOO8KSXtem7FaJ
bhC9Gqn9kPgldbLrCuu/A2L52hcFFDixWCcL4sUrxgts2yDnPeh2Hoy9xw0rs905u4F4nYBOXpaq
eVuNTzYS/9hcZwiWBEtuBXlea9lNORGpRLaNctH+GPZQBIHkiJ3Vk3RB8l+d6gRrz9fdFJYorZvH
kVbs2mFUinEVc7RF0LdNidxiBWfd2Rd+Eqv0ANa2fSxX2a3uIDTx+zrUJRHR6DIa+FxVq0CxNuPa
UQiUM/UNRA0j2tDyWpTNRLpvV/nB6e6DSIvCMkRBWhkgqBYUo1FECFeCS3eEdvmsbNf3aa2m41Kc
l7Y1NHRtUSTVGmjRpSBzjWZVZSRlU6sSRf0Il8ECAFzwA4Av+0PvD2RLlLNLksMGA0DhhcYomLhM
SPuO1fvDlOCM8Xu+lRVKHxKovibxZv1c6wzNZOhv5ZJcvDhU9t0F2xU50ojWO0un728IrZ4/3jaQ
x7gOQ8KeeLd/Xd/yz9BaXi+nGj1K9YMXxMkgBAMTiOw7Vl8ElbfMk59LZIeWtgLEvq66XSnbvojU
wkndo/Q9s5oe9JlveVa1ly+BdfZ5b3hNcoTuM3CFI9bMBNjWBmL1avBVgOtH8Xttm0Uci08MjoJQ
Dk7v1hagsZo8jpB+N++Kf5Hi7rr1LgsWEphgAW8RYxq0xKH0GHQbYu8lYQekQ2QE6idFpJR7Wcdc
Ks2vmdS4Kf8AfRenWEccDMVl8EsyxEUvx8T9LVO08TnVFrZNzyySG9w33tj9hPV9qrJsT44CsMtP
bF5nrh5TJFtyLmTWWzz0TyzjVcT/IxQJl/CBxfxXj4RGajKGUQrYbTCkDcT0BAKzB1/zKg1BJuMZ
XNtCVJ9iwKaZiVyhzS8DkBDfe6UJr848fwCl56AQBhEtNGIe9rA/8j+J1oZAj3y2B+n+zwJdRI4p
IztlMhSgKD0+vCOdeH0L3aAvd2I+zx5Dz8PuQyA2qIth7yb53ZRJFCqLZf8cqjLJyhZVCO21jhk5
/V2PG9U//XdfWmRNsezS9Tkp27Z+Pyu4jGKFLaE594Mpi+9T00baik6kbVdq2GbQVTnZgBBJ4hwF
o2KRy6hoge8NBKQERfFh0A3Ehp34cmm/2y78ilc616n27d2qKoMMZY9e9O65b9xw+2dQcTfvK+pP
ILOE7vTR+J4fWmnjO8YmXVhyWOnuFguJz86VQ1U9n+dxYuxGIaGDjcDsbdBVnzAz6Bu1aYF6VcJO
pMqmgzhrbHnshpr0iyL8cdzzRj3fGPJJbGPsDWYYl5TCgrFE0lWr346fZ1Vounxg2aGlrkQd4OvC
4958dbhZn6TIx08Dx1J0L4PbhwOHZuTaALWX+meQ9QZ5bTBCYF18yCWG4Wln1GOXNp6b86SB1qzQ
CyQKfPQ4CC3wSEzuGC3vYFXGbZn97e3aK42VrOQP0LtbdTzDKBfLhfjPFABwvaoHVTVVpLg2Ti2y
0P045KY3nxd1Mefd0w1sZZRqktudVQlwtKI09ARRJc25U77mjnz3bJMslCbuRrtzGyoxOZTSKzYU
fWUc9kTqZnqv1ZZIi2h86zvaw1lObg7I5Ho3cKl9HRwp5dVRu+5QLuc7/FCGjhY6Pq2DZBTPt+rN
R15trD1Bumwl+sUJgMWA15cu82E3YDqtS+dMmtsMddkpS1M2L4OcPL1wePRLfUfhz+6/HqqjtfRA
hNfibY+jhRMfjjUTP01iNVHjd/K92Yc+ulj74Q0ielFFTd912OM3ZQy2NoN0SfAGeseYeth4sY0l
pLZNVsFU/u3WUlg56HyH6DbgEN1NTsRJf6NFG+mmEw2essDkFTrZQRqgh1pvrWpyvHOrjkvlelKJ
1rEuYynpmloaj0faANEHjePCqbCoj9YlCf7yMwDR2zkOKZ68AwbYfbgP9ErDuUSM7IGnr0UKVAuj
SuvucmbpPwDt06Oy3k0+aCswr4yM9Vs8pm1F3NhbChFu3hmw8/eIrPI91rgYj6NBj2C/tEj6HQ2z
bjH6vh0e1T+ZmEZGdIvajkb6PWhnXs217Kr6UAQjLV09AZyyd+PQVUgvts//cd6JCzca5Bw4vzfQ
IsnfU/RJAo/EYK33rZGBJzw9KdLA1lGo2l8i9zxtjXmK7IdEd5t66auIDcn4UVg2nwrfa01buQ5n
E5ha4iaFxM8n741RE1t6BLOD7hSrmYvNE21n96lUzBJI8uTH1lYBghCFf24qBuuEgHuGymNSQzzh
C+AzFRZhfXL/qcAvJRymh0tBMN83ckJpSGERpRhVU5inaJ23Q8Dj3sFRurXlMiqJVbzK5qP6sfSA
Yt+u05wPEeIIOGdc6iLAMI5Qy1tz5MQs2kjhDSzIa8DQRO6g8nptTCe26wRcgtnjoanI0KISYa8E
pNArE2AzSshOMsq4YazmjxV4vKvPnltrLNx1/5GeS5uAb4ayIlrEFVojiBugMcRbBxKeG1q5gpF4
6UEBj1EC4ugw43UZBuKrNR63JBhiHeMXTpYH+sll2oVQAdLD7XzyxhnDY1rD+S/alka6sk0e+U2h
5bNfv5MYWmlv4//MfD7+npEyxQSO0H8hg6thJxxQ3P8Afe15qcHvJtnWIhHzBadObqAO1JjdhlnK
d9fwFYAsI0fYapAVU0ewPH5g2kxIWLJG7k4q+kRCrMhX6pGMcQ4mVojRYwz2gq7CzGIjlbXrkiLW
BeY8iSPe2x1ADFGReseiEQk0/FsxSpW8IiffnFThfcHaTRjjcLT0wbNJWWHNbXiwff8+/ir2P/Q6
3hU+fqcOIf7vpXrEnDp3ePmwi/wcwIAbYGwaI3Xff1BRXADqZOZa2F8nNwLGZ5fL1J6JBTh6783a
8DL5zI0EBbGl1gJoXks7MoYsFhqvrT4AT7dKzpC8LsnvWLpVLN+m8u9+DdbdCSUEEtX66/dk5LNc
9k0W0M9OQtWfyNVZmqhLhAyMOXsSe3Sko6Cs28rAhBxtNPWgHc6baPQjjtftBMcZE549b+00V2jz
8mfAk9WA84UX/fnWBGTpRJI3oui+9bMy1HZnrhAM/1JExT5kExkKxkDaHjL/nbT76hER6lkCSnr/
5WOnVZmXtGgGpenQQQ5VtkDWL2ovgS2tR0Oe3R5naW8xv0ap8v8F6J9mS1JlLzXJaDFpNCGwOEaS
vq5WfZ+pn8Yr6lOoHofthT6SeUODsnHhXqBSjoNbuoVfMUYt6/eThBN1r1OQ/jUdy4IENYrWfewu
0dt2dLG3jFB0ltCe0DHsDMsBwe/clNtILqPzkdfUQLFxHxxb+8HCGMfyL1ScRo9XU/5sOEFkyPqX
ns71S55n1PmHgZHXuvgTX7TVlLj0GPyqCzA1Lw7x2QFgLrD9jX5lpa2fnBf8Rih9CJhxDtLaZZgE
s3CrEt41KDVluRBp3OXtXAEF/XZtiojI9BKx8VZoGWwMJTF+Ls+SCrsjJXyim1gQncrUgybHfYEU
V/5tLGcfpO7pBFOEUQMgf9xBa+jcTbIQ6FUmGPvrOuSpacWVl4bZewIMy6IZMUJFKcCFcmSI3T+Y
isDb5DoKYbfS3breGGNjRe1bHkb5Mwvcak8yWPO4ZXF5NdteXbnox3r7bf0W8+ikKPlmpfWR9L9u
QNQfjYCij0A40zVzpEiGoujMAO8oEc0pMt19OMNxbYj/tvI2dmFE7/YSWjCZk5LKdhmYpAbNch9f
mg/d7qs9TbQkJoamewzcKAus0NTY3f4ZJqov9cmcdpFyF4bjEt2ib1zRJ7rJ9fwBpfhse9eiPWhY
Fnh/7GefeOsDeJglTzP9bjEBxQWUKp27+okcpKVpuU5RbLYBrVoMK5qaJpHWoJD2rlNsb2SZhT33
VwN6tiLzDFH1E9++v3QzCNhA4on984VY+j/6YWRMLE82xRN7ePc8kDN8wSUTGXXnZlgyzCGhVj3m
VmfMovCZGSyqM62Zf95rEuU+xNi368BNRlHgcrewuD8ZDejEH20SPO3YWPZ0CD2kMSkmSBQzaqFv
g4aHkPjF9aQZFsYH4vFNHZLotcLbzQGqIfBb1yn2KlN5HQxa4jKPq/iPdfLyCXaKoqpikvLWyasM
xqF48t3RLYgwLK5Qm9d1NODI3DRIZ9rm9asz6fg1N2Gjj2Ru6dqQn/t8thhrdENyRR8UtevAZ7Xb
5KBtCjagPesdtnRqKv2U9P3rSCNHi/CrsTpUzf+X3+mp4yzOw9vGhzcDNLPk0MtyE7fP5a3IHOkT
vXjrLIArql91I8ht7hX/4AWJbTonWsR8moT4KwiIqv6s8lcuzzTiKEEzX8Ok1GOfPPBQ6RWNb/Cc
/jpkeXY8C312sVasdHc1q3BiEMRFkGDqIAXJFPskaT1E7I2hTVQGfl6SYHBBuH/ON+hD8XuzvhXg
Q6rBecrFNrpzOoHeYFPW64DMfBHj3H0i69GvFcAtAm8OQQkLpOMf8cY1itOQkooQikDX0d+/oQSP
n1OzjLLCNpwNDhA+evu4Yajzi/KEoTPGf+xLCBOdAgOuO1i9VWIVaaFcs5lQjjfT1p89wvvHZ1SW
kNU4Ugs903K7k4uPpgEwjalMcvjhHrbt5FrxPhYIm7et1cNRhRkeRvGWfzthITQv+W/Th4P9jRqg
w64Kh2AG4zi6Om8khWWftmIOFRidONQfTvCrB7q8aLJU1VizQjyNkmwrDaVKhys8wHVMFbLe+48U
ymsEM2ryN5xXipIuxgoUrIy8FtbH4NBlHhDWNhDgGtAN1TDZMlb3VwTj4LOsGZnd0AH9hHFt0A5t
5JMWv0LrDXNPjbsk/gLU2mgVURJyN+8kqv2X7L9jQWV19gaNBoVKdNb8RIMx2LA8TPk8jDINs2uB
I/Rn8hPk5yl+BD1AshYU2TNyjk5zyXYeTrmkkZCWFhaPfh+iagX55UTNRVgXUwpLhixh+gyb9Dee
9szB11XjRgkwuQ2u0jeO0RBKC9jnwNXarjlYp7ZKFF7KIDuKVg1fzpT4a1Tv7FrcNWTmUK5CaJbR
ZnbxWeMNvqtxwudOb5hmnaQ0hxYlYSQJSborQ5WRz3P98Jw4krwNZWCCpqINiZzGu+ovNadzLkFr
x1NRv9zy2zgoXP/FWmcVk+T70zkTeHXpsxUV8B3+cjJfVjWtsA2of8f0PBOW3igFQvA8yKSmDnfB
WM+grGjd+WojkLtdBOR7xh0lPu4fmnp+cKsT4uc4f/6qKmVHD5m1X22y/7LQj+xaBMpHU1pnbE6X
VFMFrBhNHDqc28fo2pLYmJ9foOjwn8A+KNdI9X7RMUEp2YGQl3a5q3yi71QRTTCYS7JpRQeH9w+A
4JhPYmDLvPgjhOIGdJf363Di65LlfWBioUAjfsbvrxuymsd5Cs3VsHp2INgOboSu6QKQDWXMGhnC
He8WG8pWLxNv88UkcEM04x1dlr3JW/5iBQBXubgxABNp+dXV8Xv9Qap2ymN0quP3LCFkRXzUBXQK
p9GE2wLOaoWa2wWI7y8X6S74wQVKhIDUUIPxbv4qYpj4E4gYiKqyH5fWDu56W1SMgAmOfvR+BNE4
Q/O/2Yq8sMp+F3de5I+M/hkdHqUFh/AHZd7BK9SZ1RsAhnqvcUCYAoL2vdHVDa+gfy1QsKS1DWCH
gE3SG44CiebKTVfN2/M7DfEqkMb+gtRSAulUjMsPcbuMRKJj8bwPuZ22B19QuJ0m7QU1kRkKn/bK
qVZJ4U7Kjufnu6lUWfIGOiLnF72mFVh93xMgXcafvNA0YqlOO7Wj35qj/PsxG+nC78UzuAblogcb
HtfdkvyDFZCxiu3tzQftLhpcACgk22shLeUVquRB0zuU1zfEWqjEjOrE9rmCZoTxfFqf6ma3Tywo
RVxp2ekyCnmdhxjsZZ2MZHhRcxY7gEAOMewDPnHmIA/0KCxi25BdZ9JARgYoboabVP1k0CnE5ZYx
At/CT8Hof4SyZ9Y/KAUt9XnJfrOblj5/LyAgq8FAHXOTetkZjKua8dSUNRRdjqcPDe25hZchdBZt
+A4KiQqyWVi0RGltXwauN+qJOzYSPV9gnQZClO37uUoebDFPPiTk2gmsYhgd0x/evPo2YTaULHIU
ie8Rs3cbX6Uj6N857OAmmFP6US0MqB9kZ1jfARTK+6cE41EYpIASyW1H9d8cRXnZk8wRh3YwOgaX
g531sOLr/TTat3o9ofQwBgv+udhlm2DR41r58RRLgVXDa4tK2oleYOYbWnebNbdBu8vbUU+f5N6g
S+jorOg8qN+DgImkQTin/ZRl5CeBEGS2/AvHMwZVAGhLX4kaImk8RvMRRbUBz5g4XPyIjsgpE3XZ
b6Nj0erzrXaNqeiZhal3aEnwwfEhNZ22nnOQuQ++mWkQ7y4Amh62IgqpLg/TGJAf7IdAwJ+IYVLR
zq17qYITVPlcAZJKJ9Ddu68rmEJnM+HuxI+/SsY2U/XBozVnOIS2jQ+WPpt19yVOKlEjbtS0rd6g
2tKwszQvkNr1Hdc/MG//vnLSqjhPXnxh6JwRnAa962hh2cuJIrztFimpsowH6Y2hnyQnSm9ZkOL1
KIuZDN2WHks/6JxkrWhagzsi00yvaKyojbmuYLHA3eij7P0kOGHKjkBMQ/LCfs3Zu6/f0fiiMco3
6EtpqNlOwgxsZ0dVSqA146TV8RTv6w4AV+iBauXe5HI00avJAoOYtclB8jkoE2mR+7fteYn8+XSO
4rE3FbDQsFqZM4xb5XIDWqvniVb9e9nVyB0+XWmkMWtkP0RGWHA+rzCBpoZ3nLqoLb41C1AqvY5p
B53/9VTfS8mfAvyuAwFuS/B62CaN2WzIa/FrTrluPzzY73YFO7TLgiWxBuFzpe/1SmolTqygnysn
SuBDKs8F40/ZDuxWBNdBZHtr5vH5u64vBEDOdE3DlW0KzVJkySXDFkQ6lneH1xlFuQQ6ANzIwi8F
4a1By/B8UrXeIIxnYABF+HotXGpxo1Yt1jRKbLK1tWBrallcQ9ZZgH5fgZ4pBdHfCpUu5MxtNexy
IQdmEVtFPCipmOqWM2co0paKbLJmhrDlgb9wYD1QZCNnYWkVQAU6j0GhhbwYM6tgsLFHJBNfsxuu
IxmY0WU6pT9Y6Jqh2UCKC7NMJYWYz/8SFoGK8VCL/osUVrsPazVk/n8pqmZgHkK2CF65D+2xM1Gi
VMLwbK8sS2che4O7tdilGHLUbg1PCDrbw8y8XL+nzUewR9BIBd9IwZvTrBfZzR9XGbCVXBrBoLTK
0WYUJrzcUf1Lwniuaejk9jeRAOFsFMTt1eOaK0vnwdXPtiESX6RLbY6tUAPaw9IzEfE3LYrz+Uno
EzeW+49BoVkgAOYk0JNOpTqmd+eCOTQxhHERX1iXplCg7OxoyXBCgOZB+MNE6Zdw3imo1AgFil47
i+ouZ72qgVFbYY05rOBAVkOcUn4T/KuX9xGHzCM59WXQvXfRori3bqNHuOpm1vFqF2tAC3dsjgJE
U1DjqPhpjTMvcuxu7FLQv3mwMvspaloAcnNzKdgRD067RJ0I9Av7cj61ubfL1EVO7TT+iixJx0uC
n2c9tsqH0LbEMjq9/xU2TxFGQ+jnDajkQzY2JHYKY6zwX0QS85OxiQ0l5ALhSZzSLO9cOFOJbLeG
XPyWSbqi+xpKcgajfi0d+LthHmqfumYjBgYAAt8GDI/Rzel8WeLOrEC4DHCuu+oRPBaZeGTp3qcz
1K7PHba4T2wGraCqsMvPx7ysaOHfiVtXSMDpTRikFehIm60A7it9bXp6BKSUeN8OcpoVCd1g/Uw4
MPt/NeSMTl1/ODbny62xs9COKyzyjlbu+HJNgmgTUkiFR1ccpi5JAkX7O1EV64AOQedYbTzIl+Y/
ttx//mOWBH1PyxCHzW046Oj/GQoAQ0WjMUHcz2/T7bsjC9mcut5hssAxnQMW0Qq9QsXPiW4kuRIf
VEMHJXGCjpopaK5rSaT1FkLo/1b7vQYEopMtK/2uFatpiOP2apvOwAL2PBCj7ZYgzFBgotVmyw2y
jSUk4iR2TTJJu+Y9ReFA/Yh3gxiwqeZLTMauYCMYGffd2R6wgZAfRCKMSC2jRzM4J/79hfANrR2C
LmqNNrMnLDmfFpX2F1fOcos0XB7IswSboZe8YYtNYk7Cw0pEFrwN9nYwoWNWMEIzkV9ReUn/gpvo
YyzgZIe4E+j7Hhk9Zapegup+TP3bnDge+yPsH0aHplY9gTyk12qW69FXhAg0PnU+YZW4ndi1b1/3
pwYuEAvJptMNMpXmY6raJe2bLqeoA4kfExJnI/gdAf+B89d9VPEQZKapR3jDKWo+xoaRfDkt1umu
YM+uFJUaWUWXV5JMsljQFI4+eOJ0VNmEY5TeKOPK32Nxlg70aUVYFXewZdFmtr3jhTB+kMHxa/Kz
kd/ax5x5lMROtuC8tcK/IG5Wp8dJP6DBiO95z7zwUJDC2jqNSc54bR7Uca25M7FrhJ0IMXDnkDOM
2VFveGVTjCG+mkL0VAUnI25Xu4lWmkcOn/50iuGOPlL5twBaQpZWQN3sXjNjS2zMpUIE1J0scb8F
aTrkk0CPVahMDk2dViCMaWMXLExJ39fXdOkJh0tdc+hwOV6Z4RzyHghR8fCDdUBv6tVn30QSgULk
ou87s55Dhx6JskgooVzefYfzVe/uW90c/dxDwo6tKmBQUlKlbc0WExxvzjbi1IipjMkPWGL8I2Al
FoRnFwvTXNjUL+E2ONEkAiUTHbalTvr4ApBAel6biIUzeQWhzn4f5GadZVGYeHa4XFxP8g91Xrkn
Ls1xfheEuZDEkxkUiHhOip20EFlTsUFyDIs9MaHnpZDv8HCOp7gYq+dqVk93MDlwcakITxS2p1pK
2kEZ774xy8eRTNju8NUFUMMuKPPL+Nw07zH0TLu15ujhc4FL2Viq7EdaBo+uj5R5oiCQhZ80RdJc
8dxhmlcbCMkhWxpExLEri3Jmsm54TprZlse0TwxuD+PON9arrusTIl6Mzc3IjX3Q/FhsZcFUZXuy
WwJwu2FJXn6Ge9kiD2bEMTclqKKM4w7JDOtmCtPaYXwS3ylJpQDHo1njO6/j5b6c2uJQ48Qzmuje
33gunhgV8hK/F/N825YJXSHFh/AV8yvWsp/bRKLvdbHrGHpuVvP2KvJ2N5HPfM64bwQ9ZNYywfbr
gaZEOI3+rjxzi/M6xiCom3CIumivS+3bYTs6SbD6iteXfx+g1ihzR7w5qzAkfnJ56lrW2lftzJCx
5VkUkLK9is6Ak2BIS72sKHMBy+rPhmmauXkA7WzFNQIvAn/BX3EZ59eOqMtOqjIEwKgDo2UErR6N
3jKrt5yXluhxzMZEEOK1v0C9D4iwGtQjhDT7gvXxAe8Sd0u3+hTg/boNPr9QoumEcEO8hMEk++EA
69EKn/bAJOV7DLpuWT4FibRLit2oVLbTk2h7vaD9tbXaJQ0OZuFFjcgSFTxMBFm6z7I0BB7UqHEf
gsIfO2nsKg2BFQZP6uYgL2Bzvp1RHnLSpqnj/fRBCHlOpjcT1in9OPQVUPTjxrUH8GSDNVz1g5S4
wv3Bss5/tXF+hgpkpjwAhpTo01HpAm8vGohaYAJv+foH6Q3MIQ6Xb+9ME9V2hio5ZDombIEzOC+p
NNcBQJEQ6rYvw5IlVOzK2BsreVbroS6oVxNgCqb9/zy0DVSga2TiiT+Y+HbhM+8Hv2MK58+/KMs4
Rxq3A0z3GsnMfVU9M4du4g7LEJT5P/x1wJx9M/xkXnxxsBZFZH6SLRDk0qN+CAIDNLqWeMGIhGlM
0QEOKMNRnYEAjLO3C0+HELI4PvVc6jEiq+7TYPhbMskOyeRNVE4tak7932seg+h/bz/gFCi6QHAV
isGL74kWOKJBeVB7/2/Yz2ocNcxxawydfGhjU/ZsDJD7qu64ZHpwmgM9n9MZGFm9mmXXmY2RxIc6
+OLwthpWoxh/aetFJL/4H/zHhiXMmDgbXNIm7THvupxZmS/U/61ATgdKVJ5kyXeGpbtgMhXORdog
2lJXuu8nE41Q8u7srmt/nYzSUBM4NkJHUy2IEyCuzxSCgdgbze347o/CG2eIhpgYiXnavTq3ooeF
MyO62urDBHxqIlX4O0Qxno/H9G3J6QK2pvk8u35ymvEr2gKCyOKzoE/K/c96fXZNV6DSq0zBMqu1
k/VhaIFTbGLCZR65sN5zm13dWTCKKkbCY76NWyefmhbkl2oIXl/a3MYb2hQFzr436kxthRuz6pS3
QeNOjrKknSDBMtBO1ZqWzSuIXsiBAqIzFcFaXYhS3uNVwX3T3XIbh5bSeDpI9coOjRB8GleeJrLf
iMDptZBNbfV+Y7pNLrvVjS5VZZRkYGGSZ+AdVdNo37XWIi152Pzfeozdi/ZSPMsN0BpKDuSnBcEb
044cK37OxmITaoIxSE+5L4WWMgDJJh06Wr0K1jm53L4IGzoq52dn/iL86KXyIUti18Y/JD4sxv/1
37DiD53shrn/d/PygzHFJMDsDBBkfYt/ow8D718HvrFN7dnLL27zrRpIglHrqsC2mkhx6bg886aK
QGhC9zo3CrdJHtSnSKzDGJ6z7JtW+KqQ+otrYQuidsmvvvziTyUt3aJl+pC5JOSnAT5kFQofl9tC
i536ae9TttHghuHt9EtkGKp8nvwtLGYLuv8xVgA9j4W0MBivoTO9AQkYEIszDfb9NWbYo4p+cLSB
EMUwtwnd3zwZgtldCRtuBo4hWd/MpC2H4Lo6C07SCtCZYHB1WrAVMGu1YES+z6jTbuERasWuAfAh
M2455VbmdAule3ohvc38dRppA7mkWl80Ci4QZ64YOA6VvDWg2B7xJl+GSbfPVo/ERb4IaV+Qo5ML
XH3dliFEDbTKDhxeaoZOu0H7+tQqdD+4B04BZjSfmm3159Lu8mr4vH4YxOcFslY6QXg0/PqaMZ7U
JGwC6pOsptajYLRWep3iSTxO+DlCbpuy3oHvji+7Vk853f03DQacDQBLwCHv0XIUOVMDstE7PQUf
0praL/6bC1FkfEnSToX6+oPRftwNAkzdSSq1ZnPMaCl/8O5fZZBW9hUdHsp+j9fBpK87JlsDGbaO
kd1djXuLtkP8NkDpimW8UmVPHVpFyCCI0C9P+CfD/cex4WtrYcx+Kn1lCnnwPOze3EUgED/y94Qd
tO0i/nDcvjbXevMlNfeUuFNbm75EgijXmSNKoi5JL3w9tQM3j+arJp1Y6/hBolh/O4drHjS+rmOJ
ctGSviT6RueQ/AWKC9a4mgzSGoVUAmKqJvlXYp2g+XF/7OR4yGfLrsKhph88gZgXqGxX2L75Li7R
0wohPMHJY3mDqJEpw7vmMqb8Ha3YWyO5fRpjjLzbfgCksWA1CcaCwku3eyQcBQacPRs8jLC/gZ0w
+X2Chi+hQQP55PeZ8cjrhyYJswtA5Q5R9r0Y8pyUavltwY24x52f0Uk7Wi22CcH7ZCEDMAmS2tt0
EJyVPepj1sfjQboQ1cEBPKKEMg+Ex/R97NuKSkmC3UvdaDQLWRZglXU0necR7SyNKkTvoQD2trmL
dITDYsEkmTRrxEZwL4aysDwojKDdmj0gYzZPQHhwUcVU8988WVzJaqmF57G9ukqdcgqNSyp8w40y
jHliZqjXkCR5CgaX7hU94fQ4PXjTW4RAOrrx9WGqa53SsPYDjjdfZZcMcXP0S9KcSk65r0hdhGto
Z4OtHngWIwe4PAnOHMZkPB1qUGHbwLQXM83QRffLt339jaHpLy6GULFY/n5te9cTpkxcpm4mlf26
Ii7DqzPyMs3QpnkvE0P8g46z29feHlmxnPXhT5aWn0/M+zKW7OyhcqHNAKwp9qhw9e+Do1o+D4za
iml61LtIQFfoO5JQfiM5Ngari1NZAEgqHe6dIlEZHRjVdWCrhO7itwRnOErSz+t/n1KLTrtnkgNo
EIs78QosJlSvKOgXtge45SzEY/p0z6QECmCP/g1bD/RIUlq8Je/eYZkNzRArCP9LSDjbUSQg6nUA
mWADu6IqzRD00VAWO9X0LpJARBxwGf4jlQSUWEeJLm9fIIkIw13oqE2h6R8kxxZPZtRw5+SIWON5
SxzVoz8fczRg3c3K1DFlC3ZCZ7mfmuv0/NpEWwOZTCGCRX48yay0CkwTKd3drd7SnNW6MV7+fRD3
4eofTuNcINL5GNzdNSl/3asQ/VRRzdfIevqChjgEJ5gANA1rPKxjd7E+E0ps5Ro+HMdN+66NF35Y
f7WqQjLo0TjqPj+x898iYtvYYi+4zF9nfZeTw6E5OqoFXjlESZOu5U53wzopKRwAZ/Hh70B6HG4o
4SbVrwrXf/ChAFSX3l9Jaz0jf9t7gTIWRydQ+38QiKW5e/UVut4zx7UTsHH+lZF1CkeotBNFpK8A
q4X5G152un1Ay7Sy4yQRmndsGVUU2SbF8hXkiXGgIvRorebK9ZwY9PX2BQFZ1B/D2toRIn6TxBaq
6nNaOT33dXIiYXYKzyxJgAmbpZZzCZK8ptk/1NMc2y7arslVuMqehjGh6etZmqGiMOR4m6S1eajq
2NPLhsa2lRWTIa6Rr+8jn3pCVbC++KijqW0ZMu+11nhKFwWr1IVQC/oYW59pVrBmKHTrq6ZCiUJy
BMAQEvgxl0oo1I3ErSiWitOBhNat0kL+C4R8OisxcsCAwXzQFSEHmkAu0ZsEDm8eD+S9Jqa7IKMU
yIIDbnyvQsAUB8Wy0BA7qZelJQ52JP94L0P4U66mpJWXKCx6IKpJ726UMSNZLWJfH+PeePt1qQdu
Aeau6Nxb1wfsqWLBRtlR9sh/8/H9nZySOGe0f0dAejzz2fPQTfOY7EvRHW8l03vKiACQSxr1OlHH
b/Tm4mAzi84XT5Pwp+ssfIEtahUkio3iN4bXQy//RfLVVpokHGQc7pcb9tnIc/fipf+pOBMFbt8Q
vKN9fy+yErXlarKtXRL7ciYRNl6R5mchmmCrpXwmcXRBvY4h0y32T2XFcCxjk230jCTSvOx0XizZ
s3FczTEk1Qeaqxq7IooAaq9q7+ccX9PDNU3qvUZ5pQTYw2rwCC4nUqqDUMivZ+g1PkN0mKhwOGSx
5ENjF0YwS9tqtYOt9/dDdSnaek/D6myBu3PngyU70EyrYqG3QTcopdJb/OBeVnb6okY76Zj3AbRg
6cd9rjqpDmnbxSfmU/d9FUBQPM0mEejxXKQPn6D+WT+ESCfrdN/0VXfg15kfhm7Ly5sawTc1z9jt
t4WflCTylU1wWbWbVMprrzjlBJa5iCyUeNeDkiF+luNBhq25GN4WCu1xUCgiqze9uHcG8/+mKOmg
QdkKgozuTPuc96cgR5oL0QSJMLHt5YTl4/iAs2n1rm2fwj4+qv6C7lpTuNBnqZKGVHeUb2qJREOp
KA902AaiF1BdpOSdJUgXRcd8kiAkikTQIimRbZOiaSk18IX1bBHXdOLjYd2Svc28zk4QKjcWcM1f
7ZkPt+H7GOwnaowZmVTb60onWksGcdu8zUTlLN14WRvKfSGOVjuSNux+4LSjnXtxBPCwUiyUBc9n
EcVv3/e9OJMJGXPn6P48fuJvJLJt6TvGrwTq+tvD4aWsXFXFvLB4eKd+LXebyLfrgmkMX3wOGZrB
B0ndYU/dMBnAfP3NSOJSt5eSYS4Xn48yV4ttBQqhkZUPQi68FbLizMWfFW19l37Ve3oTp91ye3Wy
YIl/zGVHvWeqEjqgxZL3leABVYrupASkxw+gtOlQE9hPcm7CPlvfl6ekSdrhDABlNm0RkfETEMu/
HI/ZuL4GHfpg4KNA/aknEzHofQs2SD2ZOJz2He685fji4GVoLNrGttK4N8GyLH6Qyyi7aadLnLKx
jSEbwUYPXLGBEltTOKABRqY7n3AJXjJIyNuVXtNpmA4cYd4wTALdBmp/J3GbcD/gWOYSqFjfY9l/
a4yyZX8vrROnyufeBKIKD6ZwbkmV9MbesmCYRS/7FFZrKX+FMGiRhP64Xlyut2JpibWqsJfkyhuY
o1N+xMVs3SsGWpBZlf4X5y1z1P6P11c/sVmrfqg1HE4G5FoW01t3pUmFi5dDIY94AZg2yd2XgZ1O
BpwoI0n0tbZqwkLt06rBr7ajVPo0d2Q6d+2GtaoY6LeVAidp67AmHYZ4FNNSbGsPxhq0SmAc7H2L
lJ1atUoykv/GFtD4l68pYLXaxNwlySPhw4J55JSiShVM6R8xwRrbyvLUa0//M175VJa8d8FunIOf
u7ShcS+7eN0NsT1sgzfeHJucEsG+ujXHK5+6w7yvYBGsUkHWh5tQINjrP9wONVospDmAQhDqPT2s
VeEnqhu94+M9wjfbxcRbZjXIuMrxumLgE93cHd64Me70Prdo1y177vrEhWBs0njhYhZdI+4iLGXr
Q9y1nyUVJ1kqoqVD+k9qy67bRLxjFcbBISKYbA6e2LccdOlykPUD9wIBathvPopRh3OS3ZNtfN5r
uBlo9uG08F7sQ0ozf+FE//vAhi5/HIbA7bxTRuggcpRKmWOSfau22CKfCtw2FcaNifqJ+hSZiBqr
I4QE8W2+WEj0HBdo5VHDtp861WNsPXcPaBDwOGTX3xVEdJfonbbzXWAC5AgWf8clunuq15RBYMLK
28pE9zTySzA+kz3fOfUMK940M341SSjg6AXZP3PkxQzUarHQ42ds7ouLCOMTdbiDW79TRYarLuQG
7bX5eLjFh8AUaXV552RKMA7htxAIYRTyGaaMIO5zRbA/XIq9pClQvga6qfheJdrJEE3XVqapPrrD
7f1/G4SizwzKt3jpPDGHOTsSu2H50vXwMMkBjAOWZ/aaDIkIWgi6UMd7MGJdbTxZGzBIhbIFY8lF
EIE3ix/+5S1yB63bZtjd3w2HgK15p6plptmXO/f4IFGVzXd0YWgULt9v7ewvLVhY9PHQXOpgNYT0
u0NEi068yRgdymIsLuTCJscpiO9WG9czxE2Tlv1YXJvLEi/6YD9KK0vtToTQHQaH5MRrxCbg5ERE
6R5ePl2WC+RjvAv5ObO79lkVWyeXQREQEj/VFn8zSm5tGgfURSrv/uy+v456TeQtRf85zLmcO6p2
W8r/B5XEQPDL34ViwB1EghXY1liDoFBQimCQ+70ZGTjTVk8l9XuxfmCAZsEyYsN22w1Aqn+ur7WC
yVhopI4ujbvhdkEh6F1l7/MEwKoRzrLAGADJdznA+Sgp0lnW99sLDUg4bHt83UnUrOpsrsv+v+pB
PcMEndFRlvHHsmpPjeRWepeLFi+UEYMGG9FyviuO7t6ggO0zgxeik4aAhQmxyHoVobno6CTa9Hsu
W8U6pkhTvcu4y/G+aYd4rLD+zqrQL4hJIf4rrizQM57/291bBBZoC0Feiugmdil/PiyazVpl4LxY
bK1MyJWgeqkITqjo3l05d3KWI3oFx9UViaXF5ipoJLAgesLdnVrAriMTh420sLfExYpzyXxqMYfo
Fbc1HjLa3DNlSwvMTlITZZd/pX8gGtTljt5ogBfVCoh14j0PcRAC9kZNki33w4uwYsAhOrSlXLu7
maDZlvMILxZHps2wzZidgXO7tmwHb3tBo5UuhtYNCbf7RryosLu36abGW5tvbu9B+VE/7mhAJHpH
A7uteDMuyOGAGYTzsrg/M+8VF4vwPwb+P2yztgGYNPkAudjzNeD08PAl/iUQo+yg3mz6hnNma+D3
kHTNs/MRf6p3qPy13iCrfkFpWMnZd8W0X9MbYt6YOfU1vSXXzNZQJCemKctghNm9RbQkhTNoIyiQ
FHNTA4H6pg3GwMAYa6w5IuHgxD3mau5c+j1U7KPqt8yRMkytcBOj1jGe0pSil3T/8pGlbbHcubwy
KoBWH5jkQKa65f0swBSGIZWO7a7S2blQdcHiJ5xd7RiPaZjzCIGzSO9s8gvLYlxY8AfDpBE2Zs5R
nGdhvyruAHV3Ju5h2JXUy33Zjm7P+pCSuOmJRDcJgjA43VRkH8JCWNLug84hL0fCtGCy5e2ZOP/Z
kfXRlLidgbS0HiKN6hN8zbS7NRcNK5Y4kviBR28dliwppcmY12GVbIRQRbjoHwp6B+ZrQAF6qurC
o6ZHiA5OGLhMgGgBnLpcPUIbI+Bd3ytx/mSqRHmvy320tcTyPddXLn2Y7qX+7iSCRw3SQ53Udc3K
XNTKqJmsgGtSJAY+xzMCRYYzs8/cMcu84JVXZgRpFXpyrI8zL9PkfFrR1iL9TEjbPygoXGEOCulU
XXDJnExcbvH4dXDo4wVxNXrZh/ZpSessh246+ST6pmLEXqYEoDz1x36qyM4NowJ+eudzvBN0OGG+
HuwPYtdtBYl+hh8n2Kb5j0MRNM+tEhTKIIMPnDd/nceO7ypsrjqOQGm9Pqua5oU4fYx/G6K1MFXx
KUNMEA9nkW+A5/EfusYx81B0dpasmUsnVQ3JEUBaYjZuTKH07krFA8nfRsRv9kHbkkR3IPyCSX1c
GXMlNCvR9Yv0N7rxyU9FemerARYS3F+nJ1kMokTPP6ZarSk8TuOss7zQiP9WlIvv/Bx29E3C5H6r
RvplhQUZPr2tPNNiRHfJhxzSi7VI6EyIdz8UWsB6hjUNdkPzLSVYAjgFPMv2RnIb6d0FqVYPSCut
YKpaqBrdJWwdIjXDcWGexvSb1L8wHq6K0ai9eWRpHZ35+5ZPqR92toNQ1s1g1TUpb79JIFrh79kZ
r5p2YlZeAJe7RbXX+Cj00/NkbaWShvOKlJ+VkAibpA9zT1tqwZGR39YF+xcn10X4udoXcsSLmIwN
p9MYWv9t6Og+DFSVy3YJJJTA7i4gQ05fD89UJmFXVxBlgqEr9iqWZfA1U+Zt0UfxzFWG/9sKb5eG
5CicstWAgdy5fitJITuJacxcNyK8mv5MT4vwS7sxaL0nVg5B77QZwLHSEB/7a6EkeLh+FVV9J/3d
QZTorsd/xU73LT55n8lFuoKn/NrhRacv3sJkPHt6QHHFVS/oPfWafCwLWBXA3TKLeUZ3sVlNRove
lTyvRSNfI009V3wBa84bq9pTUXujYTzU+kgGgCmJkmxLlohPXL9C/1AlP4HbZt1cOqbEFtNP/GWA
MJ7fs8NM3J/lsEFwnCz+s6rJxjjNxQ9GCr/h6hbxZKGH0SGqWbdiroWbcyFWzVLmzdOEoOCBgX4O
wQhmXFRjnYcr4aRVYqdpwi2zaS2K1F+qL0esuhZJ/7s0+8JVTDjzo1my86MQkbajitQ18eAoGuqh
d1xY36dkfNPcog2DaOcbEj1tr9esQpCu9NdNORTGdpJ1bGEMHQo+z81Vv7FQatW7RWVVlwy4PaVR
YmUqdsKTT3uJ42xbbCBFoCj1wnrXvx3mB6gQbsKcFWRZtoLy8k6uiSW5EPy1EzfalREq7za0Rvjy
AGILtQLv520oCeB34gxovmbZxt79CkLbHmRifTMtBWYff787HZuYAcjBxun1IyagCDPKOTPiyjxV
oew5FFyvuqLF59axmRfp6pehy34BbNTrdhwWumAvqAeeMss1ekAgwE7oxZSIuUTIVUmeDbiNtcfs
nFIezY5TCRV3claBWeu9bCCSbwBFb2PRZfbm0ntpREBmUA3gxI1E4EPttFClNwutwyNrl0NwjHAi
dVao1dX0GKJmSyrXfPw7q08c3t5JAKduMeOuf4DBA1CBKci7Ul0ynZ8J+XWNmNWDE41DTMhIe7mA
1MGhsN3aythlAMjFrPJmTADJRHM8kFICYwOHu1ENGcdhfuiHjCUQvOJfM+Lu15MCkzEXfEOHb/zj
JimwEOyVFrPPZRDRYnoWHNA/3D1/BjnJWBzILTm5ltqbPQR+3TUmXbAUzRKN+H1gs80tN+pFsH07
FrNwaXFMRv7K2WxNf4GeuxJ0MSwKl19vLT9ddgwY/noQFK37ojFK9NuLA2G7DCwESU3deA8Hn64S
f6fZlYUQOy/nZ2iRKMQw/6KVqaWxyqp0ZerIDJXkGdts+igiMdMbnJugPQwswpn0Jobz3Fsb0I/7
x9wODyqC8EFNGQw2IQq4QqIVCEOuUai16iP/4Fq5L+NjCzQyaOiSVUGjOhbqS03gnxgD10B2bex1
e//oPFBAVMvHLTBQNJ/sSaauaBtliGQHctB/ETM7SX32uPbmF8wRhe6MFJBvbuaU1hctJpRY5HXI
396O8mMbjS7a+RCnKjjvaSbseTB/yMJuUA0htPoQgwMyi7oFugFAdxJIxfde5eSivckfO897MbeD
t5Y5cHmWmF7BrU3GYDaxSP8i6BNq4iWxsStJSK3AOhNh0lVTjSsDEC8rWr+lZcwdMSCEGfuabwj4
EMg7mgoZtXyxFnU7TwQdQaq76iii324eFHiMrc1So0+fSDSSt9KYV86wmIkbMBO05fSa2IdoTjuX
EAQ3HxEV+wJYWajOBoHh5eb1LQwoFHjaRNO/CgNnPkG7TB8b17WTEM2O879KTixezuZHW9xTQv4k
te1xht0CbyMMFDAKs+qJasRXNTFvxjSv0QbTaDjkDejmLJM07rDchsI4F5XbiKKB8AlpB4Z7hNRg
2kInRxeU6+F4zBbLvIN6xtYzYeiLudeAEZ+uS9/Q3IKG4C81Ehgnb+kTSjYvGbVwKjbF+ABW5AhQ
SMQn+NvQLnwC7OEuYp4wTfTQ/LlslVZuzEXHw3k1KEk6MJ6wpvxOtmsJ8sMh5F86HG25KtpLtEpr
7b43t5h4ruA7SZIRovkTB+30RFTuZsXiOTTb5LzHOf73Qfdm2NW8gYwXvV2JiCnBSx7y9q7PPwug
7zDMLsFewdNJ1nBAuRjkt3MbOSWn/GvO6sv8Un4Ball0/XomMBGVNCmzHOMdAGr05j1lbE0yZtVT
0sTW4/7k7NiDwrKEZ03CD9WpzxzQ4twjot3EdjJPXM6EFSeGduqpsd9g7hIPvNb3kXinJ4Q8jDOd
67skQGh895x2wK8o4CvSr8z7IuA1fnpshLvHfBsHECA1RhK51D7SmuzlusV0OuD9NCPExqo17mKg
tNEqfy3iF9X5TTmd5bOp+1w26sska5a64MW7W8XujLPFDx0sgIl+afg0uelGV9F0/Wp+PoBCSVS7
Wpzh7B0HNmKDGmOiHGHIvGYYL/JDNC6v35oDqv3DOsIlx01JMASV1BphQSNjaCbuOjkQBXgWOVR2
WINqG6XGf9B3jpzy7RLF0yKwTuXuo8j7VwmRwo5e8+ngvitQnMkHTkyaire4A08CvMe04qxDSndE
kYaBeoZnZ0CtapjNN53Q5TU2a+Nz3fbwhO78V4hA20/lop3y1f4pWELRMqkKJQNQIeQ5lV1N3j4K
jzZnl8L7rSbpNbnOTiNKtGHFcwricE8xYqoJO+DUYoTdHgIdvtSNGWAz+GG671lotcsFu8ANsLc/
Fb3JdzXfobTqY4wHlMhOMGBWXhp9ngJky2yCC6eTcjtrvwB9gokgD2VSCuRC+uqEijUAOM7c6FKe
8Kzbdn8CpPruqRrjQDzULGG++7Rm7CseUONA1kKmrZb3voeIYl7p5+0UBjvxsZ/f9KtxGokJXclG
Nw0LIcpO1nSpsO/62xdHCfMtF30/Nvbl3Zkn58e6qrzKWM902e72c1ZvI5yZFfs9fpz7IlpuNMey
+njEyiScKRUhUVgLpyDBM/ZIJwwIuqs5aBfPuYkr3o3S9d3pB6L14Bq4tiFRFKRM9uKj+xeScj1j
PMFZH5E5w26Vbm4ADelf4X0wqlxUTFSDId53wgC3Gh5cbJUl3GU8GDIFBCjjizlDqaAHszTajkGv
KeKz23q43kIKBeFWc/nejnenXbXJzKqP5ZAMiU07F43C8vrn4WcsroueKMR8iCQWKpKj6ouC5//O
kplQk29Q+V5NqBz0ozDL8uPwwaPASqIvtzfPJxtmrH8Y6Pfm/aNYGQ/npWB8N6v/zcYCcKJfcpjS
OpNljwvlgYXpZSiZdnbg83VbX6i1Xa3gtiVmB5+R5JwtAArYTfqOLXq+bmm8QBuudLsXf/vOeQNx
gtu0BDJpyCYdjxntgeqlpfDEG8/zhEMoiT+ENJfZ6grsc8gO9OFpnFp2k1IrygQP5OL08vwwZg/S
UHICtcsNlQZybbFd0vze8NdxMik2a3Uo8Rver0POpHT1AQtX8GsM1RbWal1eZqyjac3V9atcFOx8
fOCMHK46z2DpsrqJVeot/zdJDpJwL1CuEGPDMccS06Ip98wu8HfPhWyr5EkBzdzgH9hfIIbXS+zo
jSbVKmbKulvtxnLJEWCHVKdKATKC/4+H76wVsrBNMyhf4+d8gtlvFUjNiH9HMy3cz2Dsun/H3+GT
FNrs5Do3Z1qiIr4xJfWaQpyO+ShxkT28NPXzQ7i4tFq8b97jwoBMfFSwYMAB+B5BTiTkAfzNOOxW
GHExjhjJbVkxJxKxzsS4c3KHVUCfIChMkcI8olDKOsuNc5dLGvI+o3faUcXLHJVyC+sxI3nifqjJ
aL2VxGvNHOAljWHV0jHSMvyC2MfvzW3e2WrsqfnyoalMft2I2j7TEN3E7sXlo0T7dMhrLg8gYVew
Xhs+riDUiR+88mn8VFpOUtvWiPuGQZ2S/YP/oVsG/kGrUeDm4U2qhuUkwEU24yulXHDI9dDGmiCb
u14U8kS2HEX2iE4TrvdtH8FDuohf9MEkINxJLUxBXKfifYiogKBAJMjmDQEpYEsgLp+wsWqI6mv7
YPFRnVHmZly3J3dWtJOJhND+2lY8umxuAUjeMFIqopRpmoq+ce7usPaQ/VMC1E5DCPueWZAfYy6f
m2+jJzZT10qPjrOQo1QTkRoc/bPSVr2BSsjY7/azBnHnrbhYWuETg/XG00/iQHcW1WOun7/3DV+E
16kr2g1dSmjhj+DYhWqbtl/D3IG/OwemiQ6Kdnnx+sv+qMPc1yp9Cvy/msDcHGip5sARXRiainWg
llbaHRTwnvBVZJrzNjjw5pf1o/LrxwBPdE4oOB5iupQR45flgIaKPBFXyJB/NGmPFgSXU82oUY7e
JKpzsn53YhsBXiT1Z2Ypfu2nfICT+IzufskopirawcjnycO6trCm3RfBVkRZ+tBgyOw4FG5lQD/j
YsIhFmQK6yyPLxFswRePFkH1lK5TktYuvHnsqKDINMIAZkClPFXexoJATiG8HmqA5T0x7l+aiNi5
kFBNYqq14SzvZ3573n2rZmGLwyrmoUfuGYUv66i9KiNXcJkOCjs0ymogFRyaJTh6pi+f5ZdTsLmh
kji/doef69cDexCR+uPcaa5ba2oxI1oca1sfgXz9SLl0vDNQvDq+8RpykuJgBA6CwP5T6DGsAqqz
MIvS9SyM2BJQytQQ+06o3DbaN8nme7kpKEeHTzhwzAO02mJ7XT/1nIIoZSStMv+15Ow+OU6kNliR
aGeJ8Qrl2aC02YlBOoOCeH2LhW+/XJd5+r4+WIjEBHElibAbUuxhZjXo3HKqh1Zauyteag//ZJg/
SETUzhnkngyEXFfLzcR2YaXgfPdb8GwG5knQMvELvLqVrWL2hXZUe/bOL1OL9uXQI/RGIFIVJRfe
FMNFwth7NKHer4gXRK8UUofBpcx9mY31/v0xYXlHRdDRC0Dz+VB0bjNKo++WU4Aw4NbSRa37GCEo
4N4lAZnOy+l4sCKHeNlCgC+9OzDeaZ2I/xP/QPyMmZ941qhtfFrvnV/KzhJFHm6bktMToOlOZk71
yP+PrCdX1XRMdDk+spd5Se6iTGMQj2UJ5orLizdHwJeNZI12IaP4uBGAaV5LyWYmaSUIF9OLHbwK
iIEB7CMEyfygpPh6Axgd39WduBAI/ZPlPy/saPppl6GJ+cNQ5InyZf+Wa7gIQcdDGnYOi/1DbwKZ
lEpTTFvot1JlRmo6AiWmo9iJA98t5FcN99ieB4NYiy1APLvNyAxLHiA6lVG8HeppjJKOLOintf/2
AbdvfcToKu7s0Wht14Av7CnRYV6QlevXNgy182rgRa/G+WhcbXB5IL3kNnN/Ld4A6NFaBM9tH7AW
sdPhYg01sEd5LH7+3p0ppc4Q3RPb5JPXYAzdo9DDfM/xkZuSm9FN4PJKWlZ8FoWdWnuKkQ4AXdYy
WYrz9nx/xzr/cJy1k7uhcwn+WNhDZxCjr58JU9mSLqTJBbg/XtMHfDmJk3zjdYDPxYUaQakk9YYR
aMGaNVBElsOjc7dBy9QjMWEVX7Os+xtjaAqxhO1nfWJaLsvj4SrXQ0E+MXH/DjmtAZog1HZpBu7e
UWbrrzhdp8T0Xcs+mw3hk+ts2h0Nbh/CLbeD/oxJUi1lWmwx5gH2L3jgx9shxU10JfnXQ/HwfsPP
YeN0n8ks8UpI+vHLSZhy2xNzWi0W/w6frOuV8R0CBPKAR8rZec3zh8tVYo4zQQ+FPQSH89bYae4u
USK6JfU34JrH5P67hnTRO/dIRe0gJZLei8LNj80a5lxaVq8R5dPeuLslKo6J5IP7Uc0lAIsCpyBU
iAWv0HbUJepKUadyxh0uoSvyAg/s4dPtuNlr0QijcbivrqhYk4hiME1jEHbEdpGkgBhZ/JRw9/yQ
q/ccGxbotRaa3WVfUtRBEFgrvEMt0AH2JCZcwqOf57pMx34k2k4xO0jLT4rIZEcrELnOD4R1uInp
0P2oihQCWTHcXnWlS8qGEXpJpvLknvzogACje74Ff5Hm/43uU1DvPE0kONnU+9yhNhd722WPwwRD
D4NQ7s5ukuvjxvCbps/3depRqwBA/2UKKIfs0UfQw62HQYSaA6dO4Aa/3f1bP/tRMM4T/xjEy6Vz
+LOg2QRoWI3aSvE96XK0SE9TC3aLRLCsX1NlWmn2Y1ZJlmXqEPlOL4rDy+dHcwp5ACIoivqVwaGy
7R3LmgrwD0QCxC3qSpUpEdR7QorXMk6YEDf4N5nlKR/2lPPc1TZRS+UDFF0dZ1/T/unezRRNQ9RH
zb8KNvQ1vLdtbv9BGmq8Ka2TsuDHGURAv6NZi9usAzgcvUwrsgIzDlSqTQEatNVknQCHU8gzL1SA
ewF/yCWKUEVF99qssGa8arshSYeWdtCJdiOSGYPYbrX7Y1IXb8hWfr2II1MCiwO9YyyeqRroKhKD
uNc5VmFHllMEJ3zUZTX01WIEnQdXfFqoLkW3zatMblGdDSmDG0U9QV4JEKkL4vdfwRY2O/PmEgHG
ePMLYbleadhRPCplEEs4Oyaw39cQzQ0PH8zAXi12Pv1gsZRBceLrJgUwLLR+UyzN7CFLOl+Vj7lf
/oFuiY+GxY3C0tw9LZGmlLd8usmKV+F3z8hjaW9Fwx7KB7zBFmKjxNmySN/3AVEA1UmvHL4ZYq5K
VyVT3mOxTL47V/LBwSka7ljCSeSNrzzbKoMY9F+7qfG9rNLNLE50CkohkxyzATsN7TBjmRgG98Ei
605exQ80wh/zS9pEnAXcjmRok78+KnarhLWsy/5VFaP59zdqdUIMmgOx6ITNdWCQ8mdV+fRTM5D4
R93wxDBdWBBbsArCEP5iEyPjHaZeWVlcz1EsXJf0hD0eXJ2DmaLHO9WQzKzZKxYutE2xQdvctYOK
bZJ3s7ly8HGkhZcEfkUF6W5130rYZQxfaxyptXRuuCYgnU9gSmjnNcwTLlWG5Qxx6N5DHtk9Wtts
krVH6Wkuo3NYDJWeEO+Q7PRTvrHmYyGj1dvItHOe29jBwYefiuIAYKyYp9myCgsK7saeEer9Pa84
HXFIeZYPWtu2MtkMKZiomoBMeG8Qws7xaTL2YGjCNt4KEU0RMXiqbGtEVOP/O9MkIBInKXZQLwm5
t3eVvM/20/YcpegpPbnxg640nJkGju2Aip3fpKJQEJimmOCfyJExRUXiVa1aCT3XgNjp6Uls0nLX
mz/HpF26T3/pbxZFfJT1fQHl4yVqHEgIw0yC4665a8INTIZahE8hnI//b2B5e5Wcs6rkLguIuZJY
Na713199M86n3vO3CFZjCSVkgVDvOdXoQvV5reWw4PmDFY5DeST0HcI1eBWHU92CEhaQVqZJ7mId
Nmcf46CE5pUHIomiKWf5tGNHNoJzdn49yxfnom1iCYJEdNkkYU6zFyUBcDqmYPnH8Hu/rXLSqQOS
EJ4zn1AgpMqLQ4LH0ks/0eZNmSMtiuOaePZ66+LSNvQiooMSJIJK8dIMfbDGoAey8LbUPsSaGE4k
lxVMLMCdT2pjOv5ZDX2VoIEk3UPtAHdYThCu0uoLDwmu1rpNE69V1STnk2PlEhB7zd3AYXkVMVY3
4apaMEbj+hRn7Gg+8W2AP5RTrDH8n7In8OlUNSGRv3PXWUuJeGd0C4vy0RK9a6ZLIhzis+rDz3kk
dpk67INIsUiYp/1FNkrlvd1TDLwXbc+yS538rH3JNZMQjip9M0l3W3a1syIHuZ95H5Qkpo9mkj1c
9+op8RjWJPYHwIvfg4Y+L7LgRPKiQrq4uWOkwCtHs3l1sD7kdF+0lNAb0WxDdS63iArmiLOps1Ya
CijJ4pIYVMqYmjS9x/Jmls6cosAWzdl2Z2LQfMpIItUVGbAhlqsdzLnfcNCetP986VJqa1EdyAmb
N4jDHVyCnfQ/UaLDUsQLI0fAfEukXUWOqGmbmT1VBFQBOsGXhreDvpD46KDm1EeMWFYtQeNfxRMJ
+L8DnbfWXHWrsN+BdJOv4KvCgT3aFvmiHW7zFz/7zkx6rAwAi0ZdXIuOVEvWR5rirNM9YY3SdXUK
uDpXhuTE/TtIeDIGAoKZP/0/N5Vntj7HJNPVwtpPv1cjJD4B9I0W+S+zKxf3iSAERF2HBqKdjrhH
yglJfHv/m2t2lTwh6OWYo2HvtespCvSzsvHj99wVt/kymU1JTxI/m9+/pYX8+Ovzd+Cvy22K2IpH
oa+roLUOEhgCFLibijmMHBC/SkkAHWQTBLrgqhZCTaMWaZmOGiG6xASwnZcnPeZ/E7tEQ3exKIlD
QQb9qq8AZuYY0NBRn0cPwIxUvx9RcQk5TD+nj92gmUHII0jvU9/ytElVMBdNu5oZoVKsITUTfKN8
CrDnhSCH3PkdfCem/6Q+WPjg8e4v9ChQfStskEfxmra/MpqaFl6VUTCfqjK/effYFE/s57xN9v3H
qPPSYEMdpiVobKWZvcP7fap4CJ6YdTBPInlkNAKSMf3Ya6e1FFKclgkUp/VY3Xofo8njt5MiyTmR
hQ5xZpwNpL3a5JaXCmmwsNxRTbhQMfiX1SY8loC6LIy3H46nCcBU4ra4Ki/zsUkw18w/bqheZwvu
lOwj7jHu/JzRxx64RxjqdAzr1fAmd9TCVJsfrMsqS/6JL07WV8Dq4Ftj8hTnyaje3R+gVhBS29r0
aJbfk9jGgHHjm4VW5WcfjsMz7S8DAaXKygjnFn/o19ARFb0pVKc8blWMQ7KqA+y+Yve9l1iP9eRg
ecE9YnnWIBRsHq5u6c9T6U1X2f89PG2nafGL5/jCp/HcrMkY8CMjT0jvzsnUOxoNKGEfmO9LvL2x
XCgtrlBXtPzz1sjqwmQYemGHlOUDZjOP/E/27N1TFIx/gUz7n9ePt5Cz36u1tW+Y0IE8aOibEgSA
jHfyZqIGsZsWUwDMzUNXWAVFrZIt+KLfWdCtdkRXhL5n612mTWMG2bD1oljnjGOF3x/qBoSySdQR
HGyoTfqR5mzQK3H8DA08860z9N7ujh38k54nyD5Sid4w5Q6MKdey9E3VFrg6scyKO4Zjab8rkudd
rm9BtkAOPlnwWEpx0tAUENciilza8BPjeJ/Yf56R0HPkkzBzeOKGWGddgPFhoeMoNOGrMg0XsgTz
EN79lIFGK09Y9DnQ+YgSNnA8fELMUSiCUsri9/Gh4h6bpC3flMJIt5drMltJTL3JzHAivcrpSEk6
koFsSGz41h3NbdcwLy/T5fHU6oech47Nw91I7rVyZro7LzVBX1Oq5wjpVaqJRI9dxo8cPbNwOVJM
44JjaalZAVQ1W5kfZR2TU12xs6W6AP07hyBjRC7OqFa5ayn75wOUSca2MSfcffqSlWC9oFiyO/19
KqQNMmZvQone4Ovf8JQzp/j9GV3sMExLO1tus7igwZRxd8w5oIboqQPUcltXP3d1EipZ+w3dGjAG
+7SHHdzfpuI87zjxykV/PGTrsZqsy2qetTs6d4KLLowhCmHBTwiTKV93mK9OX1VaQTMcUGjfRSEx
X1QIk9G5tuTkBdbD/yRp+tAYaRZWOX7Yo+9VhU/amv65CLNzO97sZu4d31bwdEdSGYl2iGzv2YDO
zjs08r9jAjhsgKrGbzCsQxSuQ1jRU+DrF6M4q4WL7pSFT7h8zDpkhVo8MUuDtpAFI9fY9aWeds7n
Lr/EfWzJNLo2+FQp5zKemyGoxOS5gvh4Of6gn6+fP/o+bWDClFkQ4cCN8j7B+JzAczEV4Ik8i6G2
jRMLc304XiJ5Zy9Hv/rIU7NXhEFq2Ri2eIsIrn6MK0P1Jhfz+Pd3kt81Wu2lMbo1K8p+0prAu/z9
neqQkKf+tHQeCu6OQyMss1e1N3uzsNEyOk+Szkt1BT0LkjQlH4mfuA5mM0axhOkdxPDTKwuepnqO
xaynJI5ah1V6hjHEWAjFFwsyM6tQzpzOGymv5+RimXfIgPtJR7N9p8AhmZLmNMdA4ubd0qzPukom
cvfQVhLTuWOh6myUQHvlTwwVBBdSHvvXsz7PxMAq1eKT1fq+67NNRXPiWkQFf5BLd8wrWv9XjH4E
P2JEgEHT3KtfWuci46wT87IP4yG3W6g6WuVpExTmE1djS0sEBlWQY3nAhC6MG8sOfhZRahnIZ9AE
Pcs4bH2oImfbp6Hkmrt1t0wbvjZgK4ivEIeQm3rKNgylBWjro9LqUTAZ3fYjdmqEDWj6uMW5W3Cy
TBLLAqpj8seuVj4odeTNdzCtRro9Jt5dgOO3w7+FWDVgP0fl2zrPg1ws5XUcOgAYDSoeYuTcvkWC
qWK/OHXZPsYRBfSGMQVTCcGI7FyuRn4PAFmmqQwVlQZGDXk4023v3e/wKXEHMzVjf/GszbkZkv2A
I/984wRXplW3M5RDFkZxA4Fhmf0PYvBieINU1hLbxzBQFFrfY28jdcSyqjs0/CCAyqNTo1n8y/XU
SrKLxyfaxpcNpHp+KyuXXVFvG0WtT+gl05yjT9jsJV9VhI1soXsFUAiVzY325ahbsxEUi1OtCaA2
k3w7xXVKjdTltNcE5DUjknotXNN9pA+OuRCoJ7vVzRBfmsGbQVGG2ZUqJ0qyQIkczk9RF+bKtfoO
KARqWDNX4z/SWocDWZ/b3I6tHXDXc/U+E/voikE051EinfBQin9xp5vawKoRlpX70W0TwE4SXBUk
2dcei+ry20zTbOO78hNDDxx/tfws+IyEa+MMNUcQnB+DFVFcW0mjzAGvMcbEipLH342ut0F73OYu
fr6hp3/grq31yYba7YZcULcgPB0Q/FZDbmGnF/OFnXIeJQgId4FQO6ydp7F39PTiLr6ikjLLv6xf
jQpXw+h6/8hkr4gsgwtzDVxzLI6/26YvXMWHhReAVomHBnqI40JWDu1Y4dg5IB4C3Je1oTJxAm/8
UmgNfzpteijClNPWpeDpJ8AzqVlHxyhXoCwsVv3GcF6e76CIFMGs21634eZ5eUsiwKJxpfRk2m8F
dvwCM7zV1iVxJEMFWhG3IpJm6tMpQObXNAc6kwQT8xjUZGCCBHc4+LT9IY/NjGK8OdhOGBCCaEUU
p7A1ZLv52fhfn7gxMzhryLqXXF1nzIV9xlIUppngxTR7A7FZWrxVshMXgGSi0eIIV9dsjSmh9Lnn
eQoVpZ9KpBkAgqnOBFfn5f37KWr+ex2yRrdN8p2JeHFYIlvOvHCcZIkbmy4HIJxmWTG3TvZjo20K
2hBzGVHKJV87huvsYKOw4O9/aPL9qrLXCfaIHQ4jSVF8L+OA4hIet415Kjd5MMgtTmV87M8uGtyp
jBX2CvyLl820pk8p4wK2S60VCcDrtqJXja8mcy42OQaobXqtfsrFluu1yl0oIPPyZZ+Vo8Ngeyge
TTisNms+Ac6cTvKpRHdAmKmd2BMmjnQi7AbeehU6Zh/OBAUc/gLHp+U1eytGDCkAivd/DPuRJzf8
uv2CUVnhOtTD2Nzsc5fnZSqeUkX9mS2zomYjerimBG5aiEW/AIzp2IG3ahCqFk/86F3TxoJpLe70
CNP4ZaQPiYU3PiWkzZVbG0lOMyLTFGLcAqPj98KVlaVF2k3qmOZ+eBkMkrRfWqr+LQWK8K3bMUiI
w0gGJjnJmpLJHvm471tqKYUNQF5ugiByEMsPz2Zi1zvckzzcmTrm+xkdJ6NcBqEZ56xLsNhq/zUh
Gfmjsk0dCEqk3tXL/6FR7oiG9sOpcsCp1axOJrCDq5d81zCe4Y07BzBJ8/C9eBQ3dsLr5y7cnm9Y
G3fP8ZpQbPVSZtI8m6XIcWgS5+vtQ3/FxsEI9KsBAKodXeCTW+gA7SQ1vYw9xQ6+m03IbyzJAngs
E/MtLpoXdbfpGWBtp3JlG+7jAtcmpaZ+JWXP5TMezUfMZg+qnnE8d6iCnIphloJpFyaidJD7slCj
UjLd/j5njAW4DvrLrIqFwhw5+YGG2mua32TZbXkRE8pE9LnHxuM4577EGCHGMSofkTP7pQ4tn2YT
MIuvQaoekc4KklwUxrkAzXX1jEgDEcGPESDjMQfM8kO6uFnkEYrHnBVfzcT03rdbiOf04BpfGz7w
SWnLy87lOHIl0mpwKq+jpA1cjHWW/yPR0mzeeuQM2BFiGlJ/6jn15WOeXPvtAf3fP3Y0WBw7EQdW
yo1G6BRSgHig+u4JU8uX0hWv5tw15w99yQjCurQKuGD6ztS3Ei13FcPEMxSzkFI4BhsqRtH1wFU+
KOfEWQJg6BvWddRx2yPh/IUoqujtDpKHVLl622WLEPhWMQOaCUeGawYSEorGxJO5r41SgLynEbuK
1lnVbN7T/4Dtbz7e9M8e+gtwigxC2hI5+SZV6Kvxs0rLwOoFz45R1bHnJsA0PnNfYheQ1xvQJqbV
++2HupUoDiwjnUEvIcs1CGE2xVqoi/ivYkTmTafWxDSMMK5jTxLnenlNDPkYXlsG7hvMsWUs0JiJ
K11xmk7k3qYdEzw76HnOpAhQejBYx9XFExTD3V22IuEbbDNBAyJyeiw3V+/tdCHG+QEm0DG70Rd6
FZICYmkT7UbVCqDSz5yPFLhicNXysCg9G+My/+4qfm2xsdlXXMtyUTFX2ol5QGFt9Wyt1EoqKYJR
xgnuqRb1W+ZSTJLeedpIh3QmscoUWd7swJylFVfm1D6poBlurvsA0NmFP2tDwQKxkz+zTmr/K3JD
J6FuErNjif/J3DcVkGV/yocyVtECgIPtd3syBlChvsYyDtWEJT5lE6hD3bXHNDKPECJgRzDyrFD1
bGdiZNYFXSM9EOQS1piQrT+X9ABM7ZcABW1pWIcPN1Nu9f9qPNJoty48FkPRydyswSZo5VHexoN1
/gcfFmNaxpO+Wdl/CoA8bQ9j8B6kv+4pqSe+ViM+Hhz6NNtb2l1wZukbqJrvNYiuIsb9h6uPlvnG
Abm+b3x1FGage9MFiCxSAUpOq3d/yUaNKZPx5WygDRZRp6reQMQQNAcqaDCzapHSfIDhnm7uwXFf
e+toSTl1qXjWaRBTE0D/ByH+CbCkWziBxi9238dFoeaQwkQWmYR18A4Ovd68VRC1qE1XD3S7vuXJ
NqOf+nGUxuHGvoFi+8Brq2zqxJi74vvJBsUyHMJ4KHd/fTNrixc6wrxt1/tGfbKZdjXMx8upK6m4
VQUP3xujOFXwwSldEbLlboGNQlI1+Q9DKNjaNQ7HY5nwCz7/LweoDlG5J0pn6J5J2wIIHkgF+o19
VrIK/1o7Z7uI03JOIqO4BGAS05nPkMZEaEqusUJeJ5FcyX+oPJm2F/AnxQZT2cKXCRRI3Gzuc3Xs
skxZEOcGPDBSGHrEETFVkXOFfUDDGjcxpyXExX/rtXVBdwZZq/SV7pgK1X+P2AK+29j0LH8L1cxh
HRDhvU6h5BcsVVzErA8uahHXseelh45E1Qnr6sP5z3o0YRiaOMRqjTfaUcqKJLE7YlSdexOLOsHv
CSwqX0ueNEblMddXGf4aGXcXCNSZsoBnGRK+GdBUbDD/P8IRnVPR3ViX3KKxaw7JByfcqJyfNtJ/
i29QrucwTwRe+Ppz334i/QKTI6E8Q8ps8NUQRKBIJlNF9/UX0xE5M8mHY81yjzWBhUQ/jR3OLHUd
ynNiuHwwAA+Rpqg49WyibSD4YzoNbgnvYI2vxsSHQdiZJTvo2RgDenNYwSB8p25XCRnsQkLZxpfh
TXipk3Jq7c2cSI0jZaps8ZYTgLRC0ej7XDUuW4b3C8bGfhzWaPmd0kzwQJnD50QptklOL53/qc5s
bWXgvH1pptcHWvPbah2qLb0aYpFrmCrvZFrykHKwKXZlSfxHj7SIDZ9nwY6CkiFxHIVF1bXVdq47
U+te7q4OaHVubJD2AWgAbO2Q5G0fwU5sHkQKF8o6H0kH+Y2EU03+WBz0WNxzF6EagQgcMDwkmlXq
nNI9hAcVakCAm8gDR/SCuHqb5k7mn9YdowZaDTNkdcfAoLVJSZrl0LoMxh3yJvOlXRsUM+DBYSts
m9s6nz9XHK3ljWZPwSkWEgXdRFSOm4UEKPX3CZf7kH5ATChici9SZ7fruSXCsHaiEE2XPPm2SoNO
BZNMAtwn4HKUaG4pW2/RCJs+I8Bt3Ruo2epT5E3r8Wljhvt7Bwv8DRKNC9xksN5VMEMz7FsO6kqq
ROzXT4e9L+IlaNBFGCclZOF7X+ptH5mCEb756uoM/gl3QQSK8iZHvx4biP0+g8leU+RVbBRvconQ
9a/nKvpgYM+WASumkJmjEIKYQhDEiA4YsSh9m4amtpZRufsLQrzjzQQrS7VjOh/AdDW96NZj0y0B
4YJZeyKixWaW4DpVqg6PcJTGZi2zka4co00k3vMz1btXwAKBq7Pwx55m8T2o7uKnzRz0YihY240b
G2yzOnfwboY6IdMcjj8Or8CcAXlQ/FfFP2f/DRqFEJ5tXLd74GUJaUeu9GVmwfOS9EdesgATsj2J
ABmfqdzBBuCU3Sq6TpbS1UJDSXqWbTMG2wvIL9Gx2LT9vq3y4ZY24qzuqwoGC8efoArruTCCLyPe
1jwwjXbwKsj+5NQ9hmThPiXoruOKscoub8BFWF35uEfy7wfQjGr8O9tZNRDSx7F5iTMj6XqP/aNp
RJMpa2FjZq2OjBBFHfqrue8cpvqQbOh1nZcDS8pP6KPGacjEjN3YbLBC+90d8/qXVXAX5eLRPlSE
7/u7x+rw42UW519QlLfT3YCDX7tOuav4OnSD7F+pKodq8R+9+s+vfP4RVOFbq4+nMoeXtl5QohXd
YW1gSgXIuk4M8a9ha/EGVj1zzbCaKepi4KIopBtcLjM4qr7nelOvYHlcxXCrX5lXmPcpSKKSV4No
hzY2z1qAlrwaduVnnJW1yXuFFn5Yw+KCepH4qkTgxf47epM9yDgiH5at4RKE6WBOSLXcbFR2VhYL
+hoGdFyjMTpHwlxskuUP9VMqdSYy8tJym8NaUxQB2sQDeNrZlwLc7yNjY+STlI+SiJy1dIfk6jmI
f8kmlfnkedr3/hYbvW26MLwzDeXIzCpkxbIKqt6PPCo3Roo65R/uVYw51GPZawsyvHStAj5Eq5/W
Ja/zefiGURXPaDZA49B7YwuXgnu+QoLHyM065QtuW1UZvEGlze9IIaE2wPBnS2RejKSLNGYkHEPP
4gKjsKMwYAZdC6Puj2nUSwbdAZLp9o0gxCEpmVmPbKznhiwye6H1K3Gx4nXBjQUPe9s0GJbuzhCT
Jg/pDoX3AC4BITWjJbhNmM60oV4/Qx3Odrma6TP8GCpGfpA6y3mwdElNUuFcy6PV+dkBUGT+s+CT
apwzXiiaW4AmZB5h7cbLAv1DlOw3QgeZEegh2Czc8W//oyD5CMh8sv4zXXd9NbbnPLOOfCfCCY93
1w7ktJtkTa+wBxMhVqcOV1IuII8e39pJJqi1R4Fv7LbZBYxs7E/Xkx5KX+JralTwCR6m1F8rzOQG
KbEptUD7IBz5gB2UE2rjkyOEYmuBPmDoHbIGN9BbFzr58apj8M2T+Sh29anmi2zkL3rxqFl0fTkI
yVgSLgL8jvgMKcDUWrIO0KDKQfyqFbeXnrH4XvYkhi4O5EUl6TbIyI3iB4j7fjWBkfkh5gR5ThC1
Y0yd78oYVDyU8TwrJjOpMdAPJybaTxkh2cFaubXYK15mIY45xMnnArxOVPYBK/XZdmRZaHO0BboG
KWCtLSq/MkOTkzsCZPfWhgOri5q8yj4I4ISECoU7V3CxXVo2f28wxsyEBRMbKJelzbs9LQFBFghr
CEIQZHCfbTgYUo6ppOorM1dvBUlEDmsjdjocxZil972oGCA2EooFWPMO35xsYX2fR3sD4GY7L2aN
knybwMrDCGJAnoUc23isogXgi4/yu4GIqrmTNaKJv7pOWdPi0KyR0eberNvqhENVOeADMskA0F2b
6n68DqLWc2orp9jH18hEfS8BDuA1WyyOKZXoF5dYOBoFNiIHvgupp/4HSM0veKSyt6TCGgZCWY9O
v6fdznpTcb6nNYgCJ1rvkr0rHt2ulFk5TG0yhxbFfYTYhiVdN4qKcYcb2pp4+I/g47NeW1oY80eS
LY+PXfuLapQXCO1ykAcjjPkE/TR54c0p2VjJzbjKlBLMtflSwC7rKVHnGQDmYpY5UbQtYgPsul5n
Bpt3rqN0wQVNwod1HjdKle7X0EE/fFup6dRk3JiILwAoLknkx2ch7tu4j8BXuDriQcErD9v9KhB0
E1ERnIREZ+lbbi8PqHZzW8QoCQPkn3O4UsT8eQScgdkraJZXNs4atTSLr3Atn66vShGqMWI8C5HS
dURO2nm0JHd+0HtwLOCeGR02ndhW5upPIeDih9d2HoWQ/5Yjigp/uuoHwJ5VTRzs0s/jQFljausD
j3I+PiZ1+6Z8zMAh4pmo2sPVzVY9RSeZ9Hxvs7F/ZB3EEL6teTl6oHKik0pSHBQPK58itH16c3ju
a+5YMXZskWFxBSUIIvcug+QGY4LBI3cC7E5Rrl8TZanDI1CdXqqT1QOeYpN7sn0iNk0YhFUO5tzC
Npj7Pogq3iCS4QyZNkmjD1RHes3DCQktKeFxK/RbMGwSwd1lGi6fCCibGGXEUgav70JV1MMdisdb
kFaS866xCEnpczRCxqN57fKQr1zVFDixteIfmVL73KhPll++gdqRGahiAsjIXWFOAvt4fUhI4B2G
8M7ljgYagnaP3/z1HcH2dt36ZSqYEQR1mv7Di11sD9GbS3Jm2ffm5S7dRIeiVqA8n3/0+Qbfrw3J
4U7Fq0r5n86KOwahI+9Ktx1hMVF3K87+EsId2H/MkHG+NP/WkuJfvvArmDd9cs/ML1nNjyRTbNF3
RQYm9OE/sasJBvbT2fkushklSmkZL7B3HOfTSMz/EBWw+umI7+8Q49AKaYm1vflkV5OSsPO7U8sI
eR4F+KvjB6Pt3KLToIVdW4dbKma+KQSoIEyM8hoCghagvxtWacdFSj6tsVmqWGXT3PAk+wbWbSaV
84uqRQ2zbgaVc/jJQTYPBzQ1MTSRecsuWzGcuKJEghoNkeGvxuzEGBv0q04F8ySOBJLJc+6vm3f3
mL3MoF0Q720OFMEAIQCecNpXeR5vvSOnyn4Hy0SWbY717Z+S9VzqqAid39HfgXbzHd/rhT+kBcX6
qfALtJ0KBymlcDe7FzD1YOWJzm5wAsC3mmFYGmvCsA1+Fin/QK12624k6kCzrTRdHY8xZEDj1ADs
Hl4H8ALMibyvEMbao2h0JbHIdRatv2ieHAUxjLe2H/aR/Efpx9CrLEMTIrD5BV+K6UHihJMvaUb5
QZZdu0DsoEywSps4XEs2ajMqw7vfE54GdjbH/oj/dW9aKD0uYIc48UYEJmT0BwMWy4xdFgQ/x85c
agOoecTyUz5L0r6JeMzWdd97PoIaLtqz/HluPFFIeywZEhqYN/gjifKQ7yo+G1P7E3lP+R3fMlUO
FDnD6W6oFLe4B6aTFrx4nn+WtUum3AmnOUByx8iMAu+hDrott+0df1TVw+3Ytu7z94XB8xIw6FgU
UKKYY+Bg8XOO9CQ9/rGcc1APWUH0U5K17DrUKhCSpRXOqQ+1Z44aDQyOQKdBPUZ+nZEkFoCAmWkz
vvKmN+F1m+0VjAxIP7CIm5XO6K/OhtZljRZEpduGkPB38KFbhtjOp5Y+w6d5Tx6SuHsXAsa2l62i
/jpzaAoU6Gn80dRH3ayY2RGxzMIVw3M+JJByaHI8y4BAcyFltdHq4QgH7OLWpPh3EERa4iXNaewK
GxYAyrE0lAW+mTl4EhecqfqP6N99PpfpSNzmXJ26ak2l+QTxKqnVjFrFg3w7EX7nzwTZosDfsJsD
m+Gh67tEnhvSoatMk58cjiLxj+7F9BSiiqNRDCmqN0bxdNIw1OkKRjbZZbP+RbtfMtHsuiuI/2vB
gXmRn3OPK2kIjxWyC1rrrETOF5AK0xkZSQZDkXWVDyDl6pxtgz3beOKUwAmOJYNLOkWeNqwlqcti
UKNnCLFoVbyGxZX3eCVstfmwLr8CRrap/rGbKveLZ4rUGtm9qNzN9GluGawZ4vKKwjO2iS7X0lr5
Cpsleuz/sLEz5nZ2+Z59JnU5PprcJBfm70fCxhDxdI8DbY+n8DGcJXqVJu8iaKajXc5VWQwMWaTv
f+JQuiWFlY5tidppnYL/ee4+k4IgT8ifLy2Ld4ouaX5EBh/UinPtqv925F17xojdQs9x7b88UQsj
Cz7q3h6i2fBDRKqtHFp9+hBZyQzsIP35Um7r12BGZ0TT7tDbdolh8ZAdst3G3TcFA8Lu65+8oXY/
NIY0rEvBOBG+mhN2QyA4C/8UNx+1UJMIR7XxmRrRemt2snGq8KtmvsOwnKj2z+qXfmZstWNjc5bM
860pdymoFRxDf5unBlfQQk4+iJ2Qxo1kOFGZsJb+znA6aziZK/GUxEzadSmZfr5O4aYpWNJlcUnR
fCHnS6Z5z50wljXuIT8VSHoP002Zn5MjevzuUZ9twYhx5hs5FCCE8BOUi2jrlDeMNmeWBBsdxIck
6QuWqIpEoCGP1+hpKpCRygartqWFkis1kuGJe9FRDqN8fkWcPP+uk/TLRa1R/WRNdrS5AwH94F/k
74LdWcIFydkB1ufDLnOifmQUX3/eIs/gjBzlnTMBjrgSvFlnlsv/EGB0wEZA3m8AYUN4NPWKEDU3
EJPeG1gM3OcD2DG5AvMSSeBl/qRzObY619NWlqISE75gQ7F5b4n8pK0yFieYajPMwG7pSEQW0xqd
dv0+pe4mcp7uJONlz3PLXOXjzOCUpky+SS8vCw5kcUWmVa43JVgl27FjyHmMpa/+6RXooGDcRGOX
1tW+mz4ngzOMFHGnvNlD/673BlEDELLQLiIb/YY2KmWOLqaCz5cceAIMqR9l4i4bgX5/aKK7jLDk
52Qv+2k1DpVryhInbOxuRX+rv3FCqfxKOy1cq8jZi/Z4UDHBoJ0FUyqXIfCChaI5UJyeiADzu1ei
W4WBwaqDDm0qndrFokhq5lDn33nZ5/k+biO7t0ppxWuTiSXBqXZmVsKb7ABRBCqGch/Bdloy/pkS
ZGp/H1+pHQhPoRY2kCbPqPujCCORGXildBkgbeFBfcj1rir/HO/X24obxnXwNdDuM6Yxm8UAvjwa
IAvqaba10z7Ixikgk/iSp7OFtIfCLwXzFKY6R3LPTkbbkdkxE+jWoPJHMYLMVpS3zrVnXf7UwwuD
VjsxcN72b9sTdgqkAmsMswPnisOwxIMIvvNDq9WDlbGCR9PkM6V8eAMqS4rV54DuWx/wMlf3gsSc
wRkSnh63jCLuGQvKl8tocVJPs0+dmZ8ti1x5WOHPNNM+ymB+ZDqzsrJbx1YQ1BjKpp6KAL3FbvnF
7Sl53xavBMgC0/GxMcn/eUjJ929TuieGTE9FojMNzTO2Pn8by5PdU7KEedJZXl0dF07GuymPy70Z
npNdllboVLqe/+bN53ZnQL5JAgTViIX1bZWYnPpd++au3E73Nq2vApn8htgDPIzatHmm/ux1yc7d
0a9oNAor8X3Y8w1X2F8lS3aylJ4MDmc2ZMs5bM6s8fzCgbAp2dibdZxbdq9NtvrVotq44dhOvXTT
J5rSUmqN9k3/mu48ndqb3+9cK+780tv+HceUkabVXGlCBtFEHUyOtZ2BJk2Nd82FDLxQzpbh3c7H
QsKew0eVYUn8KDpH7Z2M2BLVbu42HDtn+95jObntXJU81ovWbwjHt+ar2EVEnaHP2fgaftX+Dbq7
8lEFYn6I3iPeGKtIJkvmSnVBZk7QVLNfITllLZWvZL++w9qix0yP4SyY58FTotY9/Rp56dJfbhuM
chX1oq9nJgc/EqBWfXBKmmYxEv4r5+l7rBHWnJTvXVW6dGUCOc911/AIIuvHMIIHRlqF/h/KEpQF
JWmfrJRA813J9JqQH3WiaHu46NRI0aGBsQEtkTc0Z66sajgiY4JVRQ1GNFazt0dla35PWJK/uKxM
j6bNTTHv9+Mbbb4ZUANAerAsYYvI/i8mA5n0ptkEbJnv5jY8F1yUcE8Z4NVymqzcS6euLoLjvS7C
4GDDY4HbZpVK+xhZRvaM8rNoaSofHXU3viBSDvAmMXSNQTQsOKHbly33NIJq/57wXTWzMAi72DXv
p9rdITJaBEUWnC8PA1Pll3co0aEuygW/OvgBgP6U5wGmgq2917k8CjWr6AfA1WbyTJERnykyZBaf
4KN67Ofox43eKy1EiJgGtDUHUVRU8Qvc5dh/Y9l1p7taIdiZ3SZfYQaAfZd5UKvdewYIj6C1JwrS
NbXrOM0lINF1ByoFRjhlI/MNPu08bIl0834hbPSXJuUed6HxrBbBCuCnN+l3Qq6gW3Boc3PhHZCe
MOEujt5+Q1hSkqASRA7ASt/WJErYymk4B2YcaGq6lQf2bkrPOzVYQe1wi+jAqaLVCwIlDDLflW0f
P+QfpkD8fl0BpO79ssmvp9o8/p0XfEijiGxAw6qx8NkBfEPKWBQmyL/l8YMA/AM0CjlGslQeWbhr
8X4Zm/geG7PpKPlr73dcA6ThQ6buTdRPhREzh61+msGvNMqegqClxMQGk1hsdRm6E8j+0Y3Rzvam
9UApjtYIZKvD3Xzsqj2gVKcsCSbhpgkPGLLMX7SwZKZc4UXcXkcl3BgEplRTQZfTomZ+6EWYOZi4
2hp+d/9c1q8MbuUvEw3EPYiY7XOLSCXlBGXaas6vatWvltGoJzqnc10KtpztrDYqP1kf8E69Mb4D
24EPvXK7UyXOOMfIvnfN30w5kkVB4Dh8A0Cw9vI5YKK3BRVZ2lyBWIgZHLqtY746nN5OFv/lzyri
Dbo8Hbn+QkbnT5JWew4GCcWh2c7WEXR45zhEMsf/wuMd5Ub53irLbGJM+iYqtY2Isj+6gReNmJbG
iuzupMEL43TaV3xDReV/kAwxOHo1NYUnz/vUh7V1bucI1qELI9zhaWdSTL+t4AmLOhbtxBDnh3z4
Rukg7Rsb1klmgf5ajQ6Dbs42HkepVzigXggLTnrda0AD531IuW7QNe+iRk2TQONuepnCycfASO73
O0FBbOSoCZkZC1BIA76K5jCuD2zfInWmwffRoLIGkR5OOFiG0X/xkl8kjI420hsIKMYYWcWxouFS
iCuM+CfYEoQIDGwwfQuSTCPVujBiTs9w5UoDA+a4u3Q4B5vFpDqVhfbSwvMrGeun/6p9ZzTKcwUr
hqI+ixR+GDOOvZwCP0tpTYARpiHjsPYRQvjHix1o2+kfUFeSku3ymIHZ0MbvjmCgeBjBBO3amzF7
M4AKF9OesYgvfKBj8r61X+ATO+MlUgpQe5ltVChrHLDEm2UcJZAOiY4tYOak6IIsMLpSnTaMmovW
RiIZQQnf/JuQg/Cb+lmRvfUYrsS+FM6hSiUjxp5rpjYXKmAJ3DocXquiq4euhPpARg0YLk1N/+lc
tqCfxJ+cYk/xHyIvnFvpzZamQHU34qrrlQp6otjBEMfvImHpIVYfyWl1qIEMOZKrVzWhrz1S2U6Q
ymlt/DP4dtR5vniQ9xUXuxwmzVopbHBF9TaWD11LGgTaLnGAi7ZDIt2YGJVbY4k9MTMRxl/vbq8x
Cc7McEunBF5J9C9Mcf8R+7/FD39TUtY8oNxRtxvKORcOmlvlKv+BJWQgA/chWkae5aj2VFVt7clB
zD6GdPDJGsStRWgUR5w/8K40fLbk4NEM63FCIn2oGUtC1r9GzgOEs9YSZ7A9pOmYwJS9OKJydicF
thAOnYFdxhSdYktxjLYaHs4WVNNVn0PgzRnF5jqHas6Jfcfo9cPZtyKFkJf3oSQyqZgo0Qd3+NT9
BxvhMubcx+GQd83UF0+GmM8aRSgGus34OeAy1bOFkuEIk2RvDTiSsMgzY8gu2FJjBGbckjz1QREw
Y1bHUW3xbKXtJyCb20JAtmLH4kGgmTpidcrN/kngkOkcikwi/wE/oIFdZN1+aZlhRA66PGxO+qFM
DIWGbg8NIXgNO/wz6VLhYWewbc8hu6Bp0BDZUdPufFbtmCCO8+Pj4EXoaeSj2ZplvkOwHakaaR1K
GhpOB18XCyS6NAdRoQNfiiedhjV0+W8lu6tbFzxjyanwtEXkHD9mZC+mOv+yT7bs+viclotgcvVF
eHSh8VZLPJ9isb5OzRxLnSlN1rNFomLPhFWhF6rFm8ZTmS0+CIAm2TAjFt1ocex3Tz7DlTYVgMYU
SQye0yk3tnXU0X30tEJeGhpcjZ7IWTFJvB/k8D60z63if/Ymi9WHoEJr1lQVvDa0tN8SPLH+m5Ai
x234vEcvdQgbiar6m45kVZmPFwmeosc9raES4pUYN3qhSASzWk/3Tei4GomQggPLIFou/gAfZfHF
O19dW4vtBaqLcxIL6JJ64IAZ2wu73NBBMXgWgpkYFm0RdJxwRgl8UANL7RmQwnnTmXXDXk00pxvd
5KrAeu2iikg7Ig/b2pQU+K/LKYR7/SevYqZH9BvFt4MKeCkP60yHzbJS4ZkVNlpGYvec6Cx1xCXW
d0KQM2Oreq2SSKaAraFXaHPoSXGQzBctAqem6XefUKlanKeavqbsftNkIgWjLPBsMpFyJeEitSJJ
afSFhGTn59DRIxDz9IumiEkkQAnOsn7q8zztWsScrkzLEJMdNVH6XYihI4st5GZfa4eaLkBzEaEc
tutHYJlrvGRSqcyjPEWMESn2yVuzM+ZOG6rmrdt4OKgfxRvRmky/7EuhGrQkb/7G/94ck4+nVO69
EG7Fj/vRYNgULhLlQppGnA8EiUwZXuRm4snWYuNSsmrcmfFDcY3+Z0xQMDgcDr1dOLKDmD2I+kco
kMA+Q/8yiSQ2GnbLMbwy6RHwPAGq2KRKPsnBKZAtwSulMRxNhJ61MU2KNh3NUvamLe/1IMF7JVRe
xFcIbztEX8UQkgWB+Ndur+KtOldzAhEIK7tadOUHUKou52NUpuT8LgkbNIOWUGD6EToilLw65bQ3
NJAa5QyUyC+5g2p9WHZsC/UCWSZJatu1oMPlqfo2EftghM+KjEINamrED7oCyZIW0x9jR/vl9wIf
bAirdXAkN7iDvO4W+uWcBKi5cCCDu91eZeePDgqVPTK8n9AQaywLHj/6lkvGeVzBZRNvLdrHem8j
mNaHKeu61dBgfc03Beb1jrGOthH+Fy6IOq8IjllXsxAZ/3iwcJHqBXjDrrzhayvdzeYeR79vHRT/
Sl+FWUtvGTjCNGQDKjwGk4pxhgaz0OptfFmiLdHtl7y5bcLCRYpn03dfUTUi9gsbKf5hISqYTMxg
ej4rlV+hjtpqXpWFJYg2gJ9kRr8RiNFufQBMNAi6V53YsS7LRnTmGcLDUbhhGjC0i5GjHNBjQHIl
HVVZe/Z1cpVbFqygQb2N8WLKBNz77Hh1PCbvtBH++ygYhfEjCzRjZbIOqWehpltYtNETU+zuVDUY
XR7tq4/tMrqGe6iciZsq7frHYXmZqrD0DTmwVHdfodlttI8p9mZ/lpdfMGLnd65ENnASVHCPzQXl
Da36AxmC5YXJOE134do5rsAWdljcNB60F5ypDfT6CcMt9wbY8GxlcfysAk3dtlZK5qHnmlgN/fpS
3Nlt9B7oWnX1BeaAVb4pLewqtLelS5KIbZUaiGKPflg1i+o2KE3a0oueEtKNTFihPc8BNsjJSHge
AZ4hh870CJbVRv+7ODCtLuwJQpoZAEyfgpUwHPbnbXjR/sKk7j/hPXEzcGp2CJccBzCRsQigDgDR
PCEnVZC+SDP/3KOScw+xPKzLnWGk7Lio4Xdyx/Abggh85gCi7bqDG4v0xK47wvfDfeDb03Gt0zPq
z+2efs7Hspug8VaHjsNKU7Eu14QEYX4rY1S7ps7mFp1mwCgSwMs75v0m0LRgAhzHr/+CNeanExcT
8eKZdViZfhF4K3HgJA5sotarLjPxOwo34M0ngdZjOiSSrtHnciPFMO5BpvfUF5dUoEJ3AzQn+siv
UilC9rnXqFcEQ3jGGEg9clVlsorYsoPi/uTk+jQLz4t7BVsVv7XyRAKAXsIfFVaCC2xzESdfvc1a
4xtfh5zNVQYkLWo3R1+vSrTfdGpwCBSIkGJf/llUs4F/XwFZpwevcX5i7a9BziRjvUjbGorOiKCb
8NvLQb12uhV0ClCrHdVI5jQCrIcDm/eSH2VnZQOk2naaYkGhRj21humL6KWDj6zoRdVgssG99pFA
2SEa6vPMFxZkTFkzKj8UZcDVy7PweGhaDhIRIvLcGQ61Tm4YVBCNSuISPeqHv7TYipjjPz5p2E+a
8iJQQvMpJsUh0Bd2JsSSwjauhopWupAvJ+G4p3kTnu361T1M1zAE70P+e7mVBG9DEHGho801BpBJ
hxeT11ULiFHQ9Jo0T4mZdUdkRZRaZ6xsNNan213xDackuDO2NwOlpDZyGLngYgMYQNUIlZJ+utlE
gZpY+k5FC8av8CF6mc1W9adfgjXqsnoFV28yylB7AbExfbpSvANsKeQYUTaWdMivC4qrh0vadhWl
mEGhLowHgb/6gGaUpoq+urzJ6exivGzfjAM04fiC6bhy37JTNDHWf8q5kdCSpRB7LDzduSMZzzU8
MCmQMv4XGlGXlPI2CrE+NQCdPaJt9O1yYJC+aeHm4mCNsyTL8J2WsHaMDLWK2PQbVKy/FvTFwzsL
DA4yYUcdQAUk/5jB4xmTklPAcO2QpO/ZzSDZy+Vk0BKq9aRrj1L2qzvgOFc8nn2jBvCHrfovmMFv
7NuYzNySSZkhjAlDEZ4NrAiMx90scDybcKc9IJn72Ihi8Y3GBHaYQJ2M2Hg2hXhx9T3tum01vNB7
J1dT4ZSNgv3cqNaIiDCWaXWxn2VG6CqZ4cdrydsrY2FTpNTIGrsS02/0HzpD9RkiQ8ZzwTtGQeyt
CEIqlGUPwoG7DvT4F46b2no49neU76Nmsw0lhdCpZqiLCNJmtJaF4yr1YSNHzNZ/e+d+qETiGg8D
abuaQaNncWrs7A3gRRZGFIN3QXh/U+PbOTMTVfljSN/o0h5DxJUPFwhOZvV/s3NPdoZLJSGx4vQc
FdB5LSZUqwoKO49WcChKO1oBogldK5SEfy4QeSVaI97GyRSOsoxNZIZYNL8jRz3WwIIOZOrBRAre
vInWVNFsgg53NIE94gWB2ACV+N/8uuNKL4lrKIICiG8fnXpPErZraJl1OmC9Gyzvp1QJx3m3V3JD
25wtsMDCgSgyyDk55mGE5SCbcGuN/gZv4giAbDIKPbIsmp9C15uBpXumMr+Q4FOU4yWeLq9NA7Ei
JFNqD3wyQDsydDNCnqxkkahlHdoJUKr/2kUYduu6GlbJiHXmzL0a8UHIYLmLbNmX+wg4ywZLygHz
ydxdZzapLEZQ5JT68D/q2XbumKrAubChS9eJFGh1N3K4F+N37LsROZU2vTSo8HJE0pMOG8yRupmy
Fo7PA4ZdHUXRp651PG9NBOPiXrCuJEsH96qkfF61VXfV4VnwwI9T0rJkxBKo4NymXVZrfBeVzUFR
MQzGPsrYPx3tmo8xetYyCjjglrDfzJmnNPiT53rz16JOlBfFamCjHiyv4swtGiz5pDCfu5+lUn3I
7PEnn6kxYXcxcI2XMEntWShfoUwvzOg8PE4x6Eeve7oF44cTfWOcbollZtntihGKS/NPYQ90DK3h
yOdPEqgMjnAGUGwW4+gvOjLqMmVjR97tYCrx1cMBm6c8N/GIUwTdi3XEnRHJkGXWQJQfuiwexuA9
RdvXzhLOf4Y1gBvkRIqdKMD/lC/eUIhF54t0vfLwlEJtMIP8gM9CJrU6fv3Q+T5b0PQ8XkWLDrae
B/R30is3sVOR1yrnw7Go42owngHwoSJmcT8IkHRSvYhD0ohHMrrZRrFBtn6YXYgTJ7J52DtaP+ww
rXAmDmVFGyomYZjIhdFPKkyJPefrYiFN/SFFN6fNRBfiQitNS3etYLh7n+vNIYWUw6OkZA3KRLYc
bTIhYMaXgSHCOLGc1hKh0cRQE8KOqVN13Ej/hKOR55VKFohCzj1AY312wnA3Aw9aBT22q+57130P
BuX9u1oBP5WpGKmrx9UWqg2Xv76M9gi0XFzTpUPSDSgJakpUkttWNWDCwOjU5uEQHafcM8oGEpIy
U0zIEiBvZyPJ5OKpT94ttGynOp0ztdM7hm6MoKE+Gwn/lX4fb79sCiZWkhIRY/eKtb0c2yOZTfkq
2kzrMT9L6Ro5Sbu/mJvDtTAlpzJdeZeuX01L6tg507bnaCA+xYYaUuyUEJi0RQ7vKxXZ+ZZp6HaU
kSs6Q7LyNCcvuwqpj4NARhEWqICaDXlssSnyZTPAqO9WEyoGQYxw0iOpZrLlP3TabPdez3zbXcs9
wimWfjToFzKzqvH6ejCATaIFTloWCdqk6cuhyZwBgMDK6otFHUW/B9vMZFtPt4GVoo8y43gm2UNV
1Str61dYQO18r8jxBxJswo+MG59ooyiKlTTm4plYeFzPKZH+jVR3a2IEpkjmcg6hthR8KopngptY
x0PFau8e9cuqZFrmUgUVZLjdaKK/fKbbrCR94fuVsXBnQjiZRUqKagfxrFMzF52Yo2v1Qn/f6JG7
iDKszvbi4Sl657yR2Bnt7tmguBeXNJ/OULjvJtMWAiQL2mB7pBnn71qDF/pcpdFamwkAbjlMie5N
iM3bn3kuoFKl2r9VZ7WpiGVgF+EEZgm0p0Bo/WQ1LdMZbKQh0Cq892OXGzPsXAu9bFMIH9KcdaQ/
SisljjfTU7Ta+og4E9Gp/AnEOXJs3hNHPTiVGlfadc2hqbRnWE7JrYyr12yLbckeaP9HykrbHRL4
UFYuBfpSCMp5sa/frjUAEuPpCbzM0nBJ8NFWqyxNnoajEMYE6H+k7GER1xBBgOyyb4Lp+J4aqOuX
d5xjvlCxQCAcm8cZIRYaFbZdf/5okXnGe177o2Sdl/N1zXrW1NQfMU2EL9AlNqVtpUmwaq/GD8BD
H6RJ/oHC3kSlE11tH6nZKN7WHYV9tntAt4SyDacCTdEJOMFIwC1S1fSwDow4G+OFZkZxXKFwbg8H
kmj+pIGbMvZNroNnMKrTeEpEPhzRvJdpc9wiReNAXHA+JciYY3jlRlqYly+lD1LgTsXwXYBpcFJm
vGn8wuajKsZJNKuFxRXcqGZtFNtXu/bDLgjlwA1zN+5QlyShvFddRO62nngur/Djw/Nz7Ifr7otr
LVyr0BxNyds9Iq90b2Doa2jBLYAu08OkBWDbSJid0Lcpn4tmWl19wa0fh2V/k4GOyXfyPfvthb/I
PTtSpNiwbvHrCCe2YiYrL0SLrnC4+0rXZm1LR0R1lCDJenTCKT4DndU3Ug9wdfH08VQjMydqPd1d
eB0qBo6q9RE62ZZ6hzVol4jMo2kHyCJOKg6WlnMs3uJPXpoMrY/vGsqSg2c/BdO8c5zhaeLS6rv9
WlS/Qfao/6U/T3vZR/h8FQDvhN4TmANevtA6vJ+ZF/SIDG8wmsWgPnZY6NjsscEAjujDDqILdtW1
3j5kr/x7wX7WDspNiC2K9OAkqxzXmzB6/mVpLAXjo/IXFwOfUrqtkAiINF/5Xu5D7vPREHWwLT5D
1YlTuDVogYds+DQN/J06qv3DIiY4o8ROiZeuc2FlO4jh/7RIuc3K2nVWxuquP8AlEFGL8ndWgCI7
m511LcB0vkmnzrMBwOy8iXN0Qn/5qqno0wQqi896wsy3TV6NDzqvVJoXCumIurIEZbG68gJMTxim
kjijm4hooPCvVLWRXXKSZSrKrS/8XRFzj7T1/NMRncMYNhcvCDHV88hLZQgPnBHDpTBP03QGNUXH
auRgFxLv9e3YhbjsI64YaofHXPtjYJ+DiXgS61XVIHwjRgVkwKClbkw1PxJ3QqBaGe4KYrbdbG4R
Tgyz1OjGAIAuNbMxHtNDZRcksyfpDrFMZkhOEpjgOr8/WYy+t7nmAmivtHMqYPPAhAgOUc5LmDpR
eZJBJvphfiOOzPDziHqyrF+W2fjwrss+b5ZigAvWN6QZjGkaw76ln4wcVcEpNNwMaky2eMZU96kq
/ggw4Z9pPxg54ZwJrQnIMeQ/csq1XN62x7F2bDmdcdsCo+LqemfCZvyUCZ0yWmpUPdKa/dQc+Anc
yJoG9SqgkIkFeuyhK9aDfhr7DXhkCGMTX6E6wnWnzZ43ZHmQ3RSflbWjWJE/puW+c4pAdVn/pEl9
JwwQKG6s1wsiluKXMcFqPiy5RcfYswX/7XhIIlmSfv1YviLkBFrYPNrByFybk26GiNKQ9X65V2gg
YouyGNqsL0wgrJ9nFWI7+tp16MKrX+cOSw5VuEntgpf02Ccp1batBnREDz91q6hrF9AtwUpTR6OV
v5mB0zCIjZyfLVqQ1pC733a7dC4vL1Eg1BsfgBWfy9kKjQ7eSeLPFifx/rDda6YAgoGnY8NqiVmd
iNldK0YDStatFQy2y2vjNVGp17yCIWV0U9l45VlWksM95v+Nj95nBSccE/Ssvcq5AFKKMkR1aB4T
FBN97F6hIy6QSHpH5ONz9qRZGjgBQx2sj/2hESrf1LwWmG68tyYIR7fEgQIzlD6a8dLZnK+05oW8
LCSUplKkIipQnBj+5kBM5cMI8ysssdkORW8GK4oMZSVonwttm/XlIovS6ddYQ5cboHkBv508cGTI
iMYL5C+TNsntAD1kIWecIgbgkKKOLll0Vz/I/lIeMsLx05+FzS8DFv4saL7L8K85KCm60OPnvDOW
VAy8L6lsqCSwZe3h90L0PrwMXuony6y4TfbkXB0Z2BGSxmq8ochwX0EegNBgD32unNvsojk+4zBq
z9TArkvkNlXRC2a4DcDUCR1gzvzv5zcDnPPCXrCBbZZsop55vgUfYQskSBjRv/m6di8hh/CJYEVT
K4AHfDLhbD9YOVGmboJHp4G6/CbwPwJno+kL9XyYmePuNcFTE74SOQQ0C5mdODkgMRDnU/jNaxPu
BSrV7rjPG/lyOP8+v6NZKl7C/TdtJRZdfxbIq/RvZ5bntfkj65VtNCV+LjW7MSpaFXMiSBRWOpPK
+I122OTbYgiEmL8BuxXI7qeePbYR+mDIRNu2h4xmNRSN0bbdlXI7Z3S9p73KSsh4rga3q2kbWxcX
whR43+gALeAQiTGPbDavcVNSe7izZDJtp63/BVra3VaXxvCQtyLG3kil9Uv792zLlqIHx76K/v4Z
rEKaIhiV9Q+cVUp9nVeqSfxXEPw7om3m8duzezZJ0IP0Qx8PPkGuHRPL4hTvIzMZZtX7HOiIzON9
ghHfGtsfKnrUxq+G8sxQV3UNI6JblthVE2iVm1FuEdDUKe7k42+eHZ4T4dWXA9YzaIGaIAxyuejp
rMrQ1nAHQaJUgfJDTVFdAelt469OGe+6x+SpSAHOLNmFhyGFEq5xU+IeVLPFlcuRk3HWMqV+oWbi
FclljdaCsbbNYOhf+GWMspwfoVDjNBqd2zs3hA0JYaQJwy3AZTa3lD+0VMKC+33FpnPcHmmaOi1a
lhuhGBI+yhL69UR7CFLna+hS7Ul3k4PUHSanh99LdcQoGsTC+elESKZKklBycj7tEnQrzMK4ovs1
qYGczpMOAs9GuqBUk6dGWblzcLGDR/w870kARXgVVMoXYTZ6L0R3BGSFxBhXEqip+Vx3lbS8u3FU
dowdfO58mtBnfEaAOSxkkdvpS/WQC+cfm11bt8sDRB78s32Xv8hZu8AObMmzEv6kxRvmK6UIATpU
7+MXMx7ayA09t/2QiWMqzjc3DtY1oFjmxVqj0FiLx+pWYBbawuAr2GPXoG/YLHc/nBi7CYpDZpTv
KwEkz/9STp0moA7Zt4fvJVP/MyjiHWNLqZeiDO7gqw3VGlvBkQNy48zROyxpl6k+eHEcV+LmHxCe
A/IfE9rj5IdimE2vUx1F5IePale9HeVFGVNaaoUrR3oc2qnMUUM2XydTqtaQF2tjCud/e4gF3MAS
OXdpDWWYAFfyLn6egOG8SWXsp9L6LFQ2pllndm2SlUXJV9HcpJADzFh1t3/UYfREEE1ogUxBGl9c
PESSYy3L7eidAK2L3+3GydHUsS7LOAdjFeERyp0QSmGeefpI42j2rvCXLmxvHLaa7UDWwyfOXpI+
0eKbq869AibUWQ8Msj3yj9s6W7/h9q0OQKmdoW4APjwb3oBOU7C801lRP5utHKiVNplu0uU5Hxzl
Hk6gAY9mzwpPAgibevETwhvnYJ+P4e6AvgeQIpG25uxnUrjGO4ayObXLDwnTIVlSsqTTdP7oP8sp
h+mFQgdbPSODCav3zx6IcWccoT65+YhOQB2ewHsJSzZuQD71pE+KxSTyNbbreKqGqu3ambFe0g6l
1B1UeWyCicec12cQAALbyPNSXLeUy2/nRSYb2qMJYaoSn5BhPacKK9fcyqnGQgdoIvuNEL/VwSEk
N8pV772XXC9wragsp18ts4NALhifhMHopqMwd2e6RxRi8cjnvNTJqIsORezADk5bW0xPjWfYViVy
3exsPcPHoXCPei9mX93DcsdgF91AXmNEz4cPJ90feiS6yZOlqnnaTvk+f88DUwwrHv+IKNsfEVJb
xXlNx/DFiznU595a4D1Zv9S/60bFuMXdXYQDI3gL/aCqWgiYLpFVrHx5p+EsgO5/ZuhDCaEFXOsv
A8UJ/HpA4Wxsc+V4aiYX1gKGxk2XBmZ5j96Mzhn93yXLwp+h3J5ji6OGKQdR4pNB/KCOY4bzxtp4
WUodujz9L2CGuZ6dZ7dewQiDRQiU9qnIzCXBaaOhBdr8bx8mTmYQ92jdOwSXfiKeWz/uZR/yzUJD
TFAhm8b1QU5KrYektxlF84uisNjnyX2SWsksNEHfGTTHDfUkk/r2zMFp1T4AKryTD0VS0bCND7yZ
aK/ADI3UKDgGt8xFuPGq7VoQohBtbEcHJ8fRn7YbR+hMOEH8mz2EbQbN/BsvLL/vHT06SzDdjOlf
ZZu27KFNdNA4vMaobSs7abfxXkTPen9TKwbQ2DphA1vcff2ufpw+FKwbHgFpUzfpn4jkjvQiwMBw
N+wYTEta9c+veWsZhGokY8zDk/yVftFDZgKprwz+YBwf3+IRcFH3QJkgwEtqXSda4AMqK6M+6ZxP
u/LhN3oreOrZqMErtDv9+Pbn1+VKWdqyDg7Y5vig5zSUfvmpudIEnuKwWQHIdwnw0PI8REeLZJdo
pqWYrULVR6RBRIRE4yI0NTmVRWbBSmF5Ank2TTaYh9t8M0m4vWDDoFyEeJhX5RL/jzeejw4WA9AM
K+GIFKdp46c54oM+IzlJStN/LtRQmO+uUAnlxg7PIXpH4andOOuoSP3fFmNFObSph/llrIvo/JVM
2ril117dyxKyHTNiLb6pQteVNuChaAVFIqLn1GvsGubSwRfe7d3iLGfwWkJaPi1b7yNlGlL/Ch30
o8kSUdajVHqTY6pqx5fBKMGH4XtXrP/mEeUxA9vzvdpqAQD5xBqQH7iNW3dKCvG6S4lp5vJ6sDE1
k5bvpbrm8Ni4RvNFgl+RHXzJnl3SmZJNqoe1A9vHozNyX3HGNXzyJcveukcO33T76bDGMT5/IkGA
KHDrtj5mnBDDNZY7V523ORu8WgHb2MJWGV8qWZO5ZaWwgaibmWoMuWrXwqtNpqcqGWtxJnAvFMfD
D/gUWPTTGSt6K96zQsSvdmX6HHzyquzfr7mGRTISX+uqfjeuB2OU9P4O7VhPC8Trn1iHNQSPB6h9
/t947/0bm8v78lHrzmJKaRTmQPtvwcChhMC9YjAtduuG3GQjoYHD1EekRpLeerTGAJsI2Kd//dxx
9tF0ILnCB4dmop+juozOnLAQZxtEO6aWELtS6Ert+aZXhIyn0GdXuaTbW2ZtP1q0WzLLoF24jTHW
H6g1W3Ys4tYNwmuOgWV9+6CHagvK2jtOhnR/cfJDFL4a+rYuofigddoHFlptgslQB3lv/iRn0SJH
CLxQC/l/UM5qQeOsTBjKI8cdGdRCqqshd6mnJpfHKroXiWTLLDc980I+/CsRaYOvfHEqLdIhv+q1
HEgxvGijToytxOUltWhQkVuxkXYiEZhwNjlrqsfAE/RGcwuYzavoyKTvfof7Idl5JKst2hMsOGl+
1WtaoY41GaeqFnXgN8X5vxt7BOLWCJeZkn7ciY7dmVnpyJa5wEDX+25Bi4HYQccxlN48EFrSOs4M
/0PqcEmEBxEXEIXf8CRv97cQel65OyRAudtqA1CBiyCmDRgErBETMPFgtyeDvzMbYIfzSvQg/ghk
zAfpLynDhIgI00+eYoWRHzEu2t2cVkSuNP0RYEtfbP7htBxslVpELXcTjaiPxKESDdxlBcd8qj33
BGVhWH0wL6qlgpbbqzoG3XPDZMC5aLOxIg3RoKO6Qqjtaml74LTIdX8My91gOiI2ent/xuMW0ynz
lErTZQLh0sDe7pmDq9VM5L7QV3aVJ8ABUvX/NMDgrxt6SJhWxkWWBhO3z0vpzYEPqc0XFUDD9mh1
aJVc9sAC1s+cjMerCQziW8WcRSiYiy57AVrEJ9keSTCi7/BTxRoIo/yotIborN90EvcHgcuF51/Q
D4XPNOl5hVZNgdtL7/7MdPqMlMIV4+OliJCgBW9MKvtjIDyvxH9fxyc2rIFevJw7x0es1ILZuvVC
Mx/mGBvuojLbB5eWqAHC7uYJ49ZgM+3X8zMTUBd9uuYJ64y85EbzW1rRupHH21kBBK9w0xCBngvJ
zXuqDUWvZapZue9fHWuSizEZQ5ebqlKcW9Bow0EAHgspRC7f+w/C0sUqJlCvv4nA+YB61IHBD74d
TV72U6tVGwiSYk8jlOxtHdWCQkY4FQvIH+SuDWihpU/lYVqiXi4RP+on+DI1AImNaGWRTn8ShM8x
fDj9kEL6VUUQE/DBL/WujtL1ZEx2VN/YTtTPX6d1AWHmBhFQRSuyV2oRVcOPjFJ/fLTRZzp2QrdV
tStXWUK8fD3oYC/uZs5KNAmhAMuWCg6K/sHHHd6sX0EY8AVDHKN9fDfCk8ENmBcS9BJCRHswHpGD
v1yr78NtxsZh+LqA8phKBV/EgGK6ymlmLjZ0IJxM6hH+zYWJANDQDxn6LxDm6KSYPwbZj5kHICjx
+LjDz1Ghi6+u/Br4PV6tiVzhuUxjPH49wTkOEH2EjZabAjTiOA+hgRDIkLg1y0R4j9lZ8wgyOa2p
253GnEJ/+F8czVfQsGac8KCTxlBHEobNSZ1z/SOYfQdnZPu5AOr8j7NuTIL3eJjm2daquq+CREIq
w34O1dI9bGGW87JcX19XtkfgLxixZibM2fVK7gE9xkoWddOOaGONh0AdUF+Dgl/Yy4jnNfi1cDNI
XarF0igwlNXgwB+SNdJ+ezhcp2rqsJBuVGM/eG0tSMHCohSuB4irKvzC7RADT/nCBKpA3trcJiwU
e2gMmLSMUi53whJhYcWoW5h2GYvYFL0tQbVa25KB/rVW085l9CxRaEOEO12DMlUbqF+xCbb4b2fE
SbC6pRMvEADZodIIiB7MaUSIYezrCt0OrymR/d1lg7T4pVgzFoY7rU2wvXMe6ROKgoobAr6N2gHg
H2c/QPW9rZmiQRoZA/qUDlqt+8x+4ah6O0jdgoD+wNoaHDU99EvNnB0kiadUEQuxEva9/OYIXcqH
aUGwcrzhlBEBCXSquO8g+LaOHcbODXYAzwAdK4CudNdk2gflVJJLuw5nVUW+eSBKP8FzDkzBitPr
tODh9oCHaimAX6+KUSguCYv9+3xTWAf4aIpxwu+qhj8V7HnzOTjmfDzTXzxH/ANwE1nLU3jnwPUh
GzGILNgSo4hZ0iTMkMbR+24JJBu38411G3a8Q69fm2/20Ksf13evXj5b3YmDQ6ynwdzp3KfQs0G/
SEzBcEWFlcXRep4cIEm5+Mv7Fdv2iQA3ORmd41T457KlHo0WMjuUXK+QbLYp7sqUeaPSG2zW975t
8fftsBUQNbntSF7kNANRJFttYOUc5MnbiSeNkGz5AVJ6iNhE85aJpgcryZnJY7ZsQ0CnsW0U5WKV
UmzNOkavmZyld9Li0Z73HGyloGmTA3+h+1EGcKjaxWXEwYriWjoKmBWk8cVgzkMHpYoUE4dBmYCV
dkvi4gGq0n6ibJWDCgZ8Svmoe00iAlURqME8z2oFz9NoohTQgbHAuTms6hjaz0GxodK5SEuJONW5
fmZT6M5BJn4FqGmFgIUCk/Zyw207za8pQ8CYncLuNi/DVQVIZfBqfhDRF/kjF3iRjbIEvFdBH+95
3jIfPge6pGFvKeTMhKyfA/61xRxpUjRUh/olxI43K9s38NercZWPlm1Z4hVITRf/+KC8YFfQH6BC
IHZllIf16Ww+ZG8w5CkRik8BGgFFECzUhzEr6pvspuU6cG0vaiLyO4RnrCTdhWBldRDlo7z6Q+jT
Akd0NqK0uEC/JE5QznDRIUJhMYPrJ/Mn2Gz749aumBgrqHGYai01kslg4PTpXtPJA4AcmB3JYHWa
HeEbPwPw1FFnusoNLklEV91zOmaA4iCN/+smMMWcEOJi3Y0ooASRoD5smHgcQ5CbCGPXNqKlZndM
CDW4sHYHjEbdeo8xg8n0BuLHtBjNxrPUqhgfn+H8jm3Hecn4xxeLB724BvMfmwgq9wSmN0YH7cHm
842RoevrEXvQG6p/ivfsqj8bGeaVmJagb1UWShG7HQi3cBZzLBhQLrNfBYu0Hvp6ggoWEJ6kmE/8
1V9DAiH2yXx91CqbQ0NehsRul2umL35GHQ5/ofppdLRMpDx5ZTsb4FaylacqD2QG9iFGv41EpVJG
PhRtNp7sOfRYij7wQuAktsCk9C6rgZ5MgxjuQddJ0saqGIZ4vNIIIE7mr7EQoclDPwerqaaYGIFD
iVXe0kry6jI3bt6mtGdAPgAdtQExHUAT64aZZeyzYR66wyJck+rp8+KcQ82IiSN74zao+En6gVXT
hCH7wUulZsd5nwbLSiN/dHqUCKQAorT1QTGikstr2D4FKSia5t6rdKQzzKFAsKczgVpIk1lGGxuV
QLShKnCnypOB1+inFP1wT9b7/FLIFdCzcPNRSLyA5QiDRPYDvwCrFjZOEIEnpZ2M1P8rBTatLGYC
8Cm0P/bCteKJ1aVqvKhtPAHTVIkPatA1UtRwW0/nIsIMyIfo4i14l5qRRDgbc/cu/lzjHw7Eb1GF
NrTnX8WbFcaTsE40Dku3KFupc1JQFSezrbmLJ3V1d24Ef34WDzw6vfJy6PeSAadYJ9zBeVklNhlF
HqQcXAMCUhdsew95CukrWYrsSIhxvMPnE4Y/QF5c/NeLyaQD0KLveAEqizY0OPvLL5HGGGK1z/kH
AmCo/jdP+8iCZDpXOQBfiuTQ4QJN1Wwdf6BWHKWaNXtUVsW1lKki8uqJ44O/evXLUWGjL95QmpCT
mVLmc4f1E3Fb0e80xnXDRMcJH3qZMCPfPehlifOLrCGqPoeVxddw745fdfOP9I+4lnE4dgc0rtSS
CD7kAhZc+i4Q9rsJUcYeqjw9/YRgsI2zzOkHM0GLqZ/vtant0DQSqiPxenXTZ4k9TYDlGPItf6fK
vHhnitA7s8OEUrxCc1V51BZDMOH3h2/UQPPpZEASKqh/2HIJ0j+784AGrQSGpKgsF46gKZGsZvq/
WUD23JdRPUH/LVymn0X1KnOP68sSs858ZHoSt6KdGx0PkuESXDoYEfWD3Nb2jjOKLdbM4yw+2sCW
Dh7+ebKUPtJt0J16wseh8lJU5CRorbKid4k2SFSeQxz1pH1lmqKJLDpjF1/k9EFgVZhdzr5O/ytd
jhYO8S4zyH5SOsZ20sRuJfysufscSdpgEObzWOGExMPobdjoxANKio1t79Wy216F5s3qulbGBXcg
J40ginQ6SKzVZoYEtAPjEllz6VKpEuL4fFqfMMRRt/z4I8l+HS2JOBjP0ANHu9rZeg9TQquJT8l6
5yqCtTkqB3v+VOHWS9KQ7J6OTtdoq0WgsIDWNSFqEy3+29JJMBqv87h2zaftJnI5vJgMmLWu2KVO
E18Jyw9wiaa9XS5Cr8I64VL+hQtjZR2UCjdW7ggHG3w7zyei9iek4j8Xum/VD5A+bGNmj8RIJslp
qnTI47+U+6nGhTaz7YUnIZBn754SGfK8ZdYcTTwH36rsuAaxNimuA5Elvf9FaQfk7tUOY6ynWWE5
DprAfflVM056JCoGohojjPVNIDPiZTjPVWg2k2PstIok7e8ieLcdookeg9uBiPTZJQ10UFbZwUWU
edStzu5njRS6qXfX1M454Hj8h1t1mhVF/n/YShcNijs5ShH5HNky5tC2+/OmJCUHv3ZXkXmi/z5p
kPe/dgkfRJ8oc30IaY/FPntlsykZ8QBRDWrDP60fraxZvFiuo4+9xWcQirF/2lH+wr6HC2cYXpHe
Bl0m9Uid9/7hjYwHligfpxNA3qIDQ9ir8EqSsmHGKlRZvWG0wxjzRt6FRFz4ma6+1IPsr1mf9618
a0qbZw+BGp4DAXeceAO8b9q8BRkkLK826lqrhcxCbwZVs1gvqkWz9UqxmvKBqFpntjfdeP0HlBh3
00T6qxs5oj4rA8mFlJKnL+/ZFBbqkTG9sah13gAdbd6C8txvJYUi4v1t5EkdpY9Eg1C0+3I+XDHC
VWSol2Gm96l09JbyKUr9aD9vLLlXr1rMCHKJjhvUBfynvqkKKMKyJb/UiFi58Z9zGr7oONQ4V9fU
ZEELPmbknWlHhMCuqOPl7S9hQAGEV1r9LbGIH6VtfpIIryWRCfh+Y540U3IEcQJQsvNpCgGCrrNi
vbYwJDTKnvVeinH3HdKE4zmFxIIFx6czFfZ2Kdahuaj97Xh5Gi7UMGQKatie04RQ28hElbHNKhhs
9zCHgAXjfW37XACmGMxlCE7E+KLOdt3BM1bghh3F1aEPW4sZIGjUdCzE912yeTBuAPF8gbvB6B/g
V/UBTatFT/H4hCwvS0bEfxRBkoXtjeaTpM33dDn/jzCz1W5g30r4aC5Y/PtFvhg5o7gvRLUMdn3D
EzA5hmt7iYKvE3WWi0Mf8fLp6csUAq4FfKsmA6h83zRKpfOraVUj26KheJCwYbxVU5FTQWMOnzY/
Z7zIc9XfL0ftYKn7Js9FP6GRt801m6huQKUCdVu0553Wa4Mfctq5Ha6rb3tk0lFDFzkI6tn/5NUf
YyQzt34ArsHZEDfp8+4kTWqSjCVoLDCyi1s0OZeXWe6JTs73oPqPFUirrhoG4kJd0d4TNaBeKV6T
t3T+APDCTg0Gq8UrPZdGm+FZXA3UVefhcMfo8E8VHZtO16fKRI/uX2VKHvesqVGg1W2mYWiQNiKQ
ZM7likM7pQSP4C9/MzHQm5caaqqCYCgSQ3Q7JbVKcpXEjvKPWYM2pl/NSUOn8Wk3dxMM8Lg+Glns
3HKrUC2xBSEgU7T1FD8g1cgcNVOvdj4okuKxo+y3g/glH8yhpIA4BMskfpPfweLdTW1i1L9Usz+o
fAxJdTQCFNW791p2J1f4xehH69zqFyZdLSq9DJtGC+r0kuWBO2WXL2nRd+kCvq0UWUax/vAdz3az
Z660D0+HrCvkNIoxflI0OVCTUMtta9rGb1PlPMpYtksqxqLLN1VUslBxvaF4bKVAXp5N4UtaXF+4
E9H7yPfekRulH5VdWquKSwoKzW1O8Ru1J+mEC2VZdqIs5m+161hFZ2b0ECZqBIvmw/DqADAO8ZNJ
urNdTtk4lxxVU9qZs7EKffmPsKOCjHcBURiIuMSVVP3tZ9pRjM+vUD9sVIzlrYP14O4UR6fRICi6
UG2YgyJCR6mlwn2CNe1IjfyUaNW4cMk6ZvO8UTzzcJ/iWqqIE6utRIcEoHXgDXpomW9zQQCa46lT
b1QrGWkc+wHQkBOM0yBDeL9EIpqlLDCU9gjdicOYiXFMeEhDXHCc61GIjPUd5zjVuTseRyvNVz8k
X7+FlVmJUnxlM+SvjVq+4E/0mAPbOmwGWraFfHIB9nJ1Mz5NHYREHj4zquFDxI1S6dR4ve5vjgyu
7ThUueGCiA04pdIGAxiM4jzmT6CZHnAYrCg667q0xOUO+ElMM8EPAwkM+7lpsuZkaAJw/02iobzf
GFNcQSt16EiVgk8GG1XsZFgNzt2m5s6LJUVAXmNDoQPA544dAOOaAR3y0d6oqq9fBDzDO6rK+ZBb
MdX336bnvziYsql0QI6NKWnOhwKUG/tLVXBMazQkBkuuCMNrKTbo15Ep3Vlbe8dC9AntJaMOaYA0
oA01nWojAcg46skUc2pWThxIbTvj5zHZI3cFRMowZVEGEuRpTr+q+lEgwSaQcYk/cIsb60oI3afW
HMVHvyF2YC4iXBLzHTG+pocEa/aZv8JXWHB22W4HDps7Z5DenCALuzdtNlos3FNFWUKUBfPNzrEk
/p9L1CMfsDwePq21v6k87Z5eqdBxn+7LvWLa+cSUW28fvdv6eUDrUeW7R5e/TPavf7rVe69r8P8X
kaZj6sK7gLbwpbhJcuscFrmi5BsuwxabBT4Igk/RgXNzbCI0KFhrE9D/RVXzSgmP7m7efGYcgshO
2j4THSv/qROZnN7cltrCTGrHsteC3GT9cIRXI+iIIRrkTPex2yKpUJFFnsgUZrzzVD2hqQVUiaXa
byvY3Sd5inJWk3zPv0TeZM4oIkefSV3MZu+bkYbbUSa7GvcTze4K1N5uJ5iQGCYx7YTCwVog0sO5
4C74q8vYNoy2sbjV6fdWb/vDN1DFvlqAOJS+2zEwaxwj953sDcJkbMyeEv87BN01H9uSYhTxNB+W
lCG2WUxqc4aH3GnYMcW/tvIp4dq1aJ7I5vj+zBHqHvBo9ACk4mKLV1LFZ1abC3S9umlLqBI0D8l4
bDjyuEkYP3F9mvq3Jjv9gHBYK/jlFFRAm5/IIIvHCcPAmLiH8BLDRO9LXQMeU3FsfHdlV05ucBma
vxorZF1nJiLYbsHggyMizbiYVNZ0zCxecu8YFc8DDUPm/hKgls4f5BChpHjM6VjwNJtNbzS/UKey
FIyFHDGQa0bF0zO+xLR1ZR/Oa5K4YkQI3uSISwaCm7IU5lW1xwJzXGWCdNdpkQgR0fTbRRSdjiCR
5W0W+zVBf5Proy9DSdJm2CoIc+57stTVBa5Tr4kZxEm5jKWqos+3/euOYX/4ZAeuCsIW/0KxdTHE
2MrV9zymakiGBt504ZlMqu8TXr4sUIS7j5rl/oNm4i8KObxduto5y0CcvTzFXt101ZROVNValQGS
rvJSNYHpyBRM/G28E/9mwdXV1hQcYHqcoBGUXQXMYWiroXCk+2rcVu1SXwNXcus1Is4sgVamVMKn
200lHGwri9ywwS+lw2suj9RfqZ4pu9WSOyb97990iE9zQj9eDfW+DI5UtgBFKRYEFnV9uli/ABiy
fvy6FhWxKXuRS89pgprpd2lnvblgCOx+nGI+7CQ8kbhq0Qj08Ji1o8dR70MamMnnrQ/HVrF3Bvps
4Ls0DbK5mk/GPNMIAWqvWgMFcLzQKauzkjbv5XyJdKwXrvUCAlmy9vBw/i8PK3DjNYXFhP4NGEcJ
Fkv7mFmSg0hJWNbUozC+z7scVe32XQhxqQKi5yZYKSQiCAXLjqGY9Sf2W2Nz9gmHxITF6nYotSBi
ZHUe7WZWb7DWlM866tlJNXjQks/hWtrkAQ9ussnTxhcEAph+0vK8QR/zDfyjS0mweWxoVLLYTtMe
PJBacBL/C0mrF8oaz67oFRkaNnL6qL/arPf9HwZlT7bCnCBEF3eCyd8Lw56onxa6N/UmFIk3ssFr
GR3bRNK8Q4xCxvtG7b2ZszbOheJmFp6EMYTHN+g8Q97Xzkk/uUfKhX4AY3IugWkzSFKtUM+Tme5R
fmsLSDZ57cKuCzzocA2nQyRdW5W9wBqaIOVczH8XVzZcJJOXrMi6DnAGdeGXeW5ikUPZxMioZChe
HW8s4lYCOS1yeD7i71vrHq73YJ9sbbWR4wjtCFcdcW96bjd1Zi1PyypcdihLUYrUgUhwnBkJ+o42
SRddaIUHhiZjy2+EnHgMqa52nemCBW2h5Gx0/K5FS7gqDHVsUe1sJM2OF9ckoWh9qxQeOp+/EdI/
11QymQ3jHO4g+WpPT56DrDhchyIY77tgrKWhEuPpX3s39GRW1KkIxtFD107WLUI28NonR+oTckTD
hmU2kQOJ9yvd4Wejegala7bmQteguwR0ahAR1nyyiEZzmMS9auljvp1tDOqPBn1weLpLM9Whecrl
IfHnM07ociTFlzZggaZNL80oU2BZwLExoBCphjAULVNC4UFg4T3b0kwElr5xI/+exlhB8skQGYH8
NrFIUgcCa+XUCCtyuw2Hg394QAv9IY91NSB3vITon04mp98uVWn/zMCOb6YLaXVIt/qVr+iItYFl
WsrFwD53RvXxLMYenQ0DrUlLaR2wM6hQbedF72R3MTnuVf5IUbDIIZp9PuSzcOBG3SnLt2vr27aH
PcJ94oQjWoupPJJtrm6JjrI4Qf9n6W7FR29jfNDLFk9Z5eCwzhEvvWJikvFA/CMFDsfPNbmnWbsY
m0d1uwSfDk9onZjCp5usQGYDdU/1+N6wRwke49a1ksqwj7MeBo2onEvhRvl/PF49891Jo+D74Le2
+mhMSHSoLq+xEPcjJtoB6JoI5EZaduRcI52iRD+jgqOD5oXBi8TppuKZwja8+gZCMl+gQs2HphSb
9DagyP7wxnCWSJrUX369H7mlbDSKi5WI+rRm01ZMfrTf+r+RBh3IbqdyjR5BbJke9YKO1chUgjhR
Je0ulVK52R5zwEU/VS4xXyVlUs3fKVRafEnsI2TLfJtJ00vLoVxq3GanuI5lM2UltYMCsaUJNhHx
FVTcSSm4SI/Ve2MbpVfGTbnLxtYv36Vm7srCUf4PcZzLylccd1AYgO4QCd1GDDmJyqgdl1A7a2oK
f2q0jN8uf1pJM8EdxaTqe0jBy/rzq2HZee8VSrU9q0xSOceAq+O/4C06gXDSxXqnQWyq07FWqUnI
FqakaCNGvRw8xqvEn1GMb4qtoZNJ4S6W+RZx1EyeKp1hMC7j5R9J6MF/4/X0yIU5dqvavQxHg46W
3cPWsaVYSSyqOJBuctpaaMGWZZFPIol4XvValbH0uSL8SOfV1F+7IQwGnmYVCiioK9r9RZK1Zxvt
bkB76LaWX+WpoCuESiA+Jfzk0S16/0Cmt31RJOqUjyXzKUxqxcqHBWKlmh66LY/hQqfBXKDlNenH
XwwIqnbHjtw+qAHh5Mx2lJ17wzo/sB4ugnBnBEPIq0zbDOCIT2LyLRu0pBFbngWifGkDBs5th30c
K+lMBLzX23cz9m016XSSnh8EZldV/sLLWlASw/Vg/LoZu0zScRkcSXuoBmixySAgX011j4ox+X+r
At70iZbwyrt+CXiU8Shc7QQpGs65WDCnY6xPzbGcXosA8vmyJzp33lBT92QMTa46uKc8f7WNl1YO
VIRP9mDCge8lzmmXB/laFTxEcQ8J31nY2OOWSoDxVI7ZhHNfTaQKR7JFvdsxI93s4KIqKWj2w2f/
TP5UEr1ouhEsz/bu+ybQKNfsF4ayQUUU7TBaMCFva88SNcJElMixeBd9OMH1bRQ2gcA1SmMbCvoS
JID7z7cCSyEwDb1RGVg/AGkJmvjEplV0H4DjumX+Z/cdwKCI+MF94G86z9oD1GHYm0pUlzWenfNr
Svz1go1P0jPJAa4E8fme4X8Lu2xn/HJlmfl2KLp7RVBwDZkqwATCJB9MLLp8D4/QmA7MHu0v4aP/
IKS5mPtFFSIbMz6c5mAnpuItY/1PM4B5u0VktdZM6Cl1W1lZrVvXdmGspUL+HYFMv3k/f38S5m99
iWIdm/HOoqO0xnIOFOPYFlSzJZJwZ68+a6UFcINjDAnUkrafjBDxDnLaysrjQCd1fL5wKRUApLA9
z22hIZcd3feIAfpBi0pBX7DNNPGNkeSm9UfGtnIw8GQG+PGjZLOCjI05tyZY93FsdiBVTedOsBcc
/fWjiTgw9CLlSyPnPH9N7+rrdJ1l05Q5RqJG6n8657umf62SokyEk/MDmIcCgMjmirmQXrYmMG1Y
iqzzlxz4AXe07R5Q5oMjgmvZZzWNkd7SwOlZN9KfuHvEe3/WdQ/iAU2toj4yAaP3EXRPXe2hyOuh
P9xhSUJAPs3aXyXu2ISk8oxE2oSVDeB8B/G79Jex+sITzUEkJ6xPZl0df0Hv7dpiEIIQge3DHQRd
VtaYvgfJa9ECVvDg7ihSn17jDE5NUBF8gZWK77SG21mZrlTA4gSNFWC+4jFUrv5gGginwXCV5/Pk
qRl2fWjw6NWxAUPXdGzP7zjLOEcTgf65QfSDJnPaBqc0kDzMdrBLGWI2zihFh3ktF7RDGwlmg3DG
ePAdFaz9tVzEi2Nk7AVxrYyTVB7173bGJkdzfWa+774skguKmVbm6GgvSVakqrVyHOPZiONz/43G
NJqgl4c2YYh9Je2xBeV6dPFh37c02sLOXdFU7AuRpZrFjc6UItRyEpITmJPDg/Zg7Xn7DSmcfpVI
ulv49ptH9IXolLR/uaD26450aZ5hYczM9IRKVl4L4d/C5+AalaVys5MAgDgKc8vQMJ9saJHzLsuf
GJcfB7QEQ5IAn46I//7bLwUXq+0VtREcxftQJ6knDNGVTyiqLUHxOz3W6/nzSbFCWBwXZzEqi92k
HzSF0cQnxwRXxbW3Qxql0uXejuAAM0VRzw6XJJLpwy3wVOnGai1Dsa3WAb76AzvDSo+WBxXSl2ri
KIWSMoZHCkrf5hTVTyxvK4P/ppgl+t+rChLm1T0Y+rwBDkqAkYKRSgHvByM2qbYU86dthpcuDtss
LnPqd/K20nDc1yN1vwpHGWowdD3kN3P69ZQGXvzmjVBCM9JOakiCGfj9kO2/2/x+9kqEnmBQ/fxT
7Vc7j2ryaucbe4zgp9s43JV/Pf8iCsvqLxr/8wZTmKqM9tFcOFm50kQnnXTWh6e/1XhfJJSIvD3I
gqDLBPUuNRuIRqqBz8FnvDKO2HYAcSzWP8PmDP8ItT0ys/kUcTZ9o9Coig8WytAbHwYrbsZqocRz
GIuxWL+9en0Zc/HyPHsYohAQ5k1E41MrCrbhJm8WgJ2Ok1K2qXXwauFT9rDwXYHtCn1m7Y1gCy8r
txV3cnRXaieLqLXXzy0PxO23scbGC9ZL+DqF6Qt04N3KmbyH3HcnHQpccFaTh1iAwNRWeCdjyJ3G
MM7c6w8gaHvIMMPY2P6OWRfd2ljs/sAC5RIc0yuDuoCkk5ppQ69ox3mt1fVq9yc2LTy6SBQL4+c0
tCffEq3/2nNl+MW42iDvDx34vPL7Iq7S+69JYd8pKPMr42YRTM6ILrP+jz/D2WliLiR6XKtLbt1e
Xfc1m2/RbCRKtBbBSqY19X/7owc755fPTG0HTmqIrnZz3ePETSAJyTN26YuONXDf02cO7ukG7Qen
hZb98eQ4Brhg3faMe9oqugS0SHa6pu3v6bz28dxE2FQlT9d4hNqVrLIeWJlefi2WBvY+ZJAaje3M
e6Cbm1ocfvWw2nxpG0j/1k7MocaeXRGWH9keGdVUBLYt5EK30GlQEiaqkblR6xru6E8ussrPn9n2
5XjEe6FzyZOjPHfNLWZHVpQV9EeKq1Z7R8uEmNqZW9Wc2VF8nq9QwetVVvSM4kGk75HP+Ro7xOsX
Qzkl0GflnnV+qJV7/LLRc3O0i0Vewz1YSFOJo+SVTyJ51S9IF8K6YCt6TbX/J73PqcMfg9AbsygW
VjWMqW7AJw4FQqGtRWInI9MdVosqEYe1/lKLCmuVjEhRSTKfpW7z5SnEey2qPOodZht+jPJubj04
wtvONpxd2l6ZC0yT5FAS5sPUPQWIVi5EIofmGOo38RvXSlXm6Qww5Cs+Xtq1sU882da/TCI/XYX5
UQXfw6OolNUPQFUjS7HNmIe3fjr1XJa1biesRixfF54KI0bXW76gFKKtvtibeQ3QHCMw5S16Fn2E
9scCnnOWjb6F9iSBUn23PC1nOp8pU0Kll3ZprJs/cvOrAQnDL4gZQX4zcebvAv65EMiEq44/zBWt
uZ0ZFTF30ou4381kzDtvybf23cR8eCNZJcDp9fcSZRfMPAB+TDmOu9JU4eDogaEefb8UeiyzR+yT
0Yna+hAEugyl/mBtFNnIBpqwkGMeyFbIee/h1M6X8GZUPrhApPVFS6f/O2NO6jn19zj/YD3jPh7S
SrSQFMq3VJZ4Rne2FG1/fP02l+EmTQMwLkYoQd+aCXLWuCq05LqbHF66LzBfHHxOsY3nfVjBIb0y
uOQBJCYIQY7YeyGMTCRECu1SZoNsdr1J0E1FARxMPiD3vY8RmXWxB8kn7jiFuWSUPd6xgVyuWAqX
FjGapN5iSxrAE1CY8KYijZaNJzA4oIfQgqsOdY4rhf+Ewz+8e8anEf9Nb/t7ydHwgDBWlvyLWe/o
KKxi4Q1C3ljpUmlMQIb1wjSdBrK3G9VKlOCTK3H3c/iuqmF9g++jBgYoFTzGUqx/WiMFdkYIBheG
eOu/8GBJ9AHJCMA+Qa+wnFIquiiyJghLklgGisk8ik2qSP0PUjaISqRkECrzYtIsprC0IBU+BsLB
8f6fRghSUDDjHlfqjrFxEirgjgHSqX3z32LaZGh5Tq35VvvE7Ad9SaXq/IsDm1TP6IFArTPJNz0F
S+Ob9mM7DqbaXsf8WQEphuuQE3jGudapg0+RMbEcCUO8C5HN2azbtrE5JRCkq6vpXvFfLXQTf5Iu
93Pacy8Cs9BSJOgz6KLCoMMKcVXwtsiOSvnHOlrVuZ8AVxVW205N6njhCD1mfmpjNXKeCG7TB87p
zgVAD+vnQO4eEZELBKNkDr32xnN9AWlB1q+0B81uXPBhFjYEnVpWUUgcTl2uw+VEVEBfyXTBY6eJ
Tf3aUFYiKilYz9VglZHU7iBy5APuVfuRuzBmk1Fgfkor9Qz4eau24Lmph6LU991MnNLEGOYhzp7x
zCKGHm9JLzTYgI93sQjQx4ArFh0qfjmZvklMQ+VwjDNMBISZajTnmv8GmKKO32KkXQ1Utzjrtodb
ZrVJk4L8tmLTiF88suy86FBesFMlR747Mn1P1UQtaCokTJjxTlMlUsiraDiC5hMNgS3a1eZHRvqd
u2LzRsEr0yeUqoSKYkWeZ+UxmdPu9Log37WduMqDysOEp8BFLYZF9JR+LuwElM7tPvZNnxW16aBr
b0RzZFWa57/ZHM4aF1fGCKlUoXVZD9ELqnSyiRbycxgINxrm0tXhRoc5kCUeJfThDR8NyYRexvCU
sbEECSyxLazg/EEi55sMkamFmvmWpPFhsRpqhlwnvm3zLgwIn6Wj4L5AehJ5iLfF0l4qBgrHItdd
4HkvuGSs50sEx3N/9DWq+jeIavYkDtCMZebO+9hB/aa/bJPu96MNnIwPaZvLZxDg8imq9tNZNnUD
eY14GQNlVhKjM8KuViYmR8w6pcQ5HiVk7c45Li4AriC0tTgb9eJ4T3pmmW1d9PYafh72BEk7Wx3T
EwzJgBO6A62YsKfO0EXFcZtfgNjGC1A8vpoiDS1Ez2tMHtknkalxnBgKUfnphdX5COcI7G4dhoyj
CnrM5uKh9BhjjkSaLdfVVsZdlNdpESExBWNQmQ1W/HgwT7l04HCqIJOlzsyrX2FQ/gVfHqsdG2+R
2tTkf7xhXKgCn09QTD9pFY4LVPREeJvZty4W+dpyB4C5sf/QnqT4Kxot0Df1A90ucJ5t8at5apZj
+pgZ7uxDyFluyNzU4/RX8VC6TDAelHNzybOfDhicE8ETiUYQlXKAE0F1ITQ8Cse2EuUA2wPEsFXb
ramq2srWmBax1WQwMrofMYbzh7nMbN7LKFTJxih0A/xoL4ONdaBeJTvgzTRPDscX4LLujq3znNeo
pudiii5cGnV1IyPG9HZfBIBG/bJLlwO9OuIAL++BR9Mg7da7GYxqitmoNPSC9LLGZqpD2oRUKIKH
mYdoXXWGLTSi8EmcR00gA2FbNvK7Dju8rVSUQTk9PZ3RmWH3qARqCpxLmumHjHvIWdxlPMLvfA8H
YOu/woBjEbPJ96JVClAprBQBmIIOWOkK+nb3/5FVhvCaH+iCbK7h8SdNIhf8CvIl+3Shtud3XcCI
AQW26L9xC8RzkVtUqPqvj73auy+Szu7+SV/GWN2ORFEdnlz1W7GVsAYZqphv83J71HYbyAPF59ih
zFdQitLFGRAaoWy2oJteGEbSSQhzg2uxg38VtMTCFy2oI5lpLUpRdTU47BBjmsPqK8UhqqSWDfmd
P55B9pmQ9kg3ruJZL2QQFrlCuFCcfvcpfSSuKVbnqGXwAVLLaW01rwuL/NIvJBC2BuYy6Rqa+dDT
Ska90a5LHbf2Qxk2Wn61/ZddWJLCHDRqnzVySRPARLSb0EnHoLO4vMcyyGIxTSlhT1ZXmv1coBqM
x3UjI8847j7VdeQNI6AlabUo9VAO2qei2xY3qH8dl8Br3FW7YWjOHuHQzTU2A2RBoKoWLwEafiey
6NRswlc4XeSa/dPmkhmBNEsQfeSJdfG3FwBRSAM7ZK1i3wczjiCeAWn3QiAB6QekBRWrkd2IP6YP
yaoAvGSU3DGqHltZa7122f8dK7uqVZZAx9doewNG5+ftBu/jiMLrT4JCmSScm/CpZ9D/LY3ir1o8
ArUI3+A+tUmu9crAHnH4VN2WFU9y0VUldrprPRdPPk9mZtYlhc6JjrILLcOriuBh0tBvclN4UWrq
9t8DnuIf7QnBiD2K3G0QPdYISdtLwLud8cD38PK+GpuTuCaL6ST5wkr2myc7dZjY7atrpdpkxBAo
QlDxDjakKDws1cGrH/h/VqQhX7pmQXaoXIxecZwiQM/Lc4KXdtTCRku5hJ1nu0/amNSWNHN7eIkL
ah0ufk5OvySvUL8H7jXwO0EHggnua/QPzqeaue09tksj+T3NsJ9rCb8MAnN/vFrzNN+Lb5ZkpN8n
u/azZ1g44yYLkXUXgD3Tyx+OlVg0QglqPp+2gaK6Wfn885qgEKUpaR2+1C6fmEKlDyTP7+12KSCn
fW84pGucn0MpeirWgBhpWPqLBa8Fex13vQg6G0xjILc6z7iM1yZ+fpVDOJSVzbAZOaNWLOU0nt3b
X7X11scmKAq5uvu+G3/M/NSMyKgf28KGHFKjegvPwzRRrJS+G3RO0J1QZWdxaFzURNKLWi0tVeUl
OEpM/+cjFOEiUUt+9DGSEwgv3jVY2TtwnRDklC9DIiDfoHh7r/RU8rf+KM2xKuuFtzyAyzPzAj1i
naX5I9LnFAXkXqNrv6vnUdPE5fdeduBRqaFZhFqgedAUe/z1vs0tgsY+xzHdD0uPZkzUWcW28jzA
6br4fE74hI9b9VJIkV83I8Qpx7wOLWKjI7hv1mw2h3AAQSZWSXad0VreIv3KKX5RTS2qZW7dfUSZ
xocyWfer++blNFKDyhr/G7KpTmDgJAxAF7iRm+Pad0MUoVJJ1UhqIOyvfmDqZzm/JblQ9HQ0esRc
NDecoLbteqiqeUHetdWTOmvOBtBw31ABoTppb9aCzombqC21EVC9n8Ojv4FdHEb5NCbe2nGC+djp
q3qoEa1it7j+ppaYhydzVofo80HyZEWjzvb2zIbCnG6IUuyKcN51oP46zuF+vxHQfGUrewXIj0nY
2VLvezuo4VyEbr75lm/pFBf9I47ib2LJyTAcKieQXM1iAJk1r+kk2xI+dI+Ap7ivyOPXbWAGnLP6
ldukbekuBeKByRQiOfQNHf4xA53Y5kDVCqm1k4PAINYZLPpfVZjwjlNn8tiPvqDpLGscG8HUkq6Z
KgsBKS4lr0QV3izvm4EFY4cfTK4J0QxxUfV3aoajhYC7iZbwz+OEg9x23weyS+iuXTuLmchkGpGA
SxEbXcS6la4bgjnGrxDNtVYTVripGNuGUg+P4XquKcj/2VGFvFw7USiDUrZmbt1QQzLcibciTfwg
LXDFUvOEdCVtJfOqY04Bk8XNKrSjzi2cex03GUFo3hXXQf52PXC5eEhSf6iPIHArfT+Lx7izOgAZ
cHgQjoaWw7odQWKIwxsOGFVMXKU3r4YsEgQZLBEMU40ZS2mVbvMz/ISvOgMBBWwJMWNhBPs7ljRR
j6joMc+76+6bY+VMWD2jcf/7HH3qFTaxJcPU9uFnlyTTbqBDTiAaep+bbI3uxdYuh26PG8BItOH3
NA1zwEiMXfqdu1MCLKhq3vK9b5CHLjV9Fwk7+Lc9kNN6eckLrxkK9yE2vkokP3P+tqes7K2N30No
uODeloIHnxU4xWNuPdRKo2AyRPPk84/eLDghiBtIgWCeVg/vxFdr10hXmw9af8vKHWAGIA23EFMg
LPnU1CxE4HXmwbs51CdyPShnV05bniOtJTW38ZVqvhogELBMyyxISNw4tgjUSZ4iSQUn52/wo6zT
PI+NoaPqiRVWkYbr/6nwNIPoLcLx2ZNBbP5dyOCBqsrDJfERFN3zhwiTeXVXt0bVwNvAxccmFsF1
f/jJJIc+fxZYVaSBnvKsEowETUUQ9s6+i0JSaFe9pBfKzkrvVX47qnqx6oi06qQ8tQTtW8rcYWCQ
OTB+ttDhj+OHx0IzH/izhi9rtPLV9PUtR55gSHA/iWmth6QkTFdkCFBxDJ+dPrf0oCnpqbZ+lYm8
pSX3kpQEtzqFk/DiCuIX5HNQaazvVObU4Edr/u5lPfFWfTWOFKuHknLjRRQLwpZErz8R5QbrylFc
mSWaDhjRurzbuoJsG87gViaTR5yl9CbHGlHSsDnUf35L0h8CsxxAi2ggWkEg7mteVgzSfG8OFfuV
ueHzUVAOAWy0zrb6VIG8rGyb8c8c/T7XounCW8yphszEYXNZpDp4dSnhjspBNV7Sydv2J0uh5tcz
Ise3oAbpEQiaB6hg//XtV/QLrQze6ob3wIO4+IfLMqRLYDbx2tFOT4TZsIidAC88JiwC2LZaruJ4
OVyFZXcrAseB0LEn/FQoaFev7Z8cIjY5EazkQEtTRYGclbm+gg3qv8xCRSBL/wb//8EGuzCwdH1r
Zk5hl2fF0I08bUQr21dKEAhNFgA4uigeaoMjAJeXsWpjN+kN2D/oIIsK/kOjAthcV46aAoGWvmeb
Ty84RU0xhxIAYkFZ8fzIfClRCvv1asj6ceC3+PY8IK7rTGY3JZ7BL4c0q+rh4pa/3OzoXyIXyKVU
10Gx3qODBXmy7Dzua/cdKd93JriMfs/t3hq7H+MT/ialIK3YGF1YWUif9f7ZpvWmcDatW7Vxe1vW
kqQ4s9aMJSd6W0g9AnQY9Bq8gb2r/7U+XhZboA+xxeP/TV5KMZEG/CoPHH5ZHUW3c4eDOfLjIZTR
KYlKQqlNRdrhIuh42ef+fXqCSq3fuj9IQL5ZcWsdj2zS8Ia6dEOM67t9cXVzz8vWujfZcgVyu09x
hXUAHtZd41/DNg8NO2hquzlF8f7TFp56ZBF75xN7p63yEdLedy1PVMkEYta15OMmlaFPzCRfEPSo
qjCO31S5PJsMUX1gHz7Q4YBowE/AKHd07OvXaCRKAmAQelJZYhW3E78wEzbPJ2CiBPZ+HrKhpMWH
koVtkbaDwnIBjP4hbtUHXbSEzCj++2FsBYEV98EhJbuWeq7oYi1eHl3pyW5t7mi5dKC1RvPSWdKD
0qg51Y8G8xeDcIjFgMl4l71m3P+jDKccMH0JQ5km3LNp3qhEh30+p/d78N83FaODf8+lRtOmi8bF
S5YJd6NjfhIPU8FW3YAdwJVPSxmzI53cvKIftC2UUN7FN79N3Qc7iKvwPvbSjdbaNS77ZzE7lbGr
6LFeuWHceTd76h5jZEY7WbKPX+gkysfgyINjfadGEd/tuimwgwinKcyacHjcZfjEZ+k5xH2FdjFI
IVSDzuCSruiyBmwwZG0OnLrNNajOt9N22J3niIWUgUvNLeOzj+r/hzsZte59w/2dJYr8TqCYWXNV
PPe0GBBFWso1of0l2/Qpeiq+0yTIMMQUCrKncA/9FZovjoMY2Zjwn9ZSm4l7+ZQgxFFVdHzhtyc8
8UAHSJEmuZNMbJsDM/O4MH9VciU4kdwOqHf2OQwbAD7XPOI/w3zxCiC1e6O/ZKMIJ9eEGCRra+xW
LvVvPEm4Vc7/hPT2n2ELjVFnq2vVam8qjG56IWZLnrER/3AWzvwhFAWJ6Rk9B9lv5+aBlp2vDZ9b
wDqRtJFMwQGE2hHLtZrJfkmmVzSzL5eggsHrZJ358HG9gKaDridapaCK8Hy6+qzKOC/0N3uhHJmO
vjaWORchfGUZshzbtNpN8ZhIyhJOAv7gVH+u2/4yLIL8LccnsgtnLn0k0sFSZjU1YvUP47fkjFN4
QyTvvgP/tOMZ9dOej7cLm97puYvnKUnuIx8iRmaSUR0sOf3/h+ct05RbGFPU8QIrrtFgsq4m5dY9
SihF5L2Jk5l/LZdb56+D+m+VBCHIorpv/3hgJoWdZxIBnYwPiDIF4icN/LrWC9CHXMMVciDO0Qpb
YFtcNa7FzotyXZb8fgFlklEhpuhr95hjL2AXkE/xpWg6BeLwwgysga/U+HSgPGyHDfk5M0p3SVxy
IZbU55EnzVH1UzH2JGWCFSXks7Hhc8qCQ4+E1jIh66wj86BQiUMnx0EPrx0A8NQ75SGPoEZhgnYN
qKG74LoR7wrrGJBZahWowHNVjcmYvdMuEP8Lm6k/Dt/4JZ45xNyTS/B8nYFcMEPm2v2jCRE+2Ur6
HAbQv3lrStg5I62clIeWQEWGkhTBKS4m1tIGKvqWTqXrNcKKTDmoiIU7RDTkuZu0cCdXPaNA5SY0
OZsKREPl5vmAKi43WRVSKcv+e0OlNCEfJO8gvo5GyAboBDnPVJoBVwAMx3kq6BGYgmgin07gbwRS
OmZ01z0ojOxAjrbT2hfK8he6uS2oYEXCnCKCmTZXiOMi2mzQG961kQ3AzT5XrzaEo8KRIG8FTBxk
FKp9ncP0QarNXYrzmYv16Y57+a1rXdR9lMWM1SMS1t7nV4FKzGYNS1kRp04qiFUTT1cauoBf0Mm9
ONYI8oDgXwpVBKOV3HjzMs4aNsX93on1uCGsNwshGrTjwSFQjyQFxFu4ANCYKGurTh54fndhU2S1
uyFIU9s/uTGBfawiive0KTPRu2XvHV/MuFk8n+WEC2HCbN3iL/NZwTGP5ggHuSDXMFwTiWiVtmiq
0AoGtj9UakKbS9cuLP4M4V/ezWUIr4o61o25Y2JHAR3uUtTPPTL2H4Pfa/QLCl9FOiEPZm8inzs2
sKoUCtz01jWzma9l6Z9z4vLnMXTDr/RNVdouk+zRLrU0xXnCIs83BLH4X0G6/PjI7z74uUE9/sEa
8mdUi+J1PtiogUUn51Vn0woi1nUeD7Va2pEh+6+ALyaxn/aZtyTAwMjzI8ScamcMQPi07f5xSdN9
oGANqgb5MB8ZpUfCMuTfTtLXBZ4vGO5ES0VrA99O6QZHNYoFMLIFDukIxtuFZ0w5dMd3fmj/gpKe
Z2uiVBcra5TqLFzO3Wa4Sobibhw4DsEyMbIr7v5BumMdMBOOMi4X1rznTi2bZuoZBLZv7hQeqil1
ZmdboiSaqiVNGCo7GkCWXhTqYsFq3rhBJ2uCXfE9Ix1ESsMWd3pTxtPMdGKajKvn0bc/L8vs4B8Y
OJH6UhSdfQxzTrPVA7f6pB8yDW/IR5HogYk45H+11XpsEqG9rBo25Awd3FuQl1VcvrZScP27RpKn
GT0qQSyOdj73AYAzesxZdUjiWrT54HsD4b93G3OkdF+rSP7efPJWD7FoTTmeaDzFVWgTFR/TqWxW
tNcK2RQPk4PXPuDEzqRSYOqqu7IYBExhgA8LbTszmttZgeLb/6WDs0Fl/5Gzxdg9UngBTk4/a1aA
v0eEvtJxXX2h3XnfqwhJV96YcRzUVhYVC5F/FhtFuKpxnKSzNmBaiwi5WEHLk7JZQEhynz2wg0sa
vzjZV2m4H/rEx1YpRz9N/XYkDlvsVuYtJTPt/1m0y2z+sT0qUvOF8z1aIuziXt3M4y+CYM+bO7WF
9/6AfzPgR2huE80gnRgYR5C/7IpgT1Cmj5fm2hgmbexHC5wo9fBrkhrRFPu7ntjOGuIlBwmt/FCk
2Eua/iYeAv8u/iwl0a48qq6X0ulqFsfQSUZnNNLXcaIipoOF590LwJ0UO8nIagx0t7xx4Hft3Tti
Bpi9UnY1qp+3d5W7oNNZC/tMw/smH8hcaIXgHOzW3jGugKUeAUEn4EfOCBuM+5FPDoY9s35BrRsU
JSGZt44OJFkWGXmToSH9h147HQ20WPJVhI+l09KT/wEEEjFAVTlnKYK+ZnP2rV/vmFvMQoOcd2JF
ILnYRcK0o4XD6VwoKBl3t24MORDthOKwGN9bLuue7iczEd/VwIc9D9Ac5LrHdtCJzlP7aHX3S31r
CQs8T3LAQEwWtFgjqfIg+HtRHli0GNiWjF8sgCoAQSBGQcQ1G88riEgSIg5yG6GJY5+F3It73Kyp
Wl9AJgNhxNKsGpU+s/3+h1qqM9u4dqSSezF6431MDmS2V3jto1zrQdygwWm+CbbaaQ+WfJbIbdrP
g5SdXvhbjAYhptWCvZ7jJIzZjAKIe1sbZZcAjN9Ag8cbgvwgIJxFVvkD237LVTxpWkxJCdAr/eUW
rVdWJ96wJWLPpxNuVjdi3H9N7aJZIxqHIsPIUMxqdkcWFlEvmd+v5jQS/8psKnVWhfbftYjMd9aV
SNp5JemW+S3CG2YcNNq9wdh2W9Fs7VmpG8r0dbziAM3HCGmM1EFsFMsTHosdjI+IbGD/sf+U6M62
MPbyQUCY+sDJ+7j8w69e8dDhLNtHCYbZs2cmephy6Gm9pxNolAEVwAUIZBHGP5+d4HnrbFgDwKjX
oc1kVjoJ45ZbSEAjOYZbfLwUXHmDVj01ZUaAfj7leVg02CRj9rmeNaie4vBLeeaBIZNhAOZgjKHB
lMLvbm2aLiumCAQSReAmpuMqSACbyZf9s9DGDwnhTBJJwdfJ5nA5T/NWKjTyWt1wp0cGPmKLaYTP
0ZDCGdUIDr+02VmrEMGsOhinZdt9t6okRXfcPoazBeKMGCrde7g4VTRiZTq7kPNVpnMyKIrYp2rg
knN+WOfVi7d1WfY4NByV710eDDs6cL7YCBpNrwPkHHwfaUCkb/eXv2Bk0DnGaP6tH9jwhw2edLzE
YZnfjuSO99dQ7qBQmzIlZT+K0ONLdxX+HUOw0tWIb9k9KyazZi3bfbbNkoG2JzstmtV6YZ9ZEwvn
mENIdPhin+lgDrOKquE6g2O5OPdnqu4wHtGEZRAGdMjltShD34MpC71tkxkiuz1Qh+WMB/Ut4lXU
z8cBHarOwaGPG3BewvyVrIe78LMlIiVgM6fQkDs4zXTf+0S64P7bsfnLZT4OZ7LERr7S6vY7PdWs
8tYi6Xvz34WOLlxDMSq68kLmYPNQdJkz0Il9ExPt/XW8chDUZ2Iss0F6lR4QtRCH/vMG7rpRmuTT
Bl88IVd/mqxtFds+3GJg0ScnQusnFM0hNYMTa+8bo/a4j4naVXWgM3kgmiUgm4vAaEgnGZbb/7HN
0Iz6x3ufTTdocaiJobQkR5vFEb/P1gqtgsaP2+oCdo4Q3ynSAmK8rN/Mo+pZOzYpY8ieogINCDFG
pkH1SEWQtPf8JZpCACo4vq7vKROU3JCGTRKBB7Yeh75/ZpB2iWqUnbzoCDjy3X8LxqgQJt8A7QRn
sG+iPTv35iBh8HLjSE0OX/3Qcz6WnykDBfvmGVbuEA9eOV+eYd+VF/WsNYRVrkJVJF6Vk6sN10AE
jkqylvBwRZ/VEgLdNKwVLG8kg23NXb64GsnVM+gkQcL60WphFSG3h/sLb15QuLMiFAGL+3xw+b30
fNRQSep/pKijcNEvk5e96rr2rvd1x+n1PfGjYZ9ZXyKNAZTzEULhGP3h9TG95KqkeAdsFkhzyb/S
Y23llwxnxy8cfM3Uj1XoZXktPV8Aa9jhkG+C/w3Uk7JIEYhczm+qdF/aD9DtB9aqxg/04LRec574
PsTZ5vkuitOimE9Vltld1zvvlqEpRFrmZjvXYVBaH5Qooee2Xo7hSOgTbtysE8naQcirMYhPBK57
mG6g3YZbXHx8u2ag/Erp1n2gvg6sLRbvlO6rwUistIDLP5u/B/19sT61asts4EwmH4l8WUl5vOU6
3qmY8jeizVnHXZumelT52+2jEwdk/x9pPyRtZL1zYH3hfpui03QRjYvfqoJPFUMbkM9SbpqG2nuD
qme2XXwVySD3pyb/Azx9iuB6i6SWCdjwSkoIf6dU6kay+ShsyrpBtNcOmThX7YNsXQ81poLb5xHx
hyvvYEyCGASHI4IWipabDnOSKlifxCAGfYgQgzlheC0p+fgcK4Nle4U0+RG2CUc+rR0Itg7FzC5T
4jcqZv12BdFA1Q/F4Tpt6BMcdI0cy/PcOBqolQnnAVquK284dLceX5rxry/URqJ9/gJrTFiJsEHn
fxPrSRSYe3pl4q98rtI99VL57gWliDDDinZXwose0zh47lCXRMa6Ka+3RWrKENCZve5MSaoOkyGH
h4GOdpQtpcUPtq9P0q6G3BPfXnSAASWz8M7fbMo6C1euXadsxMP9QjjthKu91+5VJNB30Pl/aoN+
g/WZMngxIDsO9BY5gEOcSqmxoGb6js36tjsrq+KZsCODdfiBqGrdrpT7fro5FYPtQnjtmeAeqknj
L+2cxodEU7d7hVmgB/cBv+HmM4mwtnYuTqCRtXsDIQOtTQO+nHrUbmcQeDT4+TMD/aOwJATbhjiw
s66MjEx2xWluDIaSwoNJNe0sHdRPynqVYsOg0zKFuK/Johc7mOenn+sz7rYQEDT2a/5Q11c61AeX
+QSuQD3UCtvgaC7+uDG2SlUmysAtR+9HaNsTNoPQeyiAkvimT8QFXdaPsogJb+bve4LkZH2qt7HA
PBPljebaTbWon4J5YH9NnciG8W06og65/cYJRgusbX1Uzm2cv2mncRR+jKM5DfERfbE+qe52Tzp9
W08GmyKyvLRf3hMCPsNarVOaM2ng6vPVAUmqcv/D5gmS2yC1NKkmmhH2yFOyIcoGFNZ6mbM40rsM
qjzXcC1akoU1m/jAomCphXjhyRpZNhoB5iTUAAMaCL6o8uTjo6NJznMQYsSuIbKgvXk4lnaYIfxP
/P3zKVfjBUsuj2xMIM0vjB2RPJa4eTY0s5pFqx0MbPnOu6EjbF7XHUJvEaFWyYen1l3L+58a3zCq
FYPN3Pt/ndmZkD0aq70EJRHDddhH2JU+Uz+980lA+B0QjtIj13Kf6RkJ8qHTDdmIx7dspq3iP6n3
yaXpzVa3qaYqsrX8ixZ1AC3UNboRjmfM9I7ldQhZDUuNiV3rT8pVVexuwHWybJzS5jVjumvzGlI3
bu7A5knFRkh6wJYu+XnOo/mhy0GCcgWzMLBYqJgmVKwOFohwnOFDNwfTCzeAOrUF3FEq+VwdoAli
a5fFZyuT2bkTll2/ASosMr/mki2CPnmUTODJnjSzwARy7j5mdVfX97CwmZmVDdwiTi1gWTyYwhrJ
awkTw4RiVB6qyD+rqg65iA7IFqiFAwUlJnHbusr+OU48tfUnO5iMe9yhmgDeFIr+LMhodhL5r0il
k61hhXdCFbCWNCaq24SBksRIA3GF2E3oPFrEvFOlYZZMpZMheGS5BrgDIx1VLWDZ77YjrjEXgBqn
0lZeQTt5WquhMXsbaWFLkaWZgGjvHxLPZ1snit8FXfZCKFfH2GO3xn4v23Oa5gDWI7rGYehjaA4J
iiIPvTZx+uXsexHakkxhdnFVnvm5BHUccXMptV2pQ8f5DMH7Hmx6Hh/6A7O+t6bo4eiW+j5EAbEo
WAGyDRhAzXAm2UdyYKxjbEsstbyf0P6gHTuSV0sN3cvcGdeAtDkoW7boWpCklb5y+QbmQa9vykFM
nv6h0pB5T755/7OE8BD8UceGRXU3dlTxKlBIyjr0uzqarqmFllEsRp76iE/ncvafnRbB5zJFNFxe
VquuURgYl1JYIj+voROdzjXtBsvybcv//69qHi/zQoc0Ut2efSGOz2UVZViggrR8+vFAFtDLJSDT
Lokb1uRgp5fMwsn9keSWuBQDKakarhAbPcseeiwJHU0uCEbLRAb3AXgDJo0rLvTjqV8Wz5d96xwt
mMV/UKe9wz09OVaqQL5VRnbcpYBER1PeOjiPSxVuquc0/ZnlMZ5vjUnCJzTfmRMPDSAqk+Vzy5ul
nTDSwhwtOV2e5Wca8VV5ULKronm/4tLUCIyB9AwJ16gqwQ2mqIZKNbfaTO0RYYbE+D2NQf98tYwZ
Z1NFMUOt3gwh3xUgzNCde3mziNUYDXIQIYlumuUytrkLtb4X2w11x7WvWJk+ejoSRkK5f7D1LIcc
wIWfIgw4Vd10X8dHsckjbNIWGvWqEQhPCApwVt0jVt4NimvvSKXfcx981c3bWfQ89JBc47C3a7W0
QjWschvR0TYo+YQhzSpBfY14KW4Gb9V2zl8kff5maBNBImtxBhp4zyuuF1gh95tjk0EeabIZ3BK0
h4wLd5Bb1gaI9o56GKl+VgR8y9cdCOh7k+npSCSI9DJPKjbb5kS0FaUiBLspYHcOXp7h6lGK36Te
wZZYrreax7nCxvB5EUP4kipFramjCPzhvOhzNXDPb/zX4CZYBsPQjQ1gbmPxhB56htW0/dJJhT00
fVAvPcLoJfDagH1IAc/4oQgHfrN4QDj56b8d1YmIo/Wx7ZTeBv3FB9GMZAIHuFb0SA8/8CcLeMhP
bglsbUlJ/mF3kt3hQ3q0SIGx6Pc3TwdN5Ij4QN5NGaDIaNNiBumXn20G6SD+2FzKZqLf423LCs7R
sI4F9y4/dTUyQWLgIsPvqh1fWBitGIIbjC3Gocrerbr1v0+0jP5E483FjgKhUU/b+iYpqZyQYTpH
vY0EOEVlvVqWg5oghqeZ/DejdQav3qcZ+csSqK8cIGAK/NoROT5Pv/SfTY5sS0XemV2du0tFtcEe
nDIH23Q4UKhGTWyjKsrjWksw4oVYptwB3iHysrp5GDVDAJ9qbWWYMdpWj2WHkdFx4zS9nWWcJxeF
zdiYtSnb8zMUI/zcG1+vtIxyXnUnZEtd0fhwyqCmA5OccTT6l1mnGwAtoGcthVyX58t/BYDz9wQY
sdMYrSqt/MOHn6K6dltQAdTXZwmMpvRVx3QWLiX57Z45kfLG5+55wGgVBBIa79W+EJam25c5wAy6
R42aThAYP2/TnN1UbN9ElYL0mJZpucyUanWi24aH94Shn1/8pSoHYN2BX2R/jGEvBYtRnvi+qDs/
Q27FoDFuyo10Ne+0cKAEXBCGd7rU/kkXfWoa5lqU26dBx/FTrnyt4/n4YoRlkP0t2GiOth9cN4Yr
E5Y9uPdS6WxgKXd6WFqF+VX5A96Beuz52PYzpicYI9lGDUzmm6v1Oduk/COzpps/+XyvDcoNYB78
e1ERQJ3ONRPgA4Qik+im6ydeC5SGkFtIdxN4z/b+/EtMv3s1+7nDBeKZjiA+AqUF7veAGIVLolc2
I1r1lXqhBI4rcnlGSD1eLTGoI2cc5EIIRjFiIvKDjH2TeLo5q5EyK2g67jqf13DNdNiAUV1y46N0
IncYptROnQ6pqBxVcjr69oAJG6havxYkvScCWzDm6kGDNoXHnv65UoZmRdanHGMu96n2juIVgrZk
gFsXAPH4KkxDKXlcEyZTozJMr+JkiaShu1aUfpFHYiYHkCqZ6rb0scWOHWEytnUGPS2Ugj2f4EpS
w0DIuB28Wrtt7NDfK4elR8rf2xs6jFQrAwbXVFPoQugpY6GgJ+x/18fp+XRfKGBbzaSkUZv3rezE
1tk7iDVJwcxkfdf0UsC9QNWfUSzt4oHwpCU6wuwjBodi/MIDSBAJ0/0M09m5FkS8CFG18DAYQboY
2ZwFSVr1Jy7+l++uj3W8RudZ1bSJmJYkpdYdDTdgXEx3uw9xvsW7dRE3UAlEoZOlsqs2NxCU2ZOo
a8roVYMoaDfNLx3ihWfnd1Nlz0ke0ZZfJvMPYS1TMtsz8jlWCY3sPwMjoDU0ASZGzG0mZRhYXLoG
KcJ86fB+ZA8GsiWse3zB3Rr3AalR0+vVzbg1EnONoi+V6gNhTPAqIX7/JZHWY1AbpaaG0vBUiQKz
0C7X07rsMeWmXaa9wCaJzY+8Y4+f22jjgDabDCsE0vGSpkgdtgosjJKaX/ETiLe4iKC7nen2f5CQ
+ngm6fL+zxENQRB+ZBS09RBhb7uvVceMQgJYk2pl7C8G4lhg3ihTleUh5g8dkU7oJMKQMzm1IP8+
8nEbe50vz5R+eVcHKNQfPzWg2WDx8oVpE+N686wGlMWcgxf1OV5DgQXgDc6306c78WiG939+DAG5
s1VI9tPGf3JqRAS7uLZLwdjOpW4AUKMg/fRg1IX/kmFOVRafnRLhIctrmgCAEwyWXEjmtSDQmYag
4E2BmDwPo1qV+4rpwnIC3ARSCzJHF41S4a1mGcFikDfpa1B9A3AO3j4RWOpxBc14w+bFQqKTJ2M6
GWdJI5HK4BeFGB6DxCNE65j1bA3N4ffVVYchc5sHOeBCWcsZjFelTKp3txME2dDL8R8kGqYBRxFR
nsQpwouG5mu/v1G4tKsa79g0UjkR6YjX0kfaS+naFXbp86keFphZPvBAtgixySgMnQKsP/CzDSMF
1w3I1xbu0e2tOAh15+Jy5yVBymzj620K/yjbAsODeOLI8/Ec5YpoDGugw1rJwRYDiu/ofThyrf5l
WM1NxY8Lfanf22pDe2CH6uDgjQb28FZd0GGinh4WP5ZZemfnZCtqsXjmuKJJCG+VH+4QeAGuahJa
gI2F2upughwafKtKEA3mA6vk2aZ7rM4I4LVNxYTum+kEkRD/vHQmr70odC+vqju3n4iFQKa3g49w
cF4lF+Lh31gSz1sLxRnndoj3WK0sf4T+A45QpkQ2FbvOOkJQOndaMDIxnQcoi/+hM6nSWyK+d6zC
Oo0m+jBxzrFXMahBRokxucAhWSu8wIYtseci5j60NS3g/1AOcxXdmV5sS7x1u1k9NZsy5x+z6vrR
46cepF6BiCe6XaqZkblTVu5jlFmHt3a3PCspBcj7mINep1jBNe7kzNM3H0xvOUTOP968ii84kRPh
p7vqZylP+edAbe8z0J8/he1Re0zgk+fSnFgn6YSde81nEecA9lzHzmvrcxxQZNDYLDk35DW0zhQu
bsrX0FTIvZhj36z3ZZ01+TuQiD2vmwzjCXKfB6JMAdno2Wbg0wFqLN1ry8dvlrXMdUDx8Mo6yl1x
hqJyeRC/kSTJqxJpxhrtpTh0kJsBtOtssiSA6BStHE8z3nHf1kVmile9sNlRQgC/OZ0hkDlD9UO7
PX/aluEcP00Gp8HX306u18K/FeKClXQIOFdD/WAw8k8ugMnGKoWXqDprU++4JGosA/ozsNpxz7C0
YrZF/jFrMXDg2FM1rr0KlVNqkzGToWFW6yU5KzM8CLIBcvd82Ots9teSXVKzgplJDjaq0JjPdyaV
oubEz3fX/bPseiDwsrSHiDcVyTisy84x75dSgLPnkkBpOVaNZ7zI/gcGqg9fnAssVOJDYfSp+N3E
LY3JdnBhI4aC1F1Qu1R+C879d/Q7o2j0IsSTFj7FxhxmwtjJsCD8aALF64hWYrU63zqHLdOuFPLc
6aH03+LCC2wF5E7bjaMPpcZUnikREQWDLf6E1/GqoQThdthcxPQ2KYizLGIAIzz1Q5PpeOVmuz7d
JJvJzz5+id5M4IR4+ov49S2yJtN5y0qvkoOb8BErgW9Xwyn7xz+0+/ic9PP7Jjh0pLmCOpN6bOwW
yE5r5IP2R300hqKD2Z3pE1S/NBciOotqP6PT6vwAUXMDc0yXwB3dod2ySMlKW950rkBReZ/Dq1De
f0WKCzgEFtaBjAMdSyO8HILCTGVe3nPS3ElHaKh2HNIg8BH1Eb1KK5y5pLu0rnJ3kolonbQn0LWp
c2gN/5pdjmQe+i8O/ddHUonkzNONSic1ecLz9Yp6WhUudrXaFKJcoepVBzbplbStqBVtW3lDPkK6
AqL4wDM8wlxIuOMSzHBVi/wDWtql0c5zlf7uqckmjyMTStsZ9aI4upznSWpvc8TDzqulCvUuXOEC
VX3Llt19YZLR21AOcWxbWovqFvvewS985RfKwdPiduFWGT04Gjz7JxsJZRudmfdUMSuz9MCcys2R
iX1y6IV6P+NgPXzzsjMU77ovJ67lvL2xK2ZjOjgw017s8GWEF2WJL1/05944G6GiqtWOzeflIYz5
VTXqPfhBkDzyWxYLJhKPxnLbdSNfGrkuBejRCwz+j6wJ3ZHcQ7cy/nX7iYSBw59UkWUqufShAPil
8ZJD2+VdizDX339/RpsdTfpwGFJ4N+KFLLfOIGlrfmsTSn39GfWdfXexDnV6VVX+UG04p3yFZth7
U9a9V73kV1h6d071tiosI6+VtdFBDcZTsiOvP4MvdhDlyJYg0I6cysBK2CYUv1Vr3jmz2HOvpnom
0obtcaK6lTIozApgVHeJiOi+OaJql4+3L4JxMO1gWxEQw1eLJZ0mBpfAgukhNj6m1JS0nEfTeWxS
U0anCaNlCjJ0JK7pmVA+mE2TgTWocBQt1t2wpbxaIf06TYH8JL3vFTUNCshAihXXsbKQO0mzXFiA
FHS6nfd240b1YMmObzfOqmk6yJJiDVG571OagDBLrHQI41CjKA9w59cNR/48UPRop6l1Cw4q2iua
oc6QqMLwzRkAZmvHcthzvMoZQCRFDFDwA5pQYyuUqpC0XBu46W7gBPq6YSgg2XgKi3RMvOU+DUJt
nJ6LSmkxEE8+fnOYO3jbVgaQ/RQfS4g60IqkjvIR1LlZd+5bKFQpc9bhav9tJiNlLfSGm+GfdQPJ
Bh/u2gHisGjH1u06s38Ypt/GEv7oB64uD2u2vPQo1FU55dSr4SPGdmLA86krCI+yAejUJ72Hnb5q
6y2xsl3I9pfHaVAbZJqWvTtbBwxbjVE9w3wWvQP3qzIcXY/WMsbzwDIc7MDFJ/7ZihYvXM6I8h4e
ZSUbomebnMg1VpeLfnjtUfVd0PpSW2APP6YYTLyCuoIfAJV0nNqp3hie1DSfKvyXOIkaNzD5i+6k
BrNhpCT3C2mAdHqVAHe1ydGpyaQ1JMo+IhHWUUaOOqdckhOXgirwsrBI4y1SY/ALVG09LawNdFv3
5274A6Dw8F5s5abO9I+HBMTwc5EfdNbGSSWJzVDNQirv0NROTRutLimBQwYvxKtgwjunCw02ZjIu
OwAy9QHW8Z15ujDIWixNKdq8YBFIT/y42wot4neGEOMURP167l4G3wVj+bIQtxuz0ULpvY4d/Lw/
x9jSeM/xb56sCsLvJTOiffEr5gm2ZEgAfbtN8f5acnMsd0kEg65Xx+HVhLDvCz28Lt+am35EJMTz
m80vnfycJOH+FN1ljVZ+RmwJ8+JAhQF7hL1O0YxrScrG1Gjo33UGNTBn3O5GO63uOvfLdfrcovrz
qKSpvLjcEV9QCas+PD9k/ymMjlAHzNG/GT6rlVC1SRWTC0FIix1sQ/rK0GC+lRTQa0e0sh6oAvuC
TU21uxhZ5rfwq2x0n+RRxq8qEyCrreIwPtnx4hLNM0XitHqfseDL31XchfnsCjtwvyc40ZvbtmmF
57BkSRRN2dMvM246+zA5pauTXGiP3OrufzQkKkXwpaBWsVSRQo3lMhRamk2zZCQByXkNwmEwEapK
NEF8FMllIdiinn/qzCWj9nQIVcBJS5FNs/unYAK9iqllrnCfPe+XGQOLgFf9ylJJLuhb0aYTlG3Q
c5P6moppn17IFfE0ZX7CGIDY9Ycp6Zido50fAz+ej6ACFl1Gz1K8Lxb1kzPGee1yz1LviZ/geMT+
uelAEhqD1JHgZMzmhv0R+s+dNSMO8GstqJ4oEmVFnEFgTX7r2MS87KjdBYyf1S0/mcSNuS9Kw0dl
eUZ4r/u4WnQyN6WE6H6+C+ek+tiyX+xVCg9tFfTMU+7cZ0RjJTFOmoE89Kc5Qvro6OKogfJsM4BB
fNCVbr8aLE/vuR3a5PO7+KgnuTFg6prCPwdIy6SHlVuI2Bd2ZwA+cia5wc+cfwEUp2xDKexqfdSd
yLJDDaukm6vZW8GjnAQKGuYqoE3cv4dEB+dTq6sfsvaEkql2sFdIC5/RH6B1rPBDjEk+RH2ydb+d
YEyBzwKN81wqDfNgiyJUNykctsjpLpuiVd4S8HYc9Gd4qtDh4Mv/WzHZC5HCozqMGWFduKgoyoiZ
WZGnHiyYff7WzzAWFGQsN2l4mfen0rTdBzjHzXZZwc94wDGzt1/pWRDOIvB3nfrX0vfE40X+nYkm
KXj27Fs2xrZ8/qwfCAPDTpPg39ZFVtsHMnYaOjdtPltx6V2eYvv64B0qprTZwY5Mf0ZgAskOvLvZ
02bKgpPRymhFu1Hkk/J9REpHvqjOKjqlw8tjGEx1TR/i7g2cbsOazCz7igNWTSHxcP5iLKQ9Wswn
qfkCQ1ySeopB60afwvyBnE6O8EX6uFn2LnQhvMGE8resOqgr5f7Gy61lzkntEqI1Be743JUouRkp
q5woww8kbU1JOf7l/wcTpCGJ/bspOsq7Tbxmepspth1VF/3IuMhYmWrF29a4W63wHQcTzCPsPrAH
qb5aXQPoPgaBacoMuI0DyMxSGUHqgI1qU20ty5dUuv1y3Pvd3tS/0m3jJzgVuzsrV9CAkbeG/phq
8MeZW1TusIPZu9Vv38x6j3oNfUDDPpMcaZ2kNTkiHB4QLZb4rtb/A7v2qsthBOX2lfiLpt0fe6dx
LL+rwwqZ6GDmnD6f2bztHaqxy1b5g00RKaztlEoNnwa0w5fwnM2lSQj7IjkK2udxF8ZjlcDAw4wJ
eXQYvkU0XPcedNV0DdJBMAZX3BBTB44QJJOqiBNilRqhtailKgnbmGKwQ6vyqetqY2EsIwpUKIrk
SF/U9356BvzTnJg/v196iBeGyk+0O89A9bPaR5iqWi2zz5fnw4lekjtLYnu7gbE51ArZ67qcs6T6
9LSYN++LvCNQobjcO4f4rIORaoCTUjRn3ihgNRMQET6bSautaNFQ9JBmUb9VECAjF+qeH2UTC5Ha
5Sbsjzg/KFsZwNr/Re4FAsyKGg/YexN4T0UZ64XOcP6wFeW/mFPyMROfMtbrnsevUspkmo2WBEkr
nEs2TYzrI9cfcxz+7IjnA604a2WBWdQB/Ke0NnJRgP9vC6rhyqBmFhKQ3z8Rl2SJvwcuQinRxmWe
Bofv+Px9m6qvQcO0RX8y/Rv1rQca6sUcP9joVWy6qhdv9NfT/LKt1Mb+l8kl+AkAsuxeb91DGoI5
0kF4i5s7tuILG279Fih2CE9f2xOSBhiGR9cogvuIYUktcZtVF9qJZwV8HvEtuZTwSfsUzLih9VtY
tWun32viM1eVEgzeGbe/oyFPGdrdEQw2OmBiYGNKU3bga4jruHgDZiDiuOAnvsnq6JIRixC/eVXu
xZV+W8sztjzVfYIW5HvPXEjtjy/DQ1GsaQV/z02gIA4tC1kGgWtuaBOoHS5zT2u+rlOQlIMRcEWe
VVWny76MBMODuzuPrMAGVCFgDb0UdLLr9JNeCZD0NptFHv/y98Wggz8U+ErneWQRvDy8xnVZ+hiI
1sCoAnzAoDynTFzgu5x0BFbvICGzLs1yfWkgE4EKEwq9+2cvSrHBnhxJpKb8vD/cJ0k2NCD0Qqy7
9YPKTILIo0y90dqicMw7uJmqRjmmZukfJZVsHbjiW0ikBskPOwM9V6Ax8CIbxigDfToqQIoS3GVN
aGuc/gLFJetQR/5OBjMWpd+Zm0yQVZ+3FZmZz82rPheRgMW7O5KSov9jKyIFXnHBMRJx6yU0+TDW
ljk51yDTdPGOSKCalVey1m87koiyZOXblJwdbLHpJdDNHHbtbMSe1xw8VaZvuhrszcgzGQY/SM+0
1unUCCczMcUacDNWdi77rI7g4jg10y4q7P49yikpWJWkutnsvXzqLhaaSjsCdmN7EpeDztBayrAD
hcHAXck4rY1yIwMaRJ1az2wPy/DOthrbrYZ3yAJ/QZaOtcCPBcRwuY0a3UXZyJtVQskjidB0uPjO
PVVxVoJehC8lPKdGEiX7i9bN9KHXQ5coluyVLPQ7DcPCyO897pGXMqZTQ3iOw+ONEoiKReZ7GWAF
7tILoisBmf/qVy3ZC5YfU7HiOEoXocWBeLmkCRChznPNA1+5jJGMmjtHskQf91T2xJXBVdLpy2hj
JXDYY83RTMI27wt29DLFhe4bTSCg2zPrSBGc9jtAVfvW2jWPvaY5j/H1wUtC/818ZYEeBMKTtXEb
HBWaTcPnttKlJ0/+GBEyqYxBIBwl+9VxjUwuYPh589U/g4bpvmd18EEwb2url7jrgku1RvhsVxp6
Lqe6tUpzr7jylbIxl0M4e4uUHLTwrDqdSgOl+VXP2RK7fFxExbZCTpxBmemoiZRgvpPDVRJXVHin
Et22HLeQCQVvZGXRCo5hpwhhZZTyLRmR5Stenijj87HR4ghvHqZ0oSez/tsGp3JyqGyutzU+vzUk
OYeYSfOX3UVDiMsfZyoBQRJy5SH0D0B84aIbw+W+lYk0ZB3kU2MZ3HfpMtg2A5lRtEg4zRWAEtuH
6tFcvABr6AZwOPCj7snrhub62/t+jOrfeBfVFfRvJpLC9EjhloHOaGGfPKdT8iO0BxYz1LNUBEjB
CieXwyZsWhV4TgvYXszorGUO6JCqm32d20U5/zkdQWLT33HBASHSzY4l4kYP7aE8VAxzuKcHKK7k
z3PoJqKiod5Ug7xBeRRJwDjtd7eoROO+T0grIDHyZcgU5cyJtXQuRqy7sohx2Aa8OUaHoTrcCzOb
mDM2Jh/FeHuzBZXhBT9vEnsiYRpyZ5PUNiTHh+O9PK+C/h/eQP3Q2MCnio3v99k5My6adW9Rwljy
C6xOR59TH73oo0Aztk0cfatqvEhrbY3kyX04bLnX0uLM6m87In1BG9iWMtmLjBc0Q22Mlp6yU10f
xB24fbgxdnt0oTGfawgFg7YvM/nDzbd2lzUkEH+XQGZZhKCp8eoI2Eq5xMXORaAN61D+Oyb3DSsk
WfK2yl/6DrIeNM8TwLJRLFLmCIgeh+AxgkKFui0NMSzdfQghk5iVprKtVNkqcWy7HHvzNOInRQEx
jGKBq3MpfXg96Q4WkCEfjfsPHXNkU/U3mBha57qmYG9CLVVISLD8vCrAP80zS5upr9T/Tlvz8xOD
TdJ2zbri86KO18K+dnmDhkuPYQ5wbU0GyaVlZ9AYzOSfNfpbJBYeJRrlMeepepD24ptBgyKiqLuK
7iQTmyPijCFfBFFAdCSaQuDUnRFm9xJ7N+CmlnE6qvxiYcukHswWJurJYj+hAEQZzC4QP0Hz8JuA
aGOj115LPyjXOe2/7UApf4YG6l9CbsOd+xETDdVzgIsdp7Nt9Z4gUgO/b7O1Xz7cbOCT0I673Es7
GNWZSU1fJGw7N+EN/S677yg87hXwfk8uFLvN/FhL1tiBOijS20txfHG6xan/Wy4QxgkCmPYMdiSJ
dyGpy9IE4acxWjd/kcfcb6qzTanbuOeMPBy+SQOddy4327YAqa9Q5+9g4NeiUZ8lTj1dEp9XmDd3
LlazqkSQbaLu2Z7lcnUXP0HK+G5YFswYW4aDPpcm+s/Cm3A8xDlEh/En38sJwBxuv3f8yWxHdpA5
Z5o/4/AXuuwUvt5+p7yXd+Ru2jRCb5fc0n+e22Oo7YB+8WNpa9CbLpwjQbHu76aR8CLVmXg62SKW
UbllVtvZj98s69DnFK2fbzyy6Pf3Q8jsAqAjpb5sa273sQ3dvQjGMQoJyPW665W7qpQIj2nVkAku
64xgbTuUroxJAunIsYile/V6YpwlkI4G8MBMSWaEZPUWC6Nq0ISe4mu/bkbXlXUT3g/n3Kvhtfai
UhJeiTaccCowxkv86JDEEMJba7ZuCMEbO+qF+lNEcCPccz/GQSC/lmTpFc4rlDRSoiNdASYFkvJz
pyle1HIuWlmJV1j40oQNh8Jex+yBV7OuCXgcMxV3U/e6Kt8VpN5ubX9irdBoPz+DMyzEO2SlrU03
U2VHAr35JFPfIBB3E9ymj2ulQZcm/UkwNKiMmnIfVGWHl4jVTu7wqP8ZBRDlC555lBxmD670EXLN
z2+cThjVg9HNfPagF+ccIQiEzZ8YJ4dFgW9KL2aJMRd+JeVcAaQcVAS6Koj9ZFns9X5td27R+Mnj
vzx1MdtG7c8psGcCdTSW84I9oj2nzSW4OHwDu4tEXCWseJzHOIYFlOotXlq/gkxrRHvr700AgtCf
imf3sVut4g6sxMNcUNoR0gqQlQgc+pIcvjYFZllnZGMoJJxG8v6KGXSTlSR7PsgmNUM/Z+voogB0
CBWNynZFuCa3Q7sIfs4fPR9h1T1h8ms+kkpiGjbUVUPZ+SV4XQ6eNOTisSkfzwAhKqzVXmzF8Ecd
e15Y1iWIC/lB5XEtg3HJuyLoK4WLS5IkSENN+Zk6zieTcrlC8jusYgPI012A6aTPjNTVU+S8lO5i
GMUUT+Lp5RaOlzuQSPWTB0AHniGUWujZ01PE1Qya38jGX/ck68IssUzcnNlE+Ko45X2nVgfqlAfi
3BR9XpVbN10eLFRTctx6RBtdargmh2uZXpprgE2GIEV2TUDkSm4YGa+Ow9Xo3eKl+w6xU6Vv20Dz
0uX2OCKUkxNN3qHXiwyUQm3MG2UIOg14jHKXKmlmev8MvwOKz/SCMJuCcuNLr6RcylxZbnwFaytd
Bai5QUj3SHmfEzz1EjbuTUzS6rwhGFt2dcqKGf4lpKHGJI9H9UujdSyVEyRGATi2F16x2Ut2Cp0K
0hK+Q7bYuEu3xjSWqnLCJo6ich+8y09AUPkmSentoBzlsJxfSI+Oq8891KGXsav9rMSnvUSIDHxw
6viR5BR1XmburRbuRmTFE42NtxwstoSbm7uSJB34pA45lsHbnXxn6G2GmR7ZGhQlkYMnao+aQ8YG
QgJaK40FfGiiE0a/ZkJvKO11GhAGYqhnlqAbDolGLvaGBpW6SyOktLSYpgFq8Z+RAdhnEZvW5ici
eNwT1dBZV1l53uMc2c2H/STyLWXW2W129keiPu6pLonmmYt9ybl78bIXdR4q8Y4GYCMoF67Nu8U4
+y85v4ZG/0Aw+ZaSU8pF99z7noEUb74tu8E8w3QPTU1siSC19O114ciDAEUWDDhnfVwz3HVHBtSe
mUAib/Hir5GOXTw73cy57L0b+GGt/k6lXLDPSLCWCQdk/jW4ydwHekP38jWmDHEOBKWflQFy8eBC
ktVmq77i1+G0XJ02WiLwcvGkVKcKgZJvDUnZ0nYzLo5ga4OdeiTG4JswUOOCItMORydg5OBVPyOw
/DaS90xyEvUyPivAvluSnE8B2epdbn6B5j30fuQcqckY5l7Ts9SFc5FlLSXMi8O2txmjI8qV8mSc
0eJgzcll7yKWCYAYpYABjjzzFnDFEF/SXfqAPS7xVHSlHAFjMgZBoo3aCuRugf3TjTBdTiT7Wxtg
aWpnCtztC/ac09aOzzdOVcfQh03eXQK4h5wYQeOYKG/TqfIxB+BVTBxE96iDAeLADC1017lEJEqf
r+uRTGW986CHTs/8tvdOIpgandcsQZn3V64hF4xsFQlZvyjFyu3HxuEur00OAmf7uWu234Lh2ele
/8h+RBcpUeuEr07w1Xt5Ex7ppiIkuKP/DT+bNCRW/aDo6QFxlIKsn+CYlr0MgzXs1oU4CBWMx5mq
ob/ru8YB2esm2UkP5mJnhJYrSfdCcy+7aNLEJOgAFCf6jOAj+yUvkjrGVoyPZTd9vDs78VLqbyE/
3+HivgTOIbREGCvaHmOryyq3Rf7JMgYjuQogIkESAe/6FbeOGQSOBGTWv7SAaYfv9vTOWcgdG1Yi
TAznpv5GrLOUaUF16Zz7guyzqxEDrTDp/rXpyPLrFuzfJT9sS1ourgJKuXlCxWLoAvkQ1bytP4GI
+YlKTECiEkGzmfVHfqg0gFv5W+8FViP7e079JXYidxUhCiORNW/XqkEdTleDfdGx+CcIW2yjLvvF
ze7E83hq9A3DP8myzj3tzv4BnnPtqtPueLF9bCb9s5fqceohnW/FlXSSrgVQpm4cnWB1zOxvJIrH
SzBDGTyM+otq4zlQt7dl141aAZcMLE8hag9XQDqB02NmTmGUhOgwpNZBabS7GxNFTAui79apTlOw
8Tpm9MdUcvulqNkf+RsoGD5iR5e+o/2waaWrGwrvzNMsDlbDy/esCqZDulC7SkUY3PDEx3tJUmdu
eRAMLuQyFoj0qbEUflv0emNuig+bFGq99TysURrM5mpnweWRBDYu31O44TldVilX8zItD5AXGAG1
rkGga9HNQk6+gj0ORgQW3wftEzRVt2R4L5ZWgv+G8PadlmooAl4osetideB/YUos9WvLEOXPLGUP
4rt0FCj/OENg4lVbYjGsbAWhafwDuK6g074OyxtrhfW3TtQFNr+D7ie0R1Lh+xsg5pA9jIsWGRnq
LcghY0V+ayy6dJD3KXGTVvR6mVpiW1ThHxDbXE/H+ddxiI21TrulArX+xtYZig8YVGqYDFBbJEoc
Kyh6a0+CeaYR3KQ+AQ3UU7UKJGrx7DO9qrJzDQ04o79oIuHhVNcncCwE/KUC/Sm7ku5zS0Y/qUmu
lGjaWfra3I/5sqcADC7QI+8nKDCLWdNDvWeAXpxqYn65bsPuKwOwPAIOygOR0aPLXK0Wh4dHeAfl
45IQTF5OlUSB/+gqH9pNm7Q8Weme2YlFQn+YeKjXmWNwwPaE6+cu4mq5AtCvI2/NABmTL+EjxCp2
z3Gndejtn3tIWz/YbbIGoqLQzrLA/wqtSNPmpUE0KCaVhHrlQyzFfTkhn5Ngwnb18r4r9XgRKwx4
fRJ91Zgvv2HFbCPPcOq0KLLXYMrsKMP3XCq6K+Ytk/r24dZ9PvdWbom/QoNWI3IjLaeyEs4xZCMy
ckxMMvwg4b4lgd//5EpbWaTdQGLlgk+QxCcptKG8SATuOeHPdIYOoXh7YhJdwA3TaOJ158U5xsFA
z1EEu2Ee6s8ZeIRiDt3IZ0uydTPgn5xcSdEJygurJ+CcdUuG2l6KrF9MBpm+yi1CtX3TH1oSq2ON
h50C/co2vMB5cJxcDBR7LW3j2jRqDlGcSPnDXkOPUcdMGscIdlXJfwRcUzuVCe8r6knsqu54SqPW
4akhCq7HbK93VWA8ZpKLcxt/J2+Jaegx+l8TZi1XkC7Ix4/rkATjxcCzHdX9joxI8H3RRVjVSZiy
GqUVAweRvGXUu/JF1q8c+WqjMLFlUacmMtWaerVjjMksOHVsH26TYqO+eitT1zcdFqkPiGhhvTAG
BYC7gz2BbNNNVrpevlGviGMomXRU810THOmUhLFUeryT6pO/tbKC2Muau4TTlrsNTjlfuToc9x7/
j0WbTffa7zyBauUzxpHcyoOp5DUFxgFJ/+WPs6YFwLo+8V9QRIwYAtC8l+jnzsJB5hQUyNmpAWgH
u+XDk6QPgAyyk/TJZsICzyOgCKDh/8jGTMY/25kOMrBUWfhNFTLMucbbowQ4ZNKI9ZAqRSiFpg8S
8D3MqU8FRLqFN62F+3Zzd1q4RU6qXEmwp3GwHhnGrSPiy97g8nP2IeLyiPkjzGk9Jz2BODRLFxsH
X/9OGBmCC8ItDzMEgApn0vrUaBm1JE85uc/l+zDN0ozXzg/ODt6tJBThROYVhmr66MZU7wvFvVa4
yqnCgtAWNfdJsS04U2NpTC7MRBgtz3CuvAsnMUIEGK44Uq8nSPTbodsiFp8BjiMbiSzgCvysdQy9
UZJwD9wniTxiuI3/Qf+EQh3MUrbFONvoQvMRJo47Iv5u64HC05V13FXTQKoXTd11TDDCx3nIWdDl
EWPwcYZsGixS+vP2kF2z3n+A/RokIzA8AY1MeCiuGN584voMYGSSJxFfX4tH+rmM9YopWFc8qScS
F6blhBOZhX2WsmtHMt1Vm51a/i/Cuq7trP0/lKSO/rxyOJ88MT14c2Ka1hJ3qH4E/cZZeMKoOuLv
XcS39e0gqXZIPBAtz10VFcDsShmt2ufAs+rr0KRAi/5B80e0tQK1grYdrCvV4hgyyS7r4fT7pJTR
NCY1JRjc5ksd8zm+4IFCpUF7ffwrkicBPOPUn+hTGdAS8gvKzxyDRj5azXpjhN6lyTnVII6UXBjl
pM3jPqvnFE1V0jeb0tl7SIcfvayohxFgRIcwqG1GlUdkHXnM5n2saJ6kVap2y17VPc806R0DUxjA
tedic7tS5Gg9Dxs+HoLdycWZLDYUXuOmgWE4MXiLAd+SsNrmP7vU5KHJ3LcgCtUBiv9cBcrlba0D
NPmDxLjvsamtZ2RzLlTOf+40Ae+uRcBA2d0WyadwnIBAuG1PCqqqR/tR902mo77HEkySZN9lnQM4
Tatt7uIpKLfEUUQWIlKEopBqT46knMRxNG7FusA9tv1tBHGqsmQt1OwfEUU8kB7A/xp8ZiR5rVdj
9meS9Dy15ayq44gGFb1BcaW6p8IBwXWhVl++oYfVdUgPh2BA0l8/XsAooznmAQL6mQgNgjLCRNU5
dut8BhHF1hPtqWgU72GAg8t/qxU0PGBRXNJ6OLA1tgoUJJlTJhWZj/UMCz0Mifl/hJDuRPeu7hx8
20XKYfyYuEbO8tsYOy08xyoSuwLDLaMwSob4NicaFBHHf3K1lM3BKebctl5m100NxTrNGyu7rJEt
aHBgjD1Zf9QsA0n2ZYej0qKnnW2XCR5iC4jx0QRLQpuKA3BnJJxSmka55qYh3aepIHx9W1QVFNGu
RIBO1FIOrk4kT0v6XyyJJWGdSM3SdWiPw0cCM3y9J1/Fu0eEPxeJsI20qMgoGNswTR39i1CaPxvN
PzqOnUoDbeoANToTf7pFOdlALkb5CvV+oFe4R6vZb94JIcnuCpFpcDn1ZqpE4Ihga7q5iAenslkF
QZ4IPEXBOeFHcwC8+4pFJhmaW6HxPom7KGXDRRkpTFO0MUQ25jmzhOo3f79vc1aaoChe6Om7Fbyg
p2ZhKrbnXt/q/xdfzvI77I8atZ/T5h9XscqYu7zI6ty7yBMzdWrcSOaGoQEDiFz64MiRrFpNQSlu
qUuzqKVJOdu+VFoGRzJQK4bEhaTnUrxtqzQKbp0I0ObT/o+Qu/PNEpcGQ8W5DniCRF9pSWoC2zUt
Et/fEpVxHSsTdp5nnQvCDE05zS+QaRffiQhJ7FS+GPutTq+F6O2TmISjGSj5ohODTmxsKGAUP3p6
vp1IrSND54aLOGJIlbgJr0sC6R7PtVWg/MBG+bVl0NjaxLZSWjtTAiOMcPnpZxykSyDWcNjRWktx
LOEx+2d4k2LrhDxI7+OP5jSAyF2zmmIn8eOCM3mgbU0Wj+Hy2JvzsLg3SERTtzIN9tes8x4MIcat
vE+cjoT/sOQQ5Op5G0eoJIyi8XkUghTMKnwJSefvGPPBIlyw7dhCaVD0oLfcd1r8esDB0PChTOYJ
0lGxeivvLDG2WfUw3sOD9cOh0l/Oppaz8u+cpkVit/+epC4ThppLm89NPQKjAKO3ucWj/IeSjCPa
jZVVwa+mDHRsGVh/Aig+3LWkqxer8eARW+kuvqikgGO/ggdc8uRFVye8QZItnsz8evwvc7nJ8vOS
vRw/WLfYxWWsdkhTUTUjqDnjfR/U0woRjZhsAtbFmzMIDKDQWAZwX0BeirknVRDCZk+MUmmrlaZi
FQuDNYylQJrSKMyuR1uQMaBQNRLVhnxGlA6V462TPxwlMBy0AmKSwGLJWdbEisq/9hm5/DGb/J7B
o0MbSwNYXokNqmb3NfJyCDrAPAzVE4/4Gfc129osxi5nK8YIoPEbrTsw/Tcmac0sau717sn9J52M
3a/ocrz23veAuTQZ6Dt8diEJD1HsKKru9M6oI3F828wzMxR2fdCQ4g0AxBWkteMvii+S+XxKh4Af
cdBuvWVS8zCYgmnGDGHgkkMp+RS8wUuZ59K+UakuPEe/V8kjq9yKr4bgMLoonC89MbFfGNfXV44V
BMNI+C4/dGKEztX6Q/V9FCOqR9QVNaIfzsHFafEbqRNhBWJxhyBtqsXeGFSzvuVcgh40Z52/ttmM
zixgbGAT42eC2uUAhrL1EdDP90jpew/MY9sFD41UJ9vI/XMchXvME9KvUaZH1tnAX4+vtZUqWNJ2
2jsqndZwZMPeAGAhgQn2Uh3G2SeHKLdAyRheojzBXEYM7lxl57YCcrX1TB3hsnpYuFhq4XcWXwzE
yPfQlHswhoepbsBftIhY0/MaT3KokrBXRv5BxyhIx3H+DRMo4FT0sG+gisVa2aARIz2Z17m1cqRh
82lk+B9aJTFx3FbKhITd5wgy576vvZ/cxTHDlMQBQkTORmxgiprTWIx4v29lltRvQcrrhBIhyt9M
Z6EMXFI7Ba79ngkitwfGM0h7YCgGffU5UQY++zWP9tIrHF3DtUHayMMXe2hzeCiC1yrW3ytjc8ED
7DbtaOBMV1QQzNNtdgmIQQ5wjK1OSgo4T5SquxtgTAnoYbfUo+S2IkDqzC6Csm4/dAhW0WSJq4Rp
sq1Ojs+cNiOIRPuso3dbw7vEqXc9x4h3Db3sl/xGK7Os3aE6Gmp+Gm+RktFzScdNrNS3M1dEi1/L
2klQearTUfeMmCCyQPFtx+h6dgJbcAaCgqeHZHModUCgvvlbSRjjWvF2yNa/aG1L6JyX8MIRy+TI
CPonRtEgPS6qMICD3FMm7sCrs2BE65R+A3/cMYlSdVIDzO0MJVEccPaFJ62gAh/SLCAIv3IKlz94
CH8K4L+FediX5Pc2CHOgyWDXjRqMmJB720SDyMc8vtYaF50tpK8VL7b+BrNCW4tVRvrncYILtSpD
9MdDsqx2BIgS7m8Q8qOKIwYcC5Ddotg6ViVhWQLdlpkHMjQDXPwCXYoym6I4U9/TfAD5CAtWsAN2
E0uB3Z6yQ4IeD9Nj9nL7KlCk857KPWE230QghHFoYU9nVq0RCwjIQq/kQukfiwds1MhGuSBi2yHZ
JMo63a1vKyLZZUs8nf8Biv37L5Ze55D1DTxslVgY/lB8T2OuFqKvyKzVwbq7nCy9mhWPwQFfzOgx
SZeY+fK8ctiZu31GAtjVIGXoEx/7USmKCdtQfLrT+ccWwtJjQljIwh1yJOxeXfXaI931pSpkp8Hd
cFY0BetuO8XIR/bWS1QuYHEonct1ZBJjLknL+a3m+ip8U3Po4g9cwopjI6sy2VXcvv4jJR2LWpN8
ml24rzvgpLXzIj8/QwGSKSDCKlqzMjFPK7IMTEsEjcNYrksn7uOe9cPCs7VSsbbyf+7cl4ar8WR6
UEr4GI4thdSKX3PxOVMNgTTk2uAnYjwL7E2VmtyS9rMeqART8cIIvalSaqMn6/OjjdK6HOcT3dlm
+nEyjyJPk6NeBDLyJBASxaPjsZp9AmcF4/HsEAKouGTTR//O3BFZQAhRfahYjZlv3r2Em7cG1le9
mcE8Gwsq7YPSmVVs4keX9VdpgoSN3p5VYC8nRiJXkoZV5537em+wt22h2328gMSaaPknZNJh/GN5
3eONAnAoqJNY4tZlyEEH35yrBPAiuEKLzzkC/FCcDFU0xddKFk///GRJxEqlUNnve1IJq7VmqLh/
uxgwP/fa6AmbkGcoITnRbAJ1JH4iqcSJ28u4kkYNyw5sUkrZJQ8u4XyGAH1JphvSrBk8M0Y5AtUl
vYx9VSB/OvNtYpNNHOm8Qcqq5Mt1+fmgoMxGHQBl3AJ3Q/F/OmkAsLcr5xLcO1aUhuomsGRMUTGh
vtqUgu4T2pMAoCtPf5vd3AzmpfIzD0qM5gC9toV4NAMVcGkL28bxOKrq+Fi7uZ6iSxpHuurhsC/1
SqeRRj/YvIomIMcB/YXv7w6j0gudhDUVE7u7g92i6eiC7rFuhHsNpA6mPxeluk6grFo3Pt1tAMN4
xGMxG7rndX/vUNPaSRHjx8VD6nO7TOeRiPP8uIVxql2Px3cjMO7Z+lkewYIih1mxPEAL4Mo9Gj7U
NYQiTBO1wqRH7Ol3CVFsI9L+TQzgbgXAE1RrVenxcH10QOBuXByxMjcXyK31GSeGRZYlQhkuy6lO
1Q/ffe0lrOcPcAC0rrXhYUUcZi3u8NxtwFzBI4hExjd+86Q+V7aMussKMAUHgw3h6C/HqFf7iarq
UF4+f3FVEfLWRY4britioGkWfuuh8r45w5dsG0JRAdD/HIqpqhUEjsGZAZECWhjB41jWNBZk0LHt
VEKrOnu19IPL77wC9snHbs9yaUIdg3MPtoFNzEtvxgUjCnC8RDchWbERpNxS+YILzbwEKANHcReA
umSsQ8QszVUabkqWj5iviM481xRozH8EAz69vp7f8pKGt8koUi1C+jzGImLOfLn0CDiMJZF2CpiK
5xnjJoVKHc5e3zaThKzIIdA95ZinsusFtzs1FZy5Sjq++lJ8FTenukSAQOfpp2TahBbKi0j2JlPY
YXcsj9slvpAazOubK+M2krOz0X5M3XSNCBxtA9mqRkhVPwh4fC3e4oC5ag3wfK5EqGTfwZMylE/R
IERCxRNc1CAlNCgGNuYAEqY0+8CgLarBwtcxcAL/Uh66R8bgIqBKOshhei5LCEe+Ok9QyPqz83oz
b1W0oVhQeRKpyaaKF4Z8R7Et6gJvYByL5aEjAwOB+3uo1RDyWpmvIWefmUHQrWPYXpq/mZR4rqCB
KIPdZ3iStgVsmlWTA9wUXIvKhcI7uAZzXh/MKm8TFMH3dZsn2ZC/DUF5+JGSSwgqmUmpuT8wSTAW
VrkqDk/pSBlT0hJsM0svbs0FTJQ1FeaZLcNjGC6ELqFUJJnBL3JuBkG4hS6502XJnut45gcdP0iN
ze9KN9e9Hzv1pmD0g/UGImd9iK/SoY050gkm8JphitUXfskXhUKT9XktJYwN58wluK2QnXee+7c8
/eKXzzuRlkGnjfRwMEHKJtZX2TikVNmcJ2Q1dOQdLGCIB3XntdLSvaHHN/acGJX0IEl1MjYppiMz
ke4rmXBz4JaL1uZ9DkAl8Lr+/mVWSpoLLZIF5HpwzN5Yzb18ms2IUbX7dt9e3kClTc7XL43fnyt9
6u0F9NGiS6uhVxXYdNKQnmwvA7g2rtPA3oLnm65ZCHzqGaa9aUSqp6O+el/83zDjE/YESLcUb1VD
fAQxSoUcuCXiOg8BH/C94OQKEt8JEfXNp4daZO+M94p6jSCTKzqisB6CRS5Nglld0rMmII3BQxIo
q55hMlQVJuNpiTaVMKS80mwIJPpGh8rrb3uvAtmVxTTUlSuyKmyx3GvNuFKO6ha8Ev+vQHwot9yq
U6xAcKxQjgwMvPRMhPudy1bFuK1JoZZnedQCsExuXVtMrSN9NFgmWylV2kn0A7galqf6VhBAbfcS
wPlP9eDgLK9qd6kbXh7b6URoyR/FT56+SgDAmV3WL6EH20YZ+BKjw0TUC58YVWNz+q6MBqkdaCap
k0QPExXa6FYFCkQR0gNXt+EaRh2llAbtpRhJNohTlFJL93r1CLDS6QCpsQqgtOG8ifW7zgTuwSkI
XZ9yJ7q0bItsbkAy1ojo9PwKAWQDj1BYR4bNmypgUVaF5jzDIEIc9djy7g2z5AprH1fTuHXzapX0
42geVUbwzHFDNlpq6wDq2XxX+/o2vjyC95An5yZqPLH/Z5SVSCMwlQ3gi2cboGiboklHRMHCGYr9
/pTtb0/gwCWz/Q/8I75xURql7Qu/UbGy5c0Qy9O027ewAhOGjvRtreiHkXQ7KPee0qUqAXgsDYzM
vh0OCcAyS7Jg1lgEGWWxeS9yIKrhRb/Wv3Rda60YflZ8TRr+5bE7NO7a3mDX1+Y/OFXSrB5w1qyn
F6nRt9QtljegpqlnoH/fqQcV+PK/UBJJoKCluglLjobN/ABOdz4W0RSNC9RFeygTmvpOGD+A7IH5
bJN+WCmpLmKBLc6nOZIVveeECUMlvpY4rV2u8iN898+lNk3miGjbjAYD4p7TxmdCEzcrOxR4kwNG
MYEFr6E9iZixEY/Xt4dvNYlAdBUkwlJ7nQBLcHgX1Gy2NxLh0DSZCFBLKQ0IF9XRd7OL2UhotHtJ
QEbLLbw3Fe2sRBQbjkTShvoajwfAsOK+cnToQHVkwcqUaR219ETfOI9zf51scOsBm8Pd9B3PCNLX
nryFjj3J/sf6rG5l8NX1YS2oHmaNCqWVaSb2d5GWgUyd0egewPe0N1EqaDBXmnn1z3QVIUp9c4ix
vplRGi2RhiZTzgHX28NuimgDCG3dA+PiepmAJyOkjdpROqe56q+JMHopp0KaIEJg2SDZqUs6vgcn
iwAP8XcRcQyZvRXimtR6Y/sLz8MHo4QAp9+kCnIzVgh6A/USmDJQERXdLgNmKKQbIkAnFLdNMZ9q
3z8pTyad4MLxMrIBuGgUxGA8JHn908YC9MLtA7OLmt/YBHhC6CXzMZC4sitWSc8GLW09d+HQCBoa
6wBoELXUXgp5HXIbcGhqO0ZNrSnSrGDXu93f4Ch9FzvqepTc6dxRoP7aF7SVRdy/ZdBZWbm0ZSd2
d3GHrgPGqnwBh0djNoW+qH8AiuQ1YwW+kKdd/oHOqquAIJuY63mMD9GPOi+DBOUEM1f80S9aD2Qa
MkVjp3jObzQ5llijQsuW+KV4euViGPeAanfVYEsUPCYcxUx8r6WJQLVOtZxRzlzsBt3yTjxHV+Y/
uuEuizjeiJhPPqjdF25+EWKDHA/8uUh6bdRKN19F5odVGBSOehgy5ylCuEXt58ptu+/IyXOUF5UV
LTTS4yMZz2Apv72rPS5uiEblYdlEBC+wDHqPPQ51tYJDRS6QpUwc5xhiq0JCake0/A6VkyjX9pET
KVW3V21OIngkipl2IHYsfRxgldllmkjIyyGMVj14UqyYuQlgr2dPVX6zqlf3KtoXNQwoGvZTs0c6
Po5+1mvbnH+EAWRZfDIFQB4jpLbxdE6TiyAJmiUUD7YdEf5v7ftrmdVyOmog409OyCeGsYUD0pLd
dmqSZ4df8ZuPBJ5zkBMlQ3feB3UGaCiwsL9QFCkbIqOuAWXa8H7O5Wr8jFeLToWsaUxul6A04lFX
bzgIUtyC41r4gbQF8BcUjuGMZLmuRG6i9azCN2AY2bXoO8MhQIAnDPUuLlVfMKDojJ6NQx29wYT8
9WbO7apI4iKo+lxIdH4dK0Nzxu9tYaO5tF2C6VpyJqR5zbwjzc+Z4WZQwc0vipQtm+q3orDfCg6n
rZY8byNG+K82lytX/m5vCEfN4/1/g8U6RvL6A5dljT8EXVhrM099ZKHegDK1bEp34AUbT9twIayu
JgSUwBbIEpvpnLax5aYm1lAPmUcO/p7x7ijU8x9qMwIxbrB1xZWcdhdDPWqZHOx+5ppqb2wwiM3+
Elh4tGIcQEsIKqaJ/QCxY2O6EBZ9RFfze27RrvwjJ0s3BkZxaZUoStjOSItI//4lPwPweIj7wcKv
mpqFYuxU7PZu8iwu67iT89Q/sQRPIuFcy++erUfbaInJkXZTDzlEydwippM8CMoi6i+WyVd8nU4D
DjIZjVSKxFmEi1QfAsPqcCLf7P1jnUG9U4r9Ys36+IUFmIMhF69nPDJS2EZC1V4Gi5BzsmeXPbIp
u6e5K5RGrR8KRguDNI9/EWVsamLUAe690Va8et1gd/HyIy8raz2GKj6+pHPxJgylI/8VSJ277HUa
62fbQwBcJ6Sbz0VJF2IHCkAnDB8Si5wrSr/ZNvUlgZnINoKnTPbRSdEA+kD2csD9D0XNX1FcGlhO
kx4NuhwQQlFAg0pZogLUpcnEz83MWdA5/CXtNn41vyxIBOx5qUybuOya9Wl0Ne4MKLCBwkyyZDQb
SgmO2m0lYkwsSeZXiPcOwI5YN0NGPAhdoP/kdaaYbti4d7jsG1aLxsPTlp5ka7LglDoty+Te4oNK
Z4JWim07Tq/SLERMO3Q8WTZmGl87eMe2HHkY6P5rHcwQwJ8FlBnYuNOiJlph3Q4jg6UNZ1T8Ot15
VqlEdHSafcr6izQ+BiFGsg/++0I9HPnWqmQ1T/0qiQ8bfwtBC6nUrflKGPk7qA7sMHY2LIFths2Q
nkQXFPinKHnK7NNZ0Ykao/NnCVmhMtjfUkd8tQg4Qzyrzgx6fXqlNJhLRkSzEiIWf1NczxMINPB3
D++G+g7vTkSW97ycwyCV6hhRTiAtxejQzyKEUb6FPHGtOMZHOaQczoFnNe5xDm9Rb3VgDbGibSzT
cZCBhsLMaT08OR+/hDRwEKOyLpWBfzsXLd8TXJVSuz97ufYbJtIBp4ZTfXXjLy2X6diZnp748a9w
4y7S+wIRr8rCPgdBuotRBJ0QlkE/Aj2y78Fanpp90mSBQhQZTBxqJSCwW0UssANn7JYTRpdRQkxM
9QuEo9oxn1hhGyg67DjI8ofZBcj3hL/s8kyRwUISKsXAc9Jvq+dX0bxAjZHNDTecPAzJyIKRozLg
QFBhhInRdZm5nE2rZPbRjLJgJM5rqRsKAP6XBvJxLtB3LzykDFFbjTr9yLbp+9xRiGZlDgcjNL+j
GhMnxZd7TQv5EJXluElAU0JADxHP/Hu/1HoYS911mM5AL/CDlrRvlJyf3qRJWBRhxdhP/CPIncDr
z0pRIu55lY1MNvkEW3UuERLjcjzvBeRIMzOExk8RCoG5l0455EzN7YILOhiblOvskiVlbCdZwR1e
HEGtN842y/l69dnZMU9QG9oBhPzohwtidcEhEULjF0/vjUESI80m+EcB5GiG1HS3le3TYwvxCCqh
juMKk5j8WTYCUvYDCf5U6d/TzEwvh5rfAGo+hisC1tfs6ovcoVhbT+VK7ALZB4jJzf9gqUTow/D5
cugrPAzGeOt0XkN5z9tuCV7PeeCpmEztOTZU0kY06z/9ru4KOutq6gNuirVDNqaWtRFh7TjrxaN4
/mUN1QzAQzTpsLFX08mF+fhTIfFCd4UScAwzi8k1aLByWJz8jIRY675+h7G5/ghpQiLh9yDhKzZf
y/X6jWoM45r44XRYonPHg2xABdc2yS0KO8hx+96efV1JODJI7V/jk9dZ6ysCou5G7S6pTqSjv/VQ
amYXssTSQm+Fi6HsDDjJXbbch7E7R8BiOQRshekIskQ6xm1YA50SztkjLG7yNRX2OEoiF30EdJ/L
/9QUxywCGz6qahPHyooMq4e9uFSAxwlhSQ3O+NzZHtXUKOZDaOvs57Dqq90VphLwaUFliAiTc6h8
1LVvC0NkZwXw7hJo1IK3rvOUUYrlv+PG+zmCJqFR1VwHXAxeROxYeR9qMZ3f9sfEs8kDhFUE/phg
x4dfYDoKn7eSZXAEGzroQuEJIld0jw69ED7pn5AjNH+CTTsoIahtWh5wbyq+Fi2VW6Ok6mhcDp58
JznGmYPMt3nmQWyFGQRLX+xsG8i5iMiug+QA+xEWPiu/gyoGrRx79ou5x/97ZGyp/E9yWx2AMOAq
A2lmc7PziZo3seWmqYITmXhRQPty91N279c0iMzHRkU49xEI7ZplZ4c6PWppCkK80DTDJD+110cI
ozWcok+iLHoyloGqq6K0xAqzfkJNFZPDB8bgdIzUxI88+RsY4e6u7cKgdI1pfN+RQXVsgqtpM7u+
cDKA5Drn9PQr0+QQfZ2ptMggOZBblep/3yKwdrhmilmOWKX2bjD3fTjJFUWGvGBpF7cfLgqF0VR3
BK89xqdDLWY7Yk0netZ0WXiYVVs3sonScIqLrl30wBHOepovbO0XrflDejhi0mkzg4KLM0hbw8cO
IhuVdsbTzgD0Sm1AIGKsdCOh5kLhUdsiAhwYqRWkB8fg0zCh3ey4eGSOMMpQxtz4u8LUTerZbHXg
GI+cukN1XTghcXvuRJbamky+Lfv//Sk4z2o+31NghbF6JthTzDY94vD1JMgI9hgN57DkU212FVQB
ELUcLDBkfctxmp/36U8ioXYfQ3Si2TmDTA34Ctxgtxofjqlw9F9l1BF8P7abwtxpWEQjQrUbn6q0
TrwINQUcoNWgrEiJ4e4W/dLCYr+mVxGre4rto32f83kJlNpuRaplS5b2rvtx/Z9raHHO4+moWkvk
dPwpxBQEtR+ABzQRi8PMszzpfHPuH9WjU6JRNjW/EbCs//1+++1rFNCx7Io+HiEcLZdVSEcScJ+p
LU1Vj4Z+0pAIzQLI2BDzTHtp3dVY16XKsK2X1mBZrS6oc7Ucha/0aTBl5R43s6Z3FVCB4fRMQqiB
aUznvBYeSl7nIrG66mtszlb1tui5/6u2/YVVBSZ8y0THA2DBL/KViuO2MlGjhKPOkP0SuQGf2pPZ
dK50yTgjEaKuec3Zd8c2n752GvQfn8nzj10dvuUkbHaHMZslYxlGAnwBHNOJ7iv0dJwlEFSsVGaK
Db9MAXX0XEdsrobiPZ7qZCueca3ob5uqQNsLkvkJnQ9QnR+iFIVKtw+PDBAS+2fG/esNTxbRTzxS
gWIiw47J4tLfarzUUfFTllEUsz3mJ+SF7OaKF8H5Y7dkCTR37joXlVT/2AlJ5PZfKtDIBpy1Shj7
z1oBYsgeRXp0ifaQrq3quKwa7RvppAdhVUce0zvBmLkiUCgJ/Q4rKKJkWMRBlGvfQ0jBmsmKG4hV
exyRAd+XdVp9wh0eA5Xcdvs3nd7T8RVvk/IfgutgL78fVPZUMVRtn+UTKe3A1fePZciye60mpu2g
OMWMkRdt8VwwZQrqWPJ9Tr8ZEw4VvYLy8+hYgn80ukDDRxEHVhh2nds44ZMEEc9Aw4ECCaSVjLc1
Yzq33caXR44SjCRob+4btdtTJcMBhFlkDHJ3Quk+eBCTpbVze0Af3Apu3/JZI47lA+3iDDJy8cyc
EPD83vMGEIPWHB5ouQJoDyEEU7Ug/Fg5jsbwRP2S9rvU7Ne0MuPWWxRVWGzjMKSxYqO70EnOWuv3
P67yHdPqTZQfd/1nJ2K7zbzc/qf3nCe1Ub7Be2O6RRaEvCf4QfCAttq056NRn0TjVVHE+ugqbNRL
Afrf0bvb3z8Mp1l/7Y7MSFjGFBX++M/UWAFkx1aYvVl7IBJzha/AVZCFf6I59e+H1QZSH4Y0kihx
iX/KLXyXdUXhKUV4V0Zk0nmbQKVmGksGLDcgSo5Xc5NTTt7W+JMGuF944sobRzmlXHKwyESS4yLS
kBupDFJwOJjvGvrVt6UMnnqxf/G7RTDgKk3X93n0nBsOGHHyzgiGZhOCJnhfLGqMFTTX9WBSWY4O
z5A6iNeKlcmYW8fnZo9I6TtGGtTGv0u/9jsDN8xY0qk2/7Pq4/4QBqWS6dbLhD3lyrd3kyszQwV+
swvrw9eRSkDqtKgqO5DraaMBNH59Bvh6YHZ8knLCq+M+EViIS4hv9mk7gMRUnDl1QZUo0DhPkFC4
jB1IVUIQxjt/L5/pYpVpfNKV0L4bQ8PwW3+WhbbYslqZJh+ccJHhFl2df0ASmJA5Ov53xUC7jWg2
Y8dtVjl4Cgbh60/pS7kq5IQO5/gM1/lmtVHw6w/e/G4PQqKEwclbXvZgr24gxYvOVAx6fQdsjaqk
Nw3XRU8Yv1h/t9BSBNujFb40KEspvsuEK/oSWNa5hvNv3EN9xZiBOPkLij6+ZwVvsFWY22rHu3pZ
Fu9Ef1olHthgDGCmIwZGFDYOpgQ3GKCHaGJ0Rl05acUqc/OsfsS4uOBX7GltHK8LHwsn42eOKwIW
oM2505vgrGffTg4suTas1fKiuXEXDS6SLLNyzsYl+kHS5Lu6mlY5P57WVlIcDYUzC+bpU06cQN7i
nvPLFcppsGdHe3fhsIYm2053bv9pG7usRA3f6jQcFqW6biY6HIT4j6gU1fCYjKe+6lLOEpMvvMjC
q+6JkJGaBjOLzZwMOIOPOU1jC7XzQTddGNGzJ2SJlhkT+bbjeBeNTMRGLbK03XfEsYUmwqK/sTF4
4iF883KkCTsimCj5iiJvnuPyZxC6lPmcANYBlIlm+Il43aAYytcY5mfJ9+jRc0ou+pCEOrabCmk3
cSL5sxebqX046dDGR9wpDjQvPciB/cYiQ2PgsQLTW6s4v9yvkxEFf256PYdP0dz+IyLBAQemkCHi
pmxSCoxiIFkYBz8XClvCTfHJFQXH/ASqAEF/EQcuRKzsSfqX+awOUccGWZXf3KeoHby6L/Pi8T4k
3/pcr1E47HvgRkZh4f3mJODX0ECssPOPIbqaTAS42AHzjt1wBbh/ZrSqnBX8KfeOQN8E8c64WxdT
rNaYh2o7FGqfPAyaMlhgzHFpOUEF7jgP/3y1F8ptMcUcWnr8aFnfzDQVsVmVLED3mMX2fRugbmD5
cXtXeL4LRrxA8r41DaP1Gl6rN8YBzlP6hi/UhrMxSXK7DLPf1BX7T9R6HTvGrh2HPtW3CPneqD0c
nrWfH7hBWgMZdceCIQhErHtmWXeDEwY3NWR/WaluZxmYgasn7fAwNOv4KVvqflXVrSdpvDb38GcG
n4ogNGvmEfh0xUo5ez1vwu46W40cHS0UntK0X/Dp/Igxyewjsl0xiWZfVfY2NlaM6VlY8s7fsyYC
odVs7bHIYUZp0zlDEJx3KYG6axvSeHME26yU5xZUsyvFbH4hEwiM0gwGSf+UtlpVhyWozUcM5eYz
Eq3Xdfr+o93CKRpDUY84/3b/dM3mDMhQT6zwbQx6fYe0ExYb7eWBpPxO4xdtN1R6e1TZHVPvrYu1
ENK09sxXLiZGJBxnGCnlp+stCD+germ/ei1Nolv9KXKdyMY1ud0MOf0D/VlntWXlLSHBhTsMnema
AMY+Z1LLUKpOlMx4xl5LCQpZ418hfhoIQefDcrBs7jPraLtLIlutVpE7reRmk/6e9a7S7UlL3gKm
NPXvwbDJjSPJRR2BhaakSk3NTJ6kdTMaomKQTu+GUFw+l4yweOUxFXLnv8jL5n5NN2CiE99+pJ/5
PUOYf7TMTiLdgQwOs3xovAPDkaeLIVrVlGjSihghCuH3S08axm6iJkO+Uq/UjcCiFPBsLuk10pmK
2+6He4ucVZPz/boqXJBubNcNNLba99ZB60wcZrSlSwN4XfAXB3dbyqpiRJsVECiyncpdcb67qD2N
pBZj5oQijzqFg8TEGA4F4Wc7uBXlyzkXQ3mqaE8xK7P+FggyJ99CrikxpkarTqVZi22ni6euNT0P
bF+vSJclXxj2bvZ5xhq4bYQUhrOREIH4lJawWMxlP2gV6Yxm9yEAFyxfRE/o0a4T31I6pMikHO79
GGWhPi2Fn6fOrLQJlBR25uAE4WlFl10Y71MSOdIXUO1GBN4cFDCxRBVnldCGFbiBoUVLNcxfKZBf
QjIfjTHjbFU5s20oaoFl6B+s9WjhuqLTr37iilNKGTb4LrWtn8gVQcMiZpOcO389Wxow1QbuEFh9
8odIrf2H4ta8hVpaCQWYSg92N8FtbyXL9rJfzgEk64yGB+zBQF6TGrV44FrIKUaqe8ZJ/ufB932G
S1Cl10BOCE5iOgO/9lSLc3PgiE9fQQy0EZycWcg9b5cDR0rGwUuHq5Z50l299Gk16J4PU39NUD9E
QWb8pblNK0fj9p/r4sayEhnI9uNugDoMkWfc3FwM9lI3jeG016sD+UNE6VuScDrL7wRjokX9EdQZ
IG9H6pWTJ26oSbSNsyFahPy7qoLXGe8yadjmupIAZHHExzWZOfg6LsJhi6qYZLpHT7EPlxyTLO3W
LqiV1COdtevrzTMTVETmcSCfTkr7DwM92qDwL5v0mf1XBg3CqJ5s9anndXp20RpROwS9VmEgno07
G16g/0OVj9rTJxeXgY2N2Jvm6DyvGvg+XAUaYqVuouks+iBWOc+fh4EhIGUngqS45lH0MFxX8Qri
L4HF3bAzw7P2qwjFRbrYnRj6lGtihPjb7dr/AkFhh/ILaiBc8JxaiSK4miqQdHkYmCuQe3jr0BV2
ov9FSenEZ1/H3RBV7LUVLOZDDuOyROqMg8MwC9+7VJrdM9DrLXl2FXMWG8FWuDqaFaZGT0Kid5i3
7lquPI8KQjd1GFgZFm/cEt5H4z7ZSCQaQw3CARBsYya3GQDWXTK0wKK/NgUhulnW81crowXSAGOz
iTPuJt1MyPr2g7x+kcla5PfJlNF8fztjHAxGtkgHT49UZ/wPd5XYXjVTIlEqMf7hViomQ7B27wRa
Ta4aQ4vYpHviqkuiONdYdRJnCTmFVqCnKLE4vGLaWRFl1A0J44aTmb+KR9cQ4bVessddOrrdg9LD
wJNfcONvpQHS0suk5aEWfKBngDB7yWTDi+xIc00q2kZa6ax6PVtHksD2jby8RjtoswqtKj8cfXge
HjdHrkcoEIu8I5pDDYeowKE3UiPaBeC0UZOU6XV29Fv9ubZBSC6w5MDu6A9mDQGnGgbXsYijRMca
9GSATGjU9Vww5uL3IjbUIdKj7cNpOYNtg+oiQ/LzRpUK/6BVTRUg99XGl5qV7pWGTiTNl+9ecGn5
3lDDx0vrwvY1ey+bgk1kckz5CWAX/3ptA9i2txROLF1u481MTID9CkCH33RxF0LC5ZRtnyaHgt3I
wv2Xdel0wc7CYzmwYF0JGvFxzhNxys4DMu1pxrrVl0jD+viVCXKehO4J+ToNyM6BnAXQ5CGV7yST
CKHO/qP1G3brrmltli2kBgrJD6SzrzuV8kOPsNfvqWiVdzEWtY1wNBf2DiJaN9LIlPKej3FLYmqD
7CBtd0/IDdVi9a+qfHJCF8/acyOy5RAit8kTZyDo2X2je6U2+fW6E5Jik7uXwQianj/oAuo0YSxE
/3W1M8ZO2umGU74k/1N0bIPJifoaXbuchN7DiaF9Dd/PJoh/4utMHw8WcvriZYivurkoVa+sXGh+
dJCJpQal2N/mHubdWpRhzi2EYeQriZPhyVnvtavwAF1pAt0PostcqiWx6SKBiR883qomEotD7DfU
QtK6QPopstp+LKWQ3TiNXBBUTeZnS7lxQWFkGXM9ueeBMNT1QBMcVSP2KV7TxreeSRkJ7ITQqiBP
YZzKy41xMQ0pe3qFGRQXobmMOIFOyJ6/fFCgb+FD6FKfPtLY5RI1UYCORan+IadB1BNLTMsEAg3N
Ruz75wOG+TkoeXFqF5W5ks3vQkOPVkDDrNjpmjxdCcKfgwuiDPKV5kru0yFNcGK/v9nIKiMOY81q
DQ+QIK4yyanAn0BrZyGmwMliMJiIU/0Awbjhlwt2U682+2yZBJXufzIazWv/houOzjt49BqUItbv
UixlmOAVK+t7dscMn0xmnM/z7BsiJRvG7rTCcz1kf4diQM6pQOHx+x4JGjS1pwxGawGgDgQVCKaF
aQ5GfNgBfGZg8X7Mf+483rU/hvfwoUGhT2ZIo4++vkwcLeM/8FCoQvddS9tdP8sR/czlVbg+NXrP
nFq+S7fq2LwiRQhRsEaSgpZbXueJpwg64uTccBlB/QoAT3oXGz7fj215rqx0GAbPSLqMpDJCb1V5
3GMfeLs5+GSR3Kq+sDTx5Tts1Xqm7KK5HTE0er/6JXwp58MrHkbHsTSIjaucpGicI0r2tyKZcGFW
BK2C6al8eI64CnEK+lNGVGfSIYMNsjlBWEBnjs2SfrJGWP9jGKIV6JGaxSiqjXMW0aKVKr8Qpx0L
DrwIwYaVmLfcf7vXB1aAp/JjpDQnkWnYBRXa2rV8hF+nFWEdvvdHizDbv1oajAst639ktoF6+Z9+
WpdSYILX/R5UsSoDE+btQj1xIy0mOTYSK40pe5scUnmisbSLoeroqxrk7rGFOV2jRdF126efN9Ln
xZ4zctseoRp3LSYshOP/f5+lj6mwScIPSTNWlVz5uQ2Yh+DVRKu3wyOpGAtMsXhNORHpV3+ppZm6
YXyHd3jh+0YbxP0nrzPhhZ6eG2Xlee3lKFQAxZUHUDOwcvcnP5btQTRXhJqaGqN5YQAY56+uMDoo
G9UEkiDaGckk/c5R9MKS0dWY4j7dGt4fBBmMbnioC3uGq++uUXKnfkGZqKmg9aZAjtup64DHVZEW
FwZ2M/gY0635xKsMR3S4NhvW/0RgFfCE0A9pyP9/0VF5fYQgKutm+qNyZrP5+xISSC4Ch0elorxA
aQ+5IGDeqVOW4lo/qgu3wyb5Bos7wAIz9qxAfxext3972kyDfiEmbOqr8F0wpxAbd5XyvU0XGdHO
n4taDN21znK/DvWdKlEdOCGx/pBoDieX2mKMkqTfPEPHWEgvKDBUfnChPMAIMACJN1FyxURSQK3q
VRxR5mrnMkOj5kh9/ulKWfJOzZoVKzyiILz3MqJxmvG3SXN4VLUUgIaALDbw5B+/qe+2rRH1yLEw
5VMXy/RL7Ha2JIao7cX/v10zsHlybopHI90Gr59+I/NoxqZ70PLRsjYmv46o/e+ngNpQstykOpeE
2dWrToJcF+ylNYI/l0V3NUm+b6TZ3N3JT/qcr5h5/Nvhl57wCLyASGqfABzXNUdMYHKZRlZ/6fnn
FHEasr/VwjokWla39KZZ5rR1MBXQGW0CJ9uCljVMcDiExQ65KbO0jNnMC72bQBIA+MKAKYqTDJ6J
oTrHflrudQ4vR6GTFl1Bu4+2eXaCT6kPDtNLvhzdxB3Koc3oA1W70inIvjEfdYtDWt/TMDJr6nmx
o0t4OoCCdE/+vqUnDrYwNYlaSnfG1ILS6eYCwl9pyIQBx4FACUeDgRkWgCBVCq7x348QmJHXqnWV
LwM3m9H0h5G7oKH0R0fpP453Q6ITxm1c1W19GuBtgTFiHxhTFj6qVUvQ0uk5CXuMqDEG8scPjxAr
S74RC8j6L7P0PmZKOuRC+9Fs/dva7lkq23krddaS1/WAu0A6PxpQk9m0z0IIE188P1jHJSIcnfp7
W4X20tnjjk8YTHPsMzOempViNadZFz4ZQ9yoA2Cc572bppHj3/bLH4nIsx1deG/qQSPWJBXVIN9w
D8kNq+tYN6EQ+uk8u8O1stUy24jw2fA/BsDTxQMFv9KpeX/3srZrMoRFOCJ34sck52m9zm9AXHA4
6RW3OkjW6J8u0YQH+iYMlOnvDmkiB6HYmLtkvOToIM3aaLr/eHFHLDhIq3cpiliJXqnVLixQK+kk
KFCnHD8JguEG6Qs/UbBNb8lBIWiKQK4SzNxlZEsNQqrHHymkh06jPvByXseoRclW0vrabAj+O7vB
UMtApjw78rYKF59BS8G2sjvltaYegisz++jY8LvxqkWtT941yLU06eeUVUFpbC6gCXnpiCgESl+G
UAr3k06ogxuaUQR/m0lMkRXVRC8ZTiCVRn/Su5c8HVmV+SlKFs+zvN9TYTYAn2USOf+e+MxQBLIs
I5LYJZgoSaZp3KKrgehPCJWMT3pmeUCT+NJjagVNoPMEROvUOQEsl4FnCtj3+i8DMI9Al878PXiR
z85zbFaqERrzucSl3h0W2x/HLkpDxftFePudF5YG6ESyqIPg8483O8lZ3Gw1IdYoQbPuWBAvFJC8
X6weWCYvGWMpSereIVWyQ4rmSW5XGRNaW9IQz27Eu1rMEo7BSXqaEv/2z/Tye85Yr6JD7RtUU2uv
cj91UbJRt4f2hGfEkdlBnmLEhUkY76LcBHONaajTo9cnYV+mYoXoKx+S3oIMTJ8mxftWsxKDqRqg
cqe9UwlNzX++IIPLZ6EapskegssLQ8kPayGPcxaJ8SYdys5ubN7pZEFPSyGUkNWDMVeM3eJTHIcB
oRxV1k2kB+YAxX4kKXe8KDrcA1TGIDbI87trEAiO3pE0IiubcWy7FAhXjLJgz7GbFBRscrWH7d5K
pXfwIYila1Mf34E0BTVOU74HTpKPds7RX9a0qc+AxjdJ6kTyXg05NGYd9an/iEupCzIjjCHc5jsH
RTSWK35AQYG2IfsDW+5lst+oUOtHeIeV8qvEPgY3V+jGv0Upu8WuxNAHjNldsZ8Kdtgf81o8qlhQ
bYJJLf/bI42P3ah87KW/t0kaWFgszkzTWW4XNLzX229LcbOD+poNYtbxmTFl/uxoOBz8YZS6dcN7
cqdPSFtP/kaxEMdT6QGHfGD+Ngskn2U7sy9y33lrr4CUfeTU8j0W1LRYwtxPTsJ/+jxPitahuzkt
2A9xlRpeAHr4BpergdniBuFxCxpbN+A9rEBaCTK39qu/iwLxWh0hNXNCYgIP/G1UqlFSRNqJUQv5
ALPXotwkV7pexJTl+A3bpnuxqditNmmbP0fTyEHaG4wufy1CwSuxePB0y9/YnOV6NHw8Kkrinb6E
2o+3Zt6EP3mTyqApyyXf4/txOWqnoeRp5WuL4ZCnLu12RYCZh/al6whf6KWgUA4hog0Twu3jqTk7
X+Scb9Y1POl3tDNfZXzI8fmkMkw89Ks9ZDfDUY50zKA1XR3O3YPK90FXmBcWRGYsQ7s4UiU6tIZL
uEH1Ohfv+bZVUdvwinTNjlpMfPekh+QQrL9NMDfPBuAEc1AdeltFx1agWLqN+Cth46ypAPthSfDV
JmIJ/v6vnjqchj61Ax5nEPwkBIW113J6+lYw+AAFWh2IgjeJeeRR5k5HsorrReOYJv9pUSB03SYG
tI6vKkfsKtVY90OogF9DgbrXEddCdqkZZmtbGtPd5QbT08qCcY13ViAMUGNBYhj4veQHmUrtXWKr
MWrt30Aw1LhBBwsqwlfjBqTzvPM1r/V6t5Bk4d9E/A2ZDoOv/WrChRW4MSNzcmnrLCrwcnpC4be6
7jAPiShCxx5YYt5tWo/2nU5r4mEFiJz4gmhEUVo6dis+Ei2eHJuY/VLOVqN/kk1zfWgyI/i90Qj0
1/TUUOltCoHYBdh5wuNRaNlIMtdrMwYnJyS7pisgSvQyUuHcXQtz4hH9v31ujtddoqIGRnUltGT/
fKjp8xryswozSyGdN9jdKhUubim/CYmcNlggRUNX4ofpmvpJcLOqbn6THWJqcLsnAs96oLjMdWFg
BzXktf1u10dDQmfISq7AwKjJty0TB8DTsiOC6AmzZbxCuKufCPYRf+Pww8F0S8rgJxuGYtE/yKwL
2t2YnsYDD2wrA1sXp3PgMI/YRASpXU8rbxSri4EV8TnT5obXKjhaHXYy6EJV8w9XiUY9rAiInc4F
D82zjoXZLa4z4KYPLsM19O1rWSYskPlDyD6uVQTAiojVSyK73ebw7RZwIghheAQ38IGMC2Oo+6LC
Zbfmb1qUqMGd9LlOh+kqbsAReyzx7u+Q1jhAagGf3Xxwdo0LPSfyvtjx7WJ0b4sD4Ldu/aGKnvVq
ZEl9jruWAZlw7k8jf8ftMofra0a2E1JSrMOVqQyFjgrqPBdwHSZFq+vMHMiJZDDSEYVEYT1zw5Rx
uUyjuDgyFnoQT+dDHTmZUVtML1/j2X3tO/qxMm34gbyWjcAVCSO92uqAR68YH1mjtaSIPM0tYsfI
7+e8N9KCihoBOoIPBlu7SSoK8ejNKwAV/75XZ+a3/MuNWuhVO7vXXn4UqlwGsHpV40rwgf/zLdKN
9rK9DNfsC/215qAUyA032oqD2XLESaiCmv9i02aaLMvmBE1XNDEQ90/auBpsOpmbOikZz16MLCoN
dks3+IbREQaO1igY3Eb+V9unbozR6SYhaWXQxvhlHrfFA7Hb01PflumliuD+sVxs5Ars0bw9vfvd
hbRVxLxpw9HXbOxHrvzNUX+1M1SR3K8SyJlIPcjq4X9bRCLksQxLcfh1vzpY72+tHCkJi1Xb/kZC
LDch6BM+UmQfEgGFK+zLVxFPrhhczm79NQxeNUTqKKJxX+Wumm+H2w/U5hkgvxIlbdg59YnP77oe
9XMc75FGoH2az28sbQPjs0Pk+R8qcigqohHmD+EKV1ouzssfzPHjs6u3UgoRPqgoE6RHAdaZ9tqg
yBNXNt1+z6XUwXYzzCPY/LZLrhGvZulPcFwFM9j+Iel+xzDELfclOHVx5Ed+VtnJ7ZqXFuzbB2oz
2tzQZZf/mFTehcf1FOX6DnRzstEW9MRG/MsXIoVxlKio+LKGDVE1sQ9xR8uiLvw/Gd6qCp2SylHB
VScKC5OBvmwxLub+9YqpP4h6AKU41IfB42fDk3H+36h86XfzWL4azHcSP/hIRYzhATLHk32iWYMB
F8Ifl9/B7Zo2tyEoSR4+loKvYY/KsuE/r38oVV5Ib4jbNjYhN8nGG/RLVpoiSAF6X1YVU/i7QkrJ
jM4A3Uc8sK4OD3uNYA+r/TeFuFBLFszBsDXxva70EZ7V8VikibP3TGmjt++E3TZAR0vvbW+w7x8t
JWrgbslPyB5H29fjQBAzqZqhTs9IZRP+Kgn1vycKWMArzWluQhJwhL3/6H+X0aaMg2R3sW9G8tLo
2wMvP8HvdbrwvG5v3/KB785FohMIJzy3hE1n/EpvqEaDRxC52d1fvP1iNNafDj1YixnY9GoDW3HQ
ANsIlYyN+5nAlhDvgi1nfUXrYZAmoMhe98Voc4IsGVFS1yWVMdrEyFZFNvATURQUHbNDkhYz3s8p
ELIjmDayUsN6CqatNAe3UNQ8eO2IEvKKYos7UxiWZrnompUVBTodDzqPuAiBhSaWw7L0je7zCrWb
ozVrRDEhGy/6txBg9gwfbFt93LWpwH2m9WuzNuXFlxVG8U4OYf9sOVqwbx5esUgzIS2mGV5y0iUw
NBP09aCpzLVuznRZjzCoNTUQuG3lKgtJcKmqieS8WMc64apscSx4mkjoWskV80AH/tz2ZRWHx4Ia
L6PH1jKexCM4RSb+OO66rVzfC/V1x8bf+kib5SDkN8Qg41LXTh7qcco63gskw7JBK5hbIdFByeKE
SAHPmu+a1C/6DvwA91+F91Vr+SdWdM4lxb7jxlEuYzKqLFonQbaBqW+Fr5iX6kVavqtX+c1I+8vV
QRWtmdYJdPjznWMalfVIFvntagnv4RxvCd+6ThSqZfucAPf0OSn2elx/kfoAlh/s89AOTPLiV103
jFuDus1ChIvLi/+HQvQ+kp/SWhGWHHC2ZxwJTYbGL4W+9w0vd/kyD4QC7WqLti5Iy+sd09gLFX6E
JDe5kTBq26Lz37l5tZ/Bx39ydF5FLqdpuqc8b0E76S43TlTqHoI1AcRu+buId+xdO/i87TANiOST
wkU3T7lH2SzsJw39q8x6nS+NvGl8sYDSWBHKDW/oup8/YV0x72zzeZyoAEWyOse/7sQAsDhlC+VQ
tc3QKfBlPBAeQP6i5+nL2Fq4eLWMgQbC8fuNoUdZnAuU61yeWp7/06JljMqQvjVjoQch0yvFE/9a
MZ2YtbsMDaSZuSLM8+Q0Hx8Z1c6UKPZ4RUwQcQmrbusovlQNCBIWbL6rkgRpi/Ryo1s5/hXMZPEF
O9j/ZIkzZJ2vweT/XHXS6mH8Bkeso5kAdROsj2Q5EGhIvNyAtOmIWPMIXcolrhQhsfi2+mH0wFnp
hyYeGoV9Xj8UAcPnWyh4Cv28bsMXpisTlMqNBVPUs816sJ7uuQkjyxNgvO/5KZQg1/4jf2UQKeJb
c8yLIhd/+zCIHANmch9MzroWL6q2VL0HVW0A8UsdTBFFviaBXCGha4qXbKt78ta/LnTleCtxrNF8
XADZVtfQaffe/NJBNzFcFU4lWUWx+Fom2Ahod1LV7v0fD7WU4HIkF2osdFvOep+Bp0H8zmOnuPJ5
2bFwuiX+S29KAcuEZdVFYFXthgV1fNY34uw+P5YFD5PfPNHo5o/jy4QqYxzjHbx3/hT+8534b8g/
D+FRGTUc6XdbIDZyol9xSUn6S1t9CHk7iCXx8odvu24jEHGfeCLfS97wHMJLw1+21NjQo/wIIGT7
iNlMBhq7zrjSnnsOZHYkC9HDrPiJnKExU5mCT2cuItmK4AIN2RwIuyhEdLH611fozpj7IteLUorA
xTUzyVlKl+WQrjCmFstuSufG25CIj4hJC6O9/TUn7+JQF8go/nv2e46Ij9Ys+cj3J9rScHIMa2NS
dnIvzbSpAJEgjBZksOYzdoJj6hSNkITIQG8sx0ml7NRM+XGDtXiB/KCM3mmrJ89GyHaj1tDK4T5y
tdFRVRvDF8yw5vdQHXsmRlKtx5I0fTCH88kBCWqp7xgAHKu8xAgCNKUSzuZ2hfGcQrzfPCsHSsX6
SSAWm/wJchU1t1JZ/HwbG21ueREMx7oKRIdIu7OvoIAho9+6wfKVzTxJqi/svjfJAPc450QK5/Jq
tqFQmPgqOky1tF/0hdKL3DeRGgwIxUuVD2WtjRbfrYr/pPdXwSI7AGyfYuLf941iGFmOCiIvrYBj
HSJK6TDKXJxVW8UX4KpE7CRFP9YQpToLTeIvZ+/lktWZNvCA89khS/WETe93qiRk+BQmMXk8o8Yn
Hp0lG9dXl3zLPOeaNP/5lRM7tTZftnmK4tKY+kE8nmVlfuWRW1mHJlXOGZxP1MbQA7Sfe1efcD+8
X2vs1LhVLjWwXThsk9PCtifeo0fK7GKn8EI9cvaBns9T5SXgN3/5XYzAT4/9oDJN6ed/aM0ngYyY
DVIWrPeGAFxZ2TP1q+z7zDyZzPC1VcvugdgJx/retP34rvApzCGTJNVWFQ261ujWUTCo3hTljixc
xOX99g63MSYH9QXQz6VbE9CWIOUHNRUHlkqX4Q7ssFusCN49cxGfJzR6d13LrRGjN9TXlkoiBcUA
WWA69E2IDfP9c94etAvw7wKmKhby4pq534YCUt7HwQmNWRwN3fWlos6pX8PS+mNgM4wYaNfSxOU0
8MBbJYDRs2PQLFszreYmCU0TGhcYhs1jERXB8XB5CvySDE/aiIXaU6HuDsjgdw18AW4mthNzoWrd
A/RnYwA4PY1PpiUPpjJ9Jg5UqZz0TCtGLlvy5CYjWP/Tgsff4TeNes1k76ra2zdxDbd1AYSe+iui
ERGN5AjYzMi54niBpZkz+IQ52v4E+eIYaUy+/Yyfc9EVO3q4VJSZIOp6Wbb9JXIv+jRS9SuvCuxQ
xQcnq/8DpMyXKfAai6qiB9lbuNSOMDoeU7IvfUDpFxR1XKJlZ77MxHD64UwzSmNeNWkAn2R/ddzJ
OSWi9fgDG0Kx3icqRQwAQEx98AtDGWzgvRUYj71T6pmm2Q3z6VEBqPRM8DSPAzDwhvCHbh78BIJy
m14l81xzOM/u7RBKKjIfI9ZuxEyx/8XpmvSth5fmNhHnZ4wnQF5gfObz1E7L2rkxuQtxC6d3+MOs
ZqQU5yZneLj9W8/L1uobn6dOiF1nYmoHLDxjWVtv8RbqnY1mbARYWdUIybE5o8QgQnkqHlYx/CgL
LqNhjfVQelt0eWhYdIovXC+AnfAe94sFzicQRPVdxj/sJQM32TLk2kq504CnSzh1YR+QPqtjWgq5
un6ztnY9qeIbr1r1fz/ZPNueMptdwhe4KRFmNtwLUImrcQC7cPRdQTizkhVK757i8ehTeuHMAtZc
at71Iytmnxf+JO9IJVdCr0JPSc2si1bLT+EPNZE/mBXbCJsHN5QhN9FAjldZZO2ocDVi/yuovClc
4Cr008UpDH3rEr46UgUiywgo8V7QEOZXY+F6eHAPWgECl5YGSqDUeaqa2SSntforB9nH+o2LB2YI
eUaGqkyQJu/iuCgFL/u1NBSb9a6EVpav7eaKeegRP5zIuGq4LC5Pocp8gjEHym+a4NJ0GL1cpu5H
wJqMqI7Opdat+HIFuaw8xokYoSf+rGIIEgo6+tKNGDqE9QqCNHehC0RVFRYOIjt9DtLNWgYz3tZN
Fr3P9MCJpKpcHTbu+AJmWhto2+AdPggNZVUwUZRBPo/1cXU1hCPdqcpdpsEmh6SceNwTLBXypFlJ
pbNf2PuRbN+jcyNMnGfoFFhU3Lw03AIQUSSs2k8G6nSFN4qmiqMd4ylsxWvO2p2FuW3QYAKHYFyQ
6AYhUr7aPIS4cGRSCdY97cBKgd2YY+Ej4L1wlFfQVgk62oJNK6c7c2HbKMxqe9UR1sVgDKFRt3M0
f5USyf2WYZ37SLPEX+Xo9fuE3pmek/htY/A+5Ey372MDT3aXrZ2f36zmY+l2GDbcgPV/0gzTOYK6
sWpMkZYDhQBK8ALldRU7kM9yoHVHQ6ksrE88tebje4+hiewL78WVY/NnAsVYyroO7hIW+R2LWijc
BYjaSXtOzEy8l5OMdlXcUttsUTD2frSIuDqYKhVeu6+GHeg8NhtgvGUiXTGomBalmLeRQFMVcFZS
PKOgYgJDN37lXYK0aYIUDIDEEqNPzrFIaYdFKfZfMH5KCXAjgboDMQRjVQQxbJMvhk5+Ae9ASIgo
LXyDZgSalhuDb6D+01uOLSyHyZDi26pk6Gh4M5ry493KNrXDdX4nEeTtH01ciUNj53W2lUnA2gz1
/ho5Hcl+1pvuWGn5kWEQEKL7Mdxt6FGaNvb67z59hNQy7wTPkmIRy6VwWtmfZDOOo2No1tOL0hKE
NFpRGD62GY498yHR4qZG8qup7GDwkP+BZl/Sq5opi5IR11VZw9tn55Y6oPMLXgr2JhQFQCoauApA
2JCaNF5eavTBhKPMdHeKhtV5SNv8/iIW96zJDcETOjW35WtcrBDYRsiA//ChOhYiYrnQJ6StFrhf
anrDgYxyIuMENODWMO7JWSYjC2UNyv0r13RohaG9Zfyd8XxgXlYK27jjKSCH9soBvVuin8fgCuyV
Gr9NLvR13ZUUl3JPNaJEYjP/XnLYl6eI5dVkcNt7iiYxOk5GNPzlugvvCZC/LLDVgas8E8vxetPf
xlTadZW1R0OD6HPvxTmqUcW2391APYJeMDmyOWtAoxrfctNe+M0X5E/QI6Eh2d36yHwXP5m+l+uj
968Vmo32NA/g/54G3rTDT30ABSXzvAnr0l84xk5n/EBUH+ZehniPBrhB0wTN+5rNy0LoPkaknQSL
NfZACPrw1dp2zMm7MuXlt5tLsIXBmsuBItX7iC9lChy88jC15M9CL0UEZi/wsh218a8YQjnVx6Co
rPAUv2DFHTOtWyWBe4wERj2jih9uRO6sQ4S5lINoPxcM/sj3xbiZl+cVulJR7l7/NuWVvbMegXQp
9rGasLhs6muyYRBEpVZ6Kd1KGATcx749oZxKt+1IWTM7KNOup5WbSAJ9ksUH6UI7/6LBIoxaqa66
8vTd+oY4tMDGkaX8U21DhFcRL/3PdWPNtjmQwPgDL5cpL5X2C3Eb65Mj8VoWbD+gTX0m/0LeKZFj
vfUiXKN28M9MuPOqxKRdyzYvkKqrtUwoFYxJxcRL7/TZ651b1vQFEbTkPUkauI+pDNQS7cwbKqh3
9NGC6+eiXUbLTa/qjKcaZjsfoYWGy3nc8ihQE6HdIzQQaSsjZc8tPcu1sqK9PFMz1utNPaObB3n1
D0qy6D+FJWcRsut6qrkzwkwcicprWfyvoXpRReqhG1GseqE9XSz9fEbgSTabl/u3Ij2pM75cxBVB
FlygXu+/RKZR6UjJQmyVpYHzm4oAf63kY/MvIGXVoTtQbWgtMCSk6WciRWTFlE83WoDftNMor933
ymhSo4YNVr2CBUml74xWH0LFLP53ZAG2dejWjGJvgkxpy1N+i/d/+fofaZmk0ST1J+z7yhM++vQO
QiwBPGtyv0iJPkLpVGcUmdtN4k/GUNVf0PEJDP4J0vjF1okyFOYSeBVn3bXQKfxwjMgXAp1uUa+d
bEkvKaMejiRRgOtL0PXkVL2NFht7Mz++HUnmXni2b7A+eIdSOQ/7xqrser/Rve38O770OdPbqIK/
DHy+kNx7ShGShtH42HdBjLflz4N/DpkRmUBuAmJSe+PlTTHgx/AQjw+ouZUBnG7dhwWMQza/8ncx
2ojGs6UkybAVEH6R28AAMBy1rYhroHb7Z4ycE1Eq32SHEX9n1D7qyuji0Vwt9maihZTV2XGv7CCk
3wKyRwdPr+pnobA3BwWg2pMHtobYbkbMtU7in5n4TFOOBaGJ/G2r+zQoAhj65naUYpzcFCUpvB0C
LI3MuLeDCBSTMoipnNfnOc51riWl3C1B3mDdQxbydio1sdI0vhUzhnyRQuuBu+EyKXzpcXEkdEHs
cUGXAbOibpkYL28m+dWladrLWPZ2ezOyiKk+k7E2MZWDA2ngVdzExxoNdxBJCJj1kyfVH0SXWF7j
IsTCf+d3qb3f6EBKd8+cj1jgY1UIXc0oTOY9XtGANRWbqdqUsHCp2k6cOmQWthxdJy0QZg8Lf5JM
uj4YQbxxQOeUwpnSSRqV08W3DSP/meOKlbVLgntTjRd3WM1xnSySe/3Es7G4KlEIb/asA9wMhBbV
tkEY6bXzutlSt0MqJpbhbq5lKZWKyKySDqAL5JEPPkrrDVghTXithZDmEtaFALSkqB/YX0R+ypN0
FjSOJdMVtjCWtqwS77secBpn9x0Bm7kHhK/iyyIp25RKuXfRO4vDclY492imJ3RQXShnWa/M/jgD
mUR28M4G2UCBbKFpwPuf4pN21jT9M/pioiIwDVJKLDHjYD7hJaTD+HboP86N3nI7eNtr+CuLdplu
56iadufeFYR0AfBtbZAcLTMycXkigF1RZxF/WFd56x7L+uvlUwymWDGOvEOeRLyP7fCvaP6tF235
N24+RsoEa6vuCy/KWHXWEmanSBgO/Y02XjSqnGg1Ti79gSzcQXWmraK6c4xFYPxY7lXOFe6dZVPB
uNlETN4iWQlgkXVGkDKlrWuqEV6CZ8WEbFdGag8bimVb/xP3RT7k3EOj3uzpjLh3SyQbyO3YLNZP
9KYC1gaz1y88SgTitzk6kGL4gVQkXrmEcAhkbdU54/QaTU926E0+hIw4ThC9YHLbWtfQTvQV66AV
ADExV3ayxwhNyBjUEdeqkmWB8MH+8HKmAXH1D8/qAmeDcBug1ueB/x02vw6S/eXjWrV49ApjdnYa
OmwzEauEHq0qfpafBNXIawWVW7RK68NjmH8tDJ/7eZ8/Q81QrQL+YG+6rYvAL+1I4wjwdevUgVhN
pHlQ+BKA7JfboMCAv/Oiisu7lFh05xByKn00c60yyi5k+bQSiTw9i4K9zqB86H+yDpCIi5pr96xI
rFs/i3cr1WLtgo0Hz0Q6yrWpz/OFujncpZcv5Q5XkVjkaMK0gsTO3rCVGLBH0yaeqMURr5aGudEm
Wf/4EA8VsMsJ2+0862El6hbWG2b4LQu2OY0Wvhb+FaudhcxD0BnglBQhRJd4bDVzX/wbkQ0KxmOK
vgxpD9s7e7M0kxJPrgLO7vNh0uTSYHhLvegY/dmB4sNKqu2FnFVX6rL/5OQ7xZTLY2kePe8ZMjbP
rz/kC+WFkA/dUZYGvZc1Kwc/dPWDETS6+XzsGACkWsOZaTAtVEytjDuNwrRDVBtikOpZTci1/kmA
kB+Ru6JhhyaK3Vw8tCBSsHJZPe6j+4WdKMVswLs7yBonqj4OiBQLVk1RkI0F70okxyIDWbYfKkaK
cVg1RFBZ+LeXGjzgrzV1pC0ppGKHQPaWRqH4p1gffZD3YrnyJJ2FH9nuKGwP1xbacw8/cS5VYFNP
WxypxEYmdlmVhACWXTM8DWC4FvQG56NcByuAxKBBvuy4KUJAbEkVYOqbABPh5Em8BavZx0AmIxQr
3fYKhmd3JN9Yb4rOsrBoB6Zd5blW11wf7VxMdv2D8kCZc4Z5F386lNExU6YpJnUVlW9C5gO26KGi
At1oaUlIMWz6pKDd6UwzQgZ2C3lOcBOCXImTtqwKzRM1Sg9jzUO1cYWN4DQLS2/WFBfUvWSUqH2y
LCLv/o9VuPA9NbGpqE7kC/4zXT046kkwmgGNEhIgSwocFEkarNw8kDcLXGcS5lXwehouWoSrSOay
rFmfweW3qXIQso+M87xtA4mPsabfVtm1lRVK3VhLHJKuVq7RAbV2f0SwtGynN2fF1h513Y60FXAe
3GrtTTa3wmHcI6H2CyFBvum7+cnDPDGRcg4Az1yqMAUjbWJZmU4qJP/uyNyBjK9hlus4YGQ0BSAl
aEQOtCd1RWZzGMGnWe5y72t0S4Yw16CZJD6jTuQb+XDiE3Ph/7Ch0e4/4aulrN2N92o3+ldGtSIz
Rs5GgxDEUnLX+9Imvdu67skrc2ioqeUuChd2meB2HZMowrnF5eUkt5L/eRJcrDStKZSgEK791ueq
fQTNPZuL7/Bu+HygA4h4gZK0VIHXuz3yWgIChe4vuyBMwucaE9mE3CONmp7ngUR4Dps8Iix+llpJ
mufnlsF5v0fiS000gnkGVB6gcH+e112uh/vvHUKw4Hn+R2gY37dqcF8dakcKRzfuxBpHAeVpNB4D
k0eion75e6A9dNppO8pAD6LXNP7OKTwce6fXWUKT8Csp/Xw0pVYZfNxlF//ZOG8GFl6htwzknprU
UD6e2Oc10JRK7gec7zjBVwikFcimVCJleD2QoF1epVoo7F5ncRshddhbvDRJyZ6HVopOemOFXFGT
QCEw5wQohPkjEDbrVD/9dRbjD0k0+PoVbUMRK1tEkISh9FkmTQ6AZ5ZrkawcG7DOB/QPFBHN5vIi
+oYgnR6G+ww7kucyjoTjvh1lLWZR3Zq+Qzj1PBe9NQ//WpcBLfcSq+X24yoCwKsChxjVRivCFtEf
f3fotcfaJug+KxboIaevAvXMgjQu2MeK3u0jbVrPGQtwz7pfQNe1oGMM7YfEIfnW1eY4g1XYF1LW
pZy6LmaerCn1YjfB01jWU5lOl8sECKlBGeferdOWpdzKJg3NEreaRok2kzmb84K8p9D4xBsIrhSK
AdqzfMiz4zjJeIb+8ZUKxWZrKfO5wXknhguamJNCnljJXBM3THwjUcez0ksHtStcpa4F3aYdqPNQ
AxGVU+WAs/Vr7echBFEY4rfCShffFvfKNBuWP/Lf7Rule5dR6Xmpr9CZx3mXlcZ/VsALCZ+xdg8P
mpyRJfWSOZkoaiFCoF5NxodS7vjJPzwqm6dAjYhrjr49/o/mwXHuA3plNKzWnhhbyDAql00TRvR4
8ouDNoe+1xbg1z3GWvHMZBS+V//fDdL0jFP8bcG8MFc6JX2ariFQNiDHKFLiKsbDJFIAudz1BhnQ
6H8Q+uP/vbi57RiZA0819FRTuVTq3YHtkQ/IyXpUItfajolGjD/Nhv60SWsrWpYKCKqCuIatRq4g
hrfGKytXeEzJ1scF0X7FEpduwgaVSFlf+U1BB0WxsqWIsFZZRZbmeSPtGEDtfqiCiDa+0etypX/Q
dybXTZzo6UlkWJg+70c8gvaPs2ziXln4alSeWGsCHmk+Q++NPwxjhbzXqSXmjC8vOByK9/aMaJ8z
CGvBrqVUxjvyPF7HxGR46cB43ViXJRlTnuiFLFaHefqpaXeZyB+kGkf+GZsf1zf+W7mXVbLOPm3b
+fYTNRIgHCHRDX8y3Ax/eZyXNdTnn/3gAMlAor8gD+kS1WXFn3zG1Ov+iov8SzUKZUbRSq6Z6bOj
sShqA32ZfwUZU17FqKgpumZpmymsq1jXP7rfQXlxEDxeG+vNnKLVqkFUgVzAHT1GPOYbm5TUX2Xb
VEKVtwXoyvfLH3vJZBWGHEvITYq5gPz/YS/CoGLKODcJX7MO0DmdQzClgltMdnDqgiFVcIaPqWUY
RvV0pQlXNXfMEcHgWEk/0RFyoRsz9r4VF3u0FPEXIj3qztdu9ZtaHiWYB2iGVA+JOzBzuYDfZVKt
jaVuyc9f2MdR24MnEWjvDlSHKevgcC4YcW33cV8Di0G7dhi1tsxB7tQRB0kESeKKoKtw86ZU6nP7
vqV+4jLb+X4qkKt29SqLJOfQEYv0yaVVeMBLn3qVSY3+s2D3TZRWbKNHHxUcHDDNr3XiRvavtgrb
xKgWIXBJcARdbwBt11t5ThogV+ekiTuBkgoQlik7yx/MW3zCPUfGhpDSUg+y1duLAupDrIK0eYyl
0zd8LhONEl3DiHpxCm1gd6y5kkiQKPqixaLeeaZJtGxrMHwymrlOE0YrbT71PD05ur1+7g2CTBIo
hFATx9VbrNsAyOxkr+gdJWakhS/ZBhuCHBRnShBp1eoKVfdheCRQDoIch7tlw+MQJ+KEUvwdU07z
InaAETDyqDzRJayJ9rhuXWAab1pOrGY4a6btUAOSnmJ6iAI6HFDnOxLFE19Y0n7u+9xMpRk5syaX
9w3bW6iYDU3F4AAwvBsqaE9H9YzaJW7fPFZh8orfc1Y/thoTGpMkiVF0xZAfrfR9S1krpyDnkDkD
6jLqgUBy9l/qWCqI7p2IDrAq3XjcVg5ePd29uBjOEOwVl4lSAK9GMKXp+L+lp/xWy4+SAmK8+ayq
PtcDlsTSLRhRjKlwEgY5y09YyTN+0zGNHUmFrWvkvcxSOflVuACZ7rOC9ysAml79wpMLVJuzL6NR
D3rsChs6JOLNioPCmOnTFY3UA0C95v+ayXzNiTzHSdQZTuNnc4nD4f89OCmdg/rJSkxa0uEkDQWw
QZzH6YTXyMGoOsLBBSZqJ44vy0GH1TDmNQWFQSMQ8kVTySbzl3hwhRvXkaOto5vqAk5yY4Zjk9yq
VPK2RYaxae1Ft5iCC6mfysWpnSZA+ADUMo+2GI5M9J99mcrjddegxVrG9SP79TDflD62wknCB1cQ
QM0Gqswpl8wz+WY+EttTE/t/l2DrG8FFh5m55LII1dBTgPwR1oGE5oqbFxuXXZqWNXwUFqUwUwfp
XUMor2AEyPaj8kE30t+YqlvMkVWPaxq/eSg5/Yy6a/C9VekGfLN4+4WkEHmkExJLkOOuRfQpfVC9
73BrnZFYolvZOmPBaW9iZ9Hq70xothESlbfwLU8P4ALFxH2TuLLP2RasORhjoeGIkxWoRHII4bpM
1SbyXpPZexoVX2DsFSnCMI1BUMzQERxgU40MCeaLjbA6qeZgqJ7Ikxx7Ng7BXX/K4ajaErnDdVWH
lyNGkguwYpzvMuS0BJ5Em9fIEiJJa9CSu2ctE3rchgAbAwdMMFU5On+SyPjJsSyEdOAhuW7/LSRi
1I15ty/3rVfEaF9Im1eEm0TjNbMFwWgw4Cm17y2wmterAMPgzuQQ7hyN/H2gzuEL5SiFyIqe8Ofw
VSiFzL7YmMB5IdFZry9l/HFBSwpwIY2xIGpUt1p0pdRbmrn88YmBUzk2P83fcCrmoS37OoXexK15
IBRRkudOpJX9LT8Bxvpu5wEWndII9YvsKtrkNZ9WUtkPAfq0VGz6yVinPI68AB5ZnlzOPEmNYTK8
c7tNvGfKVSt9swc5O22Q4GMQ1PtlD5a8X2kpOyxdRir+Ot4zGyVD9wBV4qFZma68DKs5S+FqQZdN
Szddn2Hiww45QYC7NccL+n4jfHmMohDJsOw7lKtchs4Ira2MRlJcn437JNqqG1dX2+0zFrisqAbO
y0t2SNv+JswvstfebJ4SIa1d6sq7rpxgzGMueYwLY9EOdcBnJ4ouTPjdFj+uKiGX2CdzUqaOoR6I
fykSWdeBy4NJaT9U/oB9xhRjqK9ePxPDTYmxHQl7XdY0vZ9Q7ZA20YZvDg5BdMfufhe21ueHLL5X
XLdXqWdRzhYqImBMTz06YC9ltEYoNX3kIf9i+1o4u6j3u86lvEbIiUJ3Kyy1C7R/pTM/mrYEowdB
o4u8bhe6LQZdIPMJ0vGxxbM1fl34IzhbB0LsORn36+D8+eVqLcBwC3xKzeMooq8Hn1HUg7zkEHZh
Dak71607l1pWnr1YQ8RSxrH8P6bx1kjgOp4Hi0XzNxVboPK7Cim5oJM3tmJyc1o4wAyXm//v56dy
/Wv2M9FOclZTrcSaK33/cRhZnzUB8als0UfdKpJXQBVrvI1o4Id/vN7iG7khvC0t1CRQZD4LMGML
3b2GawMMi4BmgsW8k7WuqC5eXiSGtQbhwgxlQSGb7a8QZqk1zuHy4YXXA5eYAi6Nk9zT0SVjCevT
kczEG9RPnqaI42CBWBSGD8U4B9ega1/aSMhb9hGKotJzUR2gWcn3P24gV8q5g0AvXlTii9QYFsPO
6CEU7FeK3XrjCbpy2wHTz2gXY/bSqyZ9MQUtIVWxbzojzSCViMhaR0ETVfKhHxsXDC4mproL6qIK
jbJob7p1UPrHGJTlDXtthtBENhPUh16SYZqYqQK4+qoZhRQXOTd0J82Q1eX861XifCYY2z9m1ttV
kB+xqYEublLz2M2uTL87Wu5FX6dxZxvNEpL7Mtk81FuhziJYKsCyOc7dDq1faykZ2x2C8P/ldNVU
x02Qs+PQt6tjoS8UgQ9hDIm0jOaL4mDinm6DTu4PS3m6HrVcBLHFssDNsJrOMF3l1g8XScgOmnmg
pzocPS1/Q3BJhyOnR6OslAVzhhgRVsMAhtsmpkYhWzO8ywpw2Pw4LNVVFQcY6UoGFvmQFPVrSBs9
2GJGpGGPBbWZGNmCZ4hmfMGJVrUwK9z28OXIfP9vOGu1Yrs4/M+lAsWiZenU0ZfqVXu8jGZAsX++
VyuRLwcjZ2DCUCzFHXxpZqASOkYLyCiAeIDFk1jvQniWMD8+RV3/esZbFX19CAxCYihkv6AQC7Fy
F8/5LKmm0YOE4I222gRMb3r1YXAig3bw8C439CYarUKdqqSK4FOnnNIeXQiuqqHjikaSAcU67dK+
Zz2zMziLtKM/hcb5XCyqsPKAuJJUpaW9wirgWi9wPZBxJ2TbcwQi3lZ5nVGA6nX/tQo0E0Enc4Kk
PBEkRtoTX6lobKpj6k8GUvvhEujcemmCvx5oaBoxaO7zIRWQ6VBZpVSLWL04XEq4h/ZHsVSGQqqo
jM0v6+hjI1fxdktlcKLC1QvP5A/SvC9q2MfBnKdFVflWPRBVcmK1YJ6EqQFqyp7BTonhNL0+RHtV
7WLB6OXSH7EJjqSRc2xMuJQrETRzwt190BwvXQVbZTXoWFG4xvzPZfFIYikeIj3+Fgs3DYLzJyaz
ADR6A5bui51cy/l3TsJ+HgnO+Meq7PQ2QcwXqCu+K9wCuIheV7yAwJzd6OVMDWIHk1vHRsYc4+HH
kKxDK47i3m21eMt+cIOWv5hkWJ7b8kjzJs5XCaVqPCdlLlGW+G3/pr1TYcKeoruhsBpEWx9cRiJL
A8yF3jN+SA6AjWGcIlk+4gdPlPxuIPVXTjxpeBx7IgaNLXGCVaeY10zUIF+223QXv5IGmXA8q6G5
lFbpztRo8lfRsdi5oA7ySOesyNN60Yuvq7OIFW7LcWph1YO1d1kl207Ng0eovjryUBsalohjTLKZ
pzDPm8uiONPIAi45DklldbwSj6bsu7h4SIDGdPvKIkE64k8k+G2r5gVoQYrPXERM8zrniV4pNC33
YPzHPzXgCPK2sxULIDH3N1fIjMCURNk0jrIg69c9mNkK+D4eOTFLTZiQy8ei3tqCNOB39gjhNR7i
WTu3ERfCaASWg4NzgUkoHRN4ACX6xC/cuZ6lgL6F0JA1azvYmzchnOsBdbzNKeAKM/Jaxz9dQahS
2MPAtBP3C24NMMyMGu5p11GWmXJ371ymgqIO4hLXPHwR0s2VeNb4F65PiM5LzKr2Whbca6SEhPyK
LqGF+h6LnIE8naBLS/VUEjFcAW6cwk/Azaqj2ZZEi6S7IxJYapZ4Z3m99jQPx3aD1Z16OIb1Jzb6
BE42fc44uqr6nlRddj48QW7GoZA4AhelFQ/IgsSyt/ebEW3aJRg8tYeWLC4LmBFERmlSeQbpYm3H
EWPvAN/E1J2Sd7ZqevCBjTfOmpDVmQBD76eigg5NxNsAf/XmdzIeaYwgpArI09dLvNJcqFWsX58j
/H4unQ8L/TGk+IbDTuWMoOo1ASlpKyTQQHor+P9JIS/zHDChZZlD9cfB+cZiYhCnc41ESFi2kAOi
nRzbNF9q4qg6SR3A/K4yibelAUPOZ/bM6Yw4Db/NLLc4q3stc541iTpjo1I9/hBd3El/mvj9gyjd
5TttxeT2DaTtuXGIjBK8hZME3Nphfvuq/5yMh7PQZhZ0NvWT+VYUj+zhFtd1we+1MH9BSDJu8A+I
4Y+a0phC3Kf+JUB1ZrpX6342Ivbk1sF9PW5Cq40mN5N/9S/U6rUXQIswTQZ14PErErofkae7w+Fi
ZufMn87DXLhgW8A6vgKdvDe9u4qhWfz/3SF5dM65uekKPBh+fDYHC7ZFIWKTLBLxbd/XULUSoQob
dTbJhPt/67vOoa0pbPMtz1cnM0ynsn8UDH+i4lrer1nmF5e6DjJyIpnufxMiQrC6WMtHOR6eioSI
sm9xZBocdoEA7Qk6NJMt8irfs3OVBJq7Ss1FT0IHEkBYnFmcWq4kE9XCCuUdIm+66cGaaFd0S8SC
5jsuJPVFegwxDudTyGaTM9AkTIF7DKpnCdSH2ls9vSDNzwk9kWxHGU1OZ7aW5tMNQPOhp15obs/3
2ZM2nsu04DAdjpmzf0SnNkTsgAg0yyP/P3oCv078YCQWsSGwtZTRUW+/ku/m1Wp8zz1OW7hK3Yd6
mZRbgshM/gQuZjDweqDDSoPCFjb42oTriYjN5L7lkLlL2YGylFGVR6lQktVKGPz4b9J5Q+G9ck1A
TiKCXYxHWd8IGud9CoVjer+kYkrw3/dhKdsXeM/Br0/If/i1y9nC3k57q58yGs1Y9f9/+fjqXmNM
vnL6hSzhcx2qBNnh1mJ7C6+95Nt9LiSN5PA8p4BsbpgSPYp2oG6PM6o4f2QHgH/87AwnsfPUr1GP
qjCxV+vcQexGquQKj6I2ld3HK0Cna+talQJnKpFUrDe0mc6ojfPSDBk+EncYfkCheYFNpexEq/th
GqvrgOUTDuoj7YE4FxIuqxHTgZsbh87Sml+Adr+gSkq0RtbNBEg4BbuUOl17/w83DSACEZbapcsQ
DQyHvPhRnqi5HQa4nJGFZlkGy5b0I0F+pye/kLhj8mQKqoLSD17KahdY5p+zIi0867qkHJQs/w8B
+GxWnzRZ0lmMBXmPIhYE6bpYenVk8Y7ytRXVbLUp6w0xBikXZNVuWCrdXV4g8L1bUTVYgLY6gfzG
P+GsrQn2QHk1Ux2qwGt8C2iM2Nxyjp5EvRLwoORZSrfavzVy/6Cep0/z8APzNIWbUdFJYZdrbRGv
ZEAWJX+1R5ceJd2NSd1FHx266PNt7psfsXtK9tWctGqsujzwYjIp4XFyPAd7+uP6n0ErbBoIXbX5
tprARWsl/l9GLHflR0hvRzNw+It67+BtARHyIZve7liMX1kzqq7u7RJ3z+Bdj/URNqRcbR/cseXN
4RL7iTmxfbn+kaGAkikc/TQG+WYYDqeJhSlEWtCmw6/sasFuYGsbhGV2TA3QIVAt64I83IiszCXE
eWuptgNoa/R7QievtMJo84x4S0tnZ0c1QHTIzIAJvmsT6Nklh7e2lTtaGImhaulN7xlMdF7jow9u
+6y1dgtBN4v1ddcBcdWS+moDR85951TqXbOh5qxW+6ezlWCiiOMD8AyT2SQPF4us6yyPhKuHIRle
TuR6c6ciMX0KLKH7aIks4jgQAKM8WJIW/mzOEni47U1jOQ+377+vAfRFtJagU4xWplaev4VcAUgJ
tu3HeyshfVKe2xRBdR7fJJhuURJixu/9AxyECb59/xDuahnxqOYU6iawVD0sSybRWQRxp8Ubwcbr
SKscKmqZ/ciS3gMO89HWBuNb3DYuuJsg+/1wgzFKLlYnHpxM1NF4c6E9Xo+IVIiz+7LQeW2mKgaT
eDcHTRcgihZClUcjE0Bl8YWOeMR3Yg94pTL1SwJehimmt1gF/iemWV0fz+CLKdz8hXUGKKWVzatR
4B/uDEH5Hncy+WNfK/fE7qP5nlMgJnPtxMgQ/4Mq7cUTmzgi3SnIwRvO/1fmtKxofcSe9TfwQjV9
hq2Ipx7CvAeXaPbx/ZnCOPQPsNiy3+jyBBjSHExplKOx9gEDvcXNV14nlmY4I9JibJmTMuu/gvk1
kFg9PUO4k1Jeg2Hn5l5i16oyA7ZqGdDy9fYcmAQeWjbXZGtX/MBKkkS6FW4xb27iV9OH3g89PMUt
NUUrxDNJo7gZpfCNeAY1RFHjN8SQCUXrVv2mbhxh+WqmBHnJ6mrKGG8CpX1l4k4XmkCR70s2a9Sp
rFIPm/AbnQViyhp4467vv0ViJKgYhEE+1hBHk60fDgwju43kHiBD4CWeevrWr8s9H3hlHpv+Dxz4
NLHdGED905AFCpgwC7oC47vpg6xiPuQ3WP+bx8ju3M5yPUMEoIyYagR4P/+bdCDtXmkaMRRsdNyv
3ZAGq4JcTuH3Gk/+fyWszX2zgy3c3l4xxAyXUQNw3MwX1Gawm7BRL7jQ7dkqXe/syZnI2tTfOcrV
JnqFXCprAQuERTcZMdaRTNFgI/lEBF+iC1IEPIxpBwO6HO9BOkfu0qb6m79nyeeA+4mgHbbCwsRP
HBitRB09/ruiEqMVgjkOJ7zzYTawVBK/v55VcJ0oqWF1ziorHLuA/G5XWJUGgTwsjGkbS+CNr0RH
gZFl2qImpR6K0y1CnrZpMfzv8/G5CT8GCa7xOhAgR04cRohN7L5Y3nco0NPeGBa7QBoXyPNPQhPH
kciPwUqpgND2qaWgjOpB13AdLdreye4eJ82PW/+6LEs4XsyUa5Qrj2Iv5kCLsOVSikQsf4YK89Gd
txnqRq8fqRSa/viT/Hf7napRqoN0+HXuNT2LX3qylE9+J56JDbnZdDfSeZRy0qkQUzfrWjCmVfFJ
9Hla00WhTTg/C2EA8lizFLmIO2WySC8+dfV7iQ1X3YGLxL++d/yhglLZErIsFOiNWqXPaeipjaGn
8y1sIWBxjCiJbO4hAEkfSuy4Wfg3rUvJrG2yy+kWjGc9/SvZnhKZSJ3FaXytkvoX+f+IoN1/A49U
fNRowWI9KoI9cgvoaNAOJphCbgTXcp3HwFr/3Z+JG3cCyGuNyIeaIKZSfaZ4CGh9knnQnfS0rELf
ACUvc2iHYEWeA6yiLHYaVIA2OK5tCHU4Yp5O9w9Hr8rzinbs8aaAxDgq7x5h2Y2iTj7I7P5OyDpb
S/SQH+t8VLCnEMTRK9FcPbdVHiUsaIGvMeZJOy9OAc/k/bXkKDqRJp13CHO13lLsoU+jcZCwfSS/
2txA1ijz9RrnLya/BIzb77KJlDy7qkdsr23gnlaHFqeiL2IJVIDiFSxdR9qTmHb3DOgoSV/ewAHy
Nf6INcYJQzKSu1mYlbxFYCxpOdnQaZCfnuh1Fyr/5njvg1WSFNoqRAFcn+8RU3dg6k7VRwyb/nOs
6eumJFPoUcQD5GyCYBvkk66Tq1yZcl0PKwg0oDhS5lixhfrPXP3qaizVmK6gt9ZpWunDr5pWgSIY
/ak2ZU+acpntHavaO8jfSJnHv44BWM9cMFek2XWBmPHZAK1iba8WgwKaFIGI2h3J423BIrvxAnx7
fR/3AqJWTEHtFKXsh8fIcu38KGH65kUq58smjE/OY5CE6KizQ+7mGlVBzdjg6MW+tlGLoxs+2U1V
X1qxe/why/121OzRrQmu91ZofXbvXLznS+gOYMzw64M5nI6nKUp4m27Ia7aK3wyXi4Gwet9ckIMm
q13qLofFMgRTH5Q59sZ4MsLQy1sxcNW1cvEj0wW3snd/+g/yOXXsR3f8ek6hhOYSC2M/dOXbrkML
DOWzaEZSwJXZOFqFHRdX9iGCxuWo070fK5k2vbDOQReh9JR8xqZC+Jo38reXWF6vvaBHaqsiVGfo
osXdUMfGxoZqA5pM18NmSnNNSLwgZqSYP768qagz97CQwyYVIt4jqga0EF+soPAEpiECcssdhzVK
Of96GF165OqjMGIVWCwLffxWYVDGFf2GXqirZLd9qdGFtF+h4RGkFsMxWZgLgrDy9kE4kK8Lya0T
lPgGUGk2mBaiX8CRWsL/XM8un/iTyjf0X9QYK5gSuTKbpdcjTPgw2AGoKi7bgaKuLJCnxTde/9vB
SKRmPz1YPXqfzG6usm4RfCvCRqQKIaLICCJyytfcPlndrScjF2hOpXWOvFhufqY5GmS5SYbz9i7n
no8CivkVzKCTp/rdBwOBlUX7RKiXdSh/k6DL7n3RwiXOxRVUtPGpDDyrP8Wt0cWsbPGTfVlwx/Ab
jVFR03pRAs3WROa400qs/Le4ywkvZw5pu0csHQGXMbQlg6yc2u6Qix19ruSr1xPYxil1PBzsX+2P
tqA47hTfKHScmA+mhThz0XSlv0pUY/Mmvg2kwTErnnUAGKlNIQngcNKW0Y5ZnGA0TuurGH9DeDYB
amqWEab7BBV23OmkdVnPDVG45JRY3/LF2b4Y8f9GE1izrO71WCrtRdfxsFTARzmkS52YdHp0OqlT
IAc45kaSb4nNFBsMe2z9VJQDmB4yAun2T0QQzfXOfXpBMbQLMp2KBjXYtwoOJjSUteGNIbPnvZlU
XSZbZWOkbJj0sao6ethALPbgOe1/cpuxTakeroHhUUQFrsCK5Fm2i73AIjBSgsrbg/DmbvT6Yg7J
fmLqf4fyAN1q7CnLrKZc7mVQ+sJQ3SOPHWfQhEhrMvWp01HfD+MHrQ0GwktOiOwsJwxiI70vMRAJ
8mNgHa49eq4j1VFyVlSoQwK43HXXtn61v1nHR3Ebr92tOWy7gC5h2lKJGZgzdat8ycmcFTb9POBN
JEJKSWX++6VoYxAv0qv3ttpHrIV8UsZRxkSMUTQX6tU4X+F1/sYWNwNnzgvxlVwnl8lpVB1Fs0UB
yngZRAxsp8CPZvoXKdyfKRAssrxAebDUe946pj3u5xcT1/nV3JtAK2HtNzkAqJr00KW0EnlAEMUB
stj5fB5kQFDCaceJOTDZF2XTdEi+QtIWEU4kHkuYQuqjEIktLZGGZBnhX808IYfL0ZgonxX21j/p
GVPN44ZiKHe3rlOTszs0VRoGyiDZTEd+XI2HZ8/VqxQQRiiXq8nDxqQhNA1vmro7PPjAmw9rrBCJ
aqDHJwf1bp5+v4S3mNPUS1lOdPNSWS29SoRLP9X6BVb+utyCgbNjT7tsVEpO5x7mB+3wyg5x3jvr
s0ROabtxRISK8KS2mOSataE1aCIEYOKhDr2QNn0HbSYG8hNkn2XIvB0zRmS6KY/kHHoYsv8paPDh
d6SAwFOQR6H4jv6i2na0KuTj17ocd2jeI4cjhZtm9BmTuBy1N4xFQPgcly3YNqz2UMfP8+PNWIp8
dIHGEG91WOIUmMPDfs2JsllWqJvQ0ysQrPDXo0S+NuyRX1B9vgMxaWmoF04G8tlvfw0rtPHoECsd
YZAf3Ewwjp3mJTIpXjTR0tAcwqMJ8E687xpI7Tr+gg/+kvQuOIAemFQN/3lKuX2nOLykndev/QLT
Rj/5qc9RMnk2Ap2DBUfzaS5xFWwOBjbKI2LzQukdLNcuhG6WdxLgvE6JlnwGRhUfWEQ1PUeu4fqG
2M2yiuddw1VumI5UUEn+wVKawxtee1c/JhKxvICFelHzQ2hyURHdwVNdpMRnmdEmiyAqc1H7czxh
QSVIb2FKOvuGiRVWTq7SdhlOOuWmgkvXQoNYy0GVDhiekVDiIjfSD3ezBRWgZ6x4jb1ZUIQop2Ee
OgRjFGlloaCSehmwaJo/otanDL6IU5lQsG3ouwDx1kS59pr1Xhz45fuLPRDLEmgwq3mv0Mp+TYzn
17gFhEi7s6a91A5RrVQGuU/7emGdlkAsSX2LetwcEtrbE/KbgSqmdz/GMQKLUNoXwLZLDTI3N9Am
I+5IEgsOE21Us96AjE5CH8tXUPTHKAVPQ9hSaS8mHyvIbwiRAC+Cf+W54qDD9lzQI03zWkexMK4L
da7hU/hmhQP2U4a1jTapFiVItFVMF/oMQM1dj4QQMcAjwBKe/97C337fJ8tl0ATpPhQznihNXmOg
eHIjW1bIndH1bootly4oMWAAZ0iAKG2Q9ntfWKMkbJgFOn6jfW46bAW8Ux1PEMvWiu3xcNxjqE2l
HjsC5wtYWSx+i+/bBjchjl+HseO+fJf6YQZf7H8rFbDg2llACTjsDtrbIkZcuJI6B/JsrKR3eLNw
T/0fRyi7GC1XDrbS7ehhEroehXCKOAND1qn7hd5l7ymd+74mom15ZlfR167nQmWzOPlhlhl4rv/R
0kHpoT0UCVWRCDyAHXRMLp/FTJEHtrhQOUF4+RUZ7ugXbIP9yXc8e6HIMr73tQyPrIkzFaJBu4jZ
JnsV5HXtUqMcEA69w5h4jCnY/chZfeWvJ8Q9D3qNp0YLWUE9UaiYmmLyPQP625cxZwFZQuz3Rkk6
OlnoCIEi+FkF31aBtVxxpxD5GleZoRJWiX9UB4NWGEm9wnBPJiZ/hg25hKnJ2Y8XAHwD11z1CaR6
u1OL/bbk2t/sP3oDMfgy3OJV+R00pMa+4C/vO6/2NpM/pB35eRshovlFG7nAfA2vZnNiLiaMKPDR
uhIFPqDDV/0F/o8ydkH2vw2/8fsBuqeaL+fcLlQakI+X1z4hUWipM7otSePMp/DVUXpQVxIogmCt
NahhWG06v+Sr2m51HhfPnzbCp8bgTwuTapAjtDrir7jBrYNtFZXnRfH7/DTVfzkHPetX2VizS4Jl
GqKASo7QAaWTyj/5m7FpqypJMRECjyxk2gLbpS3xUrTHNMi5kp2W3vmysF/66vxb1BBHhXsgI7a1
Ba1tc7Zmdy1+DWjWTihQ1Wl2pcO3N2J6ADeL/L+haIwytqgwjLakoy70GtJ6iACkJFB8epZrVGcy
d5MIX4PYlVCYLhasmLFhOHUdyqkjtLc+0QeVKhAgarF2VgeQjmh1wAKRndbbsNcg+lO+MA1ggZ8t
y6WUKBOJal8pcZCZovw4DK/2RPK+yVtOgOAQXHa6maIymqpOljY8fDtCOWfyO9n6R4qlLySHr2aC
/HHpxInEvcDGiEakRThKqh8SsGI90tr/nuWMGA3J09WXgKDUogMTfaG20O5MYP9mNdtvzUJmyNvu
h54gQJgxNagQ4hW3nQV+XP/jKDL3941R4I8h4snRwYeTieuDkUN+FncrATZkOH4Y/o28nNEpWQbE
sOq9JuqTsLsw5a/kR6iXQjgupkWmM8IC98ziyt4zhDSKLsUEAIXE/xN8d2WHrHu3dGKsytiz1Red
YKNR5hWAd+U4jK+LImH/o6huA9ZXPA/GQRtJe7H9Fyg2Sx0QDAU61MOKi3R3XTznhjNY6GtIhrKr
6uFH+XmPmUK/F4WVVscD0WAGLUY8QjHwH1xOZnqEtBML815rxm54nM0lJyt3iTUc/mIchPCQflhC
WnAF1YsVidtdybZb9crrr96rnBVROFehyqCoDuEXqp/rkj5WbI43FIUGWy29peHSFVfDjFTpasKL
uMu0X3eNJLYIRAg+vVPsScsnLp7BE/0alIo3x9HhgcoEsoBQ10FUt0oy1Mt7tQLENHSDifIpaGeM
+JuE/m66KN+I6KQGiuGcqHFOmKz8xrVyAHa2jagxDZ+/BtQY4J1BiVnPemM2jmC66UmoU58VSVWe
1AsxA/SSRdQHLGrx1XBBIDSF6D9/EXz15ZsRXijFkJ+ot0xfMFBN3xFiPH+GCQ+bkk4cBuaslZe0
44crYe+eZYzGin30gDGh8wKBCLgOSUf/UN1bNJsN90HrXyzTMXT8ZmaU/nV3O+PE2wMmV6d0mkfA
yXp8rSxol6t3+XVhloZbZClLmOJLjeeM3g9QY8r8JAY3m3gKIxnFtjxdNJSf2PaTo58F8MVOI2c9
FwQBRtDgBqw4/hs4AWKI0tqLZ3grAqMrnw81MgqQBRo6lh/qP0J2IhwCckzr/2bi8O0QgKhYkhw6
Jl9lvFbM2YADnsUWmkjjavgDDgn7FdMLJwEyseVkb/T1qnIgkRM+BipHxPnAfb822CpMX3NCk6Kq
yo8Z5OwrwXU4jf3RUVKGwp4HeZSMWmkxDXF1W5WdyTbKTCRWZ4krKNuN+W4OskZ/fvdyTMLsE2MS
C6Gryf2zokU5BECKD9GiFxm0cYYFMejFwgABL4MRRQMT98/L/Bi63dIPz2XJQhJE3mf7TMpj2m4F
REsNTQkIuH6fMWz5RQYj19g2hJjqpQXplQOf8fBcwU+IdGmxWt3okC246907lsHMYJJ/MD+V8CWS
u/lwc80L2S1Qb1+1dqzSQYm+TpiCgMvW/Ej8Z1YNvpwtNseMYmQkYMg26AjMWXd+SSLSBBLOlGre
hk7jQwrKrwXM1YlfeCk7WopEjd+ciTxHkDlDQzZ0gl0Y420/lil9oDDu2GEAx1m6wJzt/nyEUIbB
fr7wloA+vH/QJlDIc3VGZNC3H6utZG07N1uSFGDu1nr2OX6xYlu4E4BoLK/CaOQ7IujJWAEXL0FZ
V6syIY0wORKuitzEFo5ETNKTS0l0Q1k9qTF5kFvCcMMBDlmHHbEpIBg6DPuVTjvQmivS8YVNUS1K
PShHtd+8AQy9JZlc9A9nKkVt3nAnAIUjrx9wQhTHQf3SXF/1Lwbh2uZ0pIlZ6Qg+n9HsqUlwXlL3
b/ZCa1RpfEUUnrJ4/vFKK7EUmhNA+OdPtbOqJgI9BIsKvuNd+garCdlGlVfm/PHQMISSZyWaFZsj
eNzgMo28SlCC9RB1sTtwAuz0DTIwJiyKElVjoydi9bm9XENpCLPdeqiUtgWIfJDb3c63Cf3Bua1d
IcqKZcULPpddOoHovWErqLmjQqacE3wX7EzxqpD+cX/H1au0s1kyYuee5Gb9KNbF4/S/FF/EY645
SQ9T6otaiXxlCiJwrbAwh92oB9xvQyJfhADTlz8r1p1D3wuafGQNfAgzH51jWGAoHAENslXO0zm0
MoCtR7pQGIDNZ5rob+8yCRZffahk903+b+3ubDVMSUW5xoSBBR9ul8SkSA3tQaVoYajVT65xWMYM
JLgu4uNsLAh4RHL+BOXA90eKSsx501KTShlFCoe9KoLFHHstRs8mQ80lPnHJWC100kw9laLS7rhk
b51tMYdF1xasC7OItdaeYErTIdePhiVK5Hs40pQGEvxMPVoYI1f0lWEyBDNwkNGEDuJVp5xDiP92
nToJrYpwS+CFZ8y2AD461Dxgy5hIavXTlToA8h8HNCWz4cGiV5IHsNShYXFkTMm7+LENrDIO5WQQ
34QnGwQSa2VJS8tlm/E1B7nEeQ2IwPzmx0zV/seH6sOXI1vzWVdEI/XhIXmtG8vZgHw8vXHYBvpf
SWF8BdLw49JNghIyi8I8KUCNoSdE591y5z2fEG6Hb3NP8T7r2BS1pf4mCvF5EMF1TGxRnKjzESrG
24YTg0fJw/CDVJqUQLWfkymUGNM9G9QtS9Mb3a7G2Gm2JymmK3jKYPkeiIeOg3T+sBDW5P9mhgZW
oUjqht2UqFzUdb10CP1E/rcbPupHxIrhPMWQtRcD9E4tvI+x3/VcK3w/ZyR2kF0ARa2/XbzeR5Ik
2Dt7iNZV5o533aaNKApQZdOqpt66xz8kPNq3Vw+sqVasNp+YzmleUK+1Noe8e3qColEsuJ4HDOAV
5z93xRqt7kG/9So7JbUPN1xXM0nUjk9uWrSrL0g6rdCZ3gZwpasx1P/V2Sdn4fqbReBZeQZOvhjY
28r4XgdNb0N0E22WEoQhQmsWhK48PDr0Btqihudc4I5gkK6qOmJWJ9xAhVJ7pjeXUW0nruhadfxX
yg9UPILKpIylzdYcEPu7ax9/gfQDwfX/E2Mydkk+TqY4P7D/z9OHw2/RyWBVCWR4yZJ3FKr3Hbpq
ICbcD/ji8FVSxNztVOottbXWK4hK7VqX/KdGyxwRnL0/Vmo8uTWGoFpcwkqCmb4a4xeBN9IV7mXk
TBlKOH8GiGOD/nCUuJE18SCIGrWmJC00gHT+SnEjYR+V18h2LO3AV4KJyOZkeu86j3vhfd1ozyfR
AELRK/eRHOMpx/HX78vQkQ2RaeDVSy0TaB1YBj89MsEx1yhQd/B+Kr2Vc6kEkgzghnCBFM1JNPqs
eTiCCHHhZbiLSH58v9CW0IpTOUBooxU+W0/o6RVgJPLSpfiroUXOXlbP/n8RM9N/cATmuLh33l3m
yZzpRHpvTzIUagvDgUixmUOVEZFBKLWnPR+xT8mRSLXc2OA6MTLsKBt6GF7m6oyiFYMejED+MLKl
gKK+2FWIVzd9PFvKzGWGl1h5teZY3xLxAzp/c+D1k4T6D938/OMpZzRO+R8DbVmTUORhNDiDWhIA
y3tBUDAuTlBb/3LaOQZ9juwPkZE9jEv/lTVTsAV8rZKs4tZtY5O73tZTWCvFP9YZ06Jp9Dws8LAv
mY5HPhv4Hl6jhaw+qzbnPppNFR82aSO1FJIOvLNfVK9AT/J2yTAJ5OdIujy69Mvlijsni0+gffhW
fm0tBMlr3Y/vReUpN69VcdSOYWjYUjidhQfrWOvC2mr/bmN2hUcIh/SVI3Yk1R6RSMwLI+5H3JYn
7G2crCUJu0ellDLyrVIYyWU+azYlcrUN/qfQ/r+lXCVtX6HlJkSzSwFWk706WSTr6Mjyw0QX2+lm
NID8RY51lb5eSimz5PCsmEGS45BF/2E4op+sfd/Ea4jcY7wfBE8dvmf4qkq49BYN3Yphas95eY83
eB7EH8PEY2Z1HS1JmxoTuQLpaoKhgtz5KtGJPqHTMlWZofdVDIlHRzrjakxIvpr+FxikVCaueoz1
kk7eg2qEaz+ZMVEUfo8LI9Thk/JdZlZz+Yte7tjEx1qmmynOMnzX6OsoK6TOM2ukZZRBRu06aWJw
Tp3JXQBmwu2e39UJ34v/qnr5Ae0zoigLH5x6Vtg2I1fp9+VVtXeN6hNQGs1W489SnpMTB+MGsPWp
W6h9TpYvO+m74GR4WAWmdaiwyZoshxcc5vRQ5+2ylG9W1cozvmVLJa3afJwDALS+XUn1zJAWdRBy
Br1UN4oDr8JzXIua7aTKW9BC0cF3sbaSKg6kzwFv396kKVouRs5UxENTLaDJN2t88s5Auh+1+EXe
mNrdijXqvv5mX6hMu9svsAC6iPeGKRmHexRDZzLuTCIio2c9RZf/RMvy85J7uwN4MsLjNB/ivPG2
hSqFwL16BZyhUtnySXyC0ONZVaRW46ecN2n4DF80MUEbZnizLIzBePmUe421GTGiSvKTrj4qAJTI
IEKQKzJ6vnbFZHrhSfZxcQLsjIe31W6n/Xydm9F8vwUlL7yVl7149Bf6HrJcnPzxiQVtbOJnVZg6
1ZuqsyZt3j0wOX9Fdgi82LTN9N8tPJEgqMt/1xgRIA2KT1622Dr9ShF1j0RpL0sd5aI5+581GzCr
FNiTxJL8aBwLbNSMmtRVbWxwUYWjkF4/Ii9dDU2tI+2TYV8p5PnARX6vJXzHOHTk+NwBZpIKcOxh
/fGqY1nkVszg00+ysObH9FoRyU4eexY5h5O674Qv+kJiptGcfT1x/w2xhGe49fBAAyvnJE/F8lft
CmaBKZ+fkvvc3o50/bW/aw05J504N6vjmwx51f91HfSoo4QGjhe0pOOBTZON/mnoosNsrcHDw5Kt
zIihjbtMAcVR+PzCY61fqMTujYx/91WQV33ZzprSVygJLdvCo4JP/tjyIGq4p7QVpY+xq2wUKJO0
nnus/KknEXTYTL7LsPd5eZlMvLR76BbK2Y7HnVL5SQ7cdsRUF6wSCioRCUiVPlQqt2hCAsShsvx1
+NGBS1OE7i05EYjuUslA/PQ+nybu1nj7jYgWUR9LPTMhUHtM1CBoWYcd7B5e3dE5fxun8KkoZSka
irhHJ9yvfeoT6iM2i3dOnhRwE3qx3HlH6bCdZOp2P8DqBTRFuiQ8nVfyB2yr5m5ZwyDtR+rTZI01
CH4/kwT12F5XpPB93Wr6evE1WgQa2wXpzsXgldVPU+qfAjO30o0GEo0QVrE1H7z/Wzbz4bLCbL43
dyW1tDMyiFuQ+UdgCaZgLipfCe+6+RZ74JcjhAITRw8jbxi4HYcmbhFPeS5P+hqSvdRuV5ju+2U3
jcIbcMbm/zGu+pPMjc/a92Uga0A7cKogqMrzc14gocu33knm8t2nH6h7vzfGih8rrwEpYr0aBryH
Qd7DzRVbdHRFDpOQ8MxL9Mp0zO1eUmex5BNYBh9U+ODJafEO4mDDs7oL4NPGXM9ultEVK488T6rN
PWRs4bXgLaC9MBH5NpnBTRPqutvbDTKZxs1iQ0vJDzjAVaJBIyI1i3mXto8Fb/4KmwuJFkApX4Dl
70F0KWALMJsUOFc8ten1CHzoWP3lPBaAigtEODM+p+rIQXWgdgV6W95aW8Spdfn9oH+fgzxqKicI
RkVv1KfaiywP9NdhpXrEJTbK2Cv9b8HulGAiQ3JotYMqXReiLp/ex+ZFIvwmqTXhH1q1yqKK+GTA
I6dCkazT+SZcN6wEHDkDaB5CfIUe/66lFAYIm0sbhKsNnO2FRlXPC0I6oOH83VJ1EqmIkKgfJJ6h
T6kBvJ6A8/4k/ApZ8eI3uCTyL5wBEPp9aCyEaEcz+LSvZNWgaPtbL+Nxsnec9POhoij4Ctj8Mfar
2vqjGCwcY4IYXegxi58qXasgvacGlcYkHJpNU0ZvEfq7QzRM9MOtVFJ1QOLXUTaH6KTGXegzgPN0
GkvbgCzyDRgKsWr64lEGgIzw0S4doGP1b24erPzF+F75m/FEZmWSqoKMeqh9GeQybxj0O96vYeZ3
rmiz2WABDX+JRnHVAQzORDqP7pBNGLc2wGqF6er6KY023X3HICiDCiOO+fsyOUez62KwIZ2OwXzI
dg+JeAXLvFLu3JWuYiDEJV3idtxxiY+sIjywxmPTRJhdJo26CNPqR3CtZL6FGh7tHFeLH0Zd/3FA
V0OVB0HSlsNmeh1iIpcWg0WzjV2hBB6StQGcADxQtDDSnxma9Z7xEHbJDHtLqRtfr7+quuQcdBWm
i0ePiUVFHDFFIGRQt2G9/S7dbGHmhZEmlvwVr+aebUfF/QzZDHu+6r3Y7hOjN19XWi9vBM43ySSt
L3iglYjTRfSCZ7gbndGFXsxKm/cvX0dp9NsB+G8iR5AZopRAZ9IN9QBNw0RmuCqFPCC0v+8Dtpcl
FrITQfKQhOX66d+oZvnk28rEuO0rkeplNkBGXTxCL/KKSjFbSIo2D8PUK+uLAJIiKJQDVHpplp9P
ixSe38agOGzC9RPX3ZYNfalM24TquCyNDoviKlYBMKcSLaavYc5YEHZYpkX/FGn3KpH564xf2HpM
E0UMAdT7ODX3PY9oWhfWNDAyY2utgjUnHPHDi+oL/Z6FL2iahwjrmku/iPF9csN7PfmK+kNUnwqY
Wbj/HBOnErYrxGvHBU+nLEBE4pozshQoVXOYLAda/dz2RF1jTtEAvrK1wqk06Ie4/F/rYEealTFw
mLtI0i/TyzVosYxPZopvGeNKt+Muf69HnQHVrm1z6ATffpvSzMIqdXskqT2byXtifUWHWceZ/Q2g
aEwxIYKDU+MhS6aQl6CI9fTjI2wREnasA+zuo7BgfOtlbGiBasDEYz7sdlOxGMHyfXToWbe/066T
43Gv20SxC+FE7H0DFUiDSRozT/wlglKCgCVudk1LoX1akiwq93x+piXem6fajRvE5fz0Y6YGCkfw
ZsCBP0iPSege6F5gYBfb6BIFE3Gu2A7VQokwj3TygcPJba/koCWWlCi1f9cndZT7rfUnSbef/yTr
8PeReXR6J9RLix6SadYeGeZwbTfk0hIi9q8DNumtbbWp4+8yi+oCmfcNey6M9mRF+YAM/5rDpaIt
YYKDHUz2udvloM4SMuzWWVk5oGiAtBpaGB5cstrxs/qWh4kwEzv8e23rtXwp9jRf/mB7ZME2lpDB
QHp7s97Kr6Kmb9MtmFFgK3O+acdZwks3GawfJj/lvCGU5Eoq2R/abXta0Z5GYqNl9pwE/N9yWIzo
Duclu8lyXmO+jGV6G0xVSozznZAbf0sI/RPlAOYGPIttABhojxdXZi2HYh8C832FxvkYfmfISHea
d8ZNGMps4ZOcO8W8JqdKtKI6zE1+sKrpwUXBUniTIFaiP8iWfvKZfdCeKHoWflX7AFLnobG5535s
XEGruqYFgVXB4K0Z9H0KDZNjuTXO3OHZlWYfnTeEKjOUS38lA/z5hCl9sBxf2iJCSEH3mbtLQ3M6
ttSDEQkaY746vFc09/5hXL2tc0AFfvz0umnzMsDn1zlFw9EKQNJuiqm5AUTQfAg2K7O45JYYUqfd
ZNU0B8c/Cp3lOMCuEaad/oe4fzRj9JWZnnzq9wPLLkgJvtw3DnRWOWiIAJEqq/W/md3stfhhoLuV
Z++PA9TaiG7+fYYlIAEB2A7Wx9ZqSTXqz7AGuK4ANGue7Z+uuAMpPc8Mx5JZrezVbNvaKzHZQ5Ge
BFCAVccO6sosw0sdNbMl9kCTReel0mLLQbNTz2KkVXf3/kHN+WsMGomTzKd1kYgeAOkVSvCNPZwe
n7xqcPjD2j6avCDFCZ08k69NFokRFYecRTY0vx21rpKgWj1NCxe0l03N4PWJLbNRXQX1E8lN8+d9
DPzQzCRhZqd5Y9AdOD9ZbzcnZylUHtO9wG7uUUyA/nH2imjoby1zjTKunz5IMgYZRZ9v+l8hC3ts
1A2o1mrw0F2ZHRrXo8I/DSplk03uGp1rGkQHW1/4/RmbDq0CX7Gj+cywHezGwL/LaU7VJT1ITmR1
oebLT5X0RB0wwI2zvCrarIZOzKWuKCifZVh5y7ldQ5HDHSLC1V5qeX4pbgzuSsu66cDwiKDetlXt
f07e4C+PB68xtmEuhZoZN+x8XmWqilGppupcmYWiIEASOiJzVQFEP07FNrcSFaHE6dz9tvhJ4sch
2AliImohhILVWPqrP7wJVwg+H0sksXIrw8fdhItg8e6Ivg6/psTNxmGFsI4ooOxcSQCvxRcBJ6d3
IeDMyDNSGZJxPJQ8GG6Gz2n/zS+XpfnVQiapAv2AZrGgt4QYWuUuk7RR4HdWfegQXy7kaBrEcgYH
DTSa7EDDJmUZ+ZFlij04Ps5qCkOp5TaHC5sCLUcgu2hzkzzwexWTCz4uloykpHoay3NCxBtcyMYX
e3GNg/NEeqsfs5mUKrLYlZE66nBk4lHgevuY22g5Ceo31uz5qiVtP9xN+kLvUkG6e9RHuWj7xUld
w1muJc53sqyWObxnPsBCqUJhDCb1LKQEfcGOqDyxXG5Y/EULvLTz4owgv0ZzXrbTSynB4naNv41E
4REdFa4KQTUxtIdcrgI8zPrCL+YQE+lJHwkjgFhIhBsHHlAZNgsuYSJhUUgTsI5ZQsly5ermsb8S
tXXNafmIbYRBbfGAinWDqSVj9TmHwHihkD0tYOcrJwOJ6DEQ9Dz+9zAyfekL/MzzxjRyK4NbeFnr
giLmWAmFt06jVJl+0JOStlPMvddeHDkosWMNIL6BCSkWlmjIDtsjxPFUyWEPLUWueqZMDkQ83uXX
Q9GFoQ6mPfekZ6sg8yNlUlouFuwpClP5rrmuflLP9XZgSaQZ+A7ZPTL9YdaAgBz51YrFvz6FYhKt
6z5KBBzMvkut7ocm9KxCBBrgK8XfGzku+7/w+fJmOeWWQAPbngEKt4R8WKiGoqiUmxNHPiiDWYPX
GeTvbhMl8VX69A+ujsT5xzI05iABCQdpWtm17D300wQNw8fl5RbjzSKnitcN03UEh8wdtQ4baEIM
fCSl50ZtFYEarHCc3TYZ3Ngy19f6UaeIQJsqFU6L5O5+DAeKh5dnRDkyOxKUNIvIvcd3KalP/PZ3
M7W5/gNCU5gcw9y5KpDqsVHXX7AT2knO1Kn8o6NmB9exb+hwGoO+BiexbHtWDFSGreePjMY5OTjF
9AR9Jy0OuqA0wmGcvqbJ5QEc8BkSfWDL4m2kqmWbIRsg0iZRKqzmb4VRhvPlMHox/qARG1RLOKw1
BHDmEETMrENmRMED+rPJI+0IyI2SydgoYpqlbrIVO+qQxaf8b6wFIveNhYdqzqxYNVhIM591opIg
BJRe/HeUbmpJwX9PqcpmtmHE9wfZLHPdcAk0O/aZqIIkW3d+1A7mWOjnbQ3gxvMYw6/Lr9EK8TT+
nEQAlwR/S/jKGc1FTmhVGJiT3y7LO3RMaZZXX9qr3C3PAOu1aSWx6U+w6p/ctGxNeBEghHx6SKNf
IuVpQEf9ygitqWBZnPyq6On+2lJVYr+MgKeitzi1UZ+0dtWePcCXDVEuMEjDpw0+YaIGNWqSrbow
+cKC+lYBnZpGZL2xDQXUKpuMbwq6VlYbQ+L8wTNfXwQ/hdVaEpio3q/L2UI8VTWk4/kCqGcC3nov
qVU/DqRPTpVEeU3O172d5eSAegBdWYemO4v4yQTKVeSfepNuZLGsyDs6GeVvVlCXsMe8eIRu6bJN
N6pgVqCh1xjo84SRG7QjCx1+cqBc32bmiz4f97cZ4K7miElbK2RaNtZuzR+X1aEbneib5gRkdcwW
/fq7CVvS9aV6u+mXCLWT8y5gR4yuaFlgeTI6gya4w/5ViqvFZbu6OLh021N77+TrrHftH+Kd7fuI
ebQUFT5VK44oBp1aQdtOCv1cD6lWS/dRWgElF8+EwpimdvB7x3PU/MQ8xOSZVq0cN+0FD6ADXmrM
G8rQ71Ycru5ak99FAnP3wfKUKJ6xyF+3yhiasuFtvA8ZD0IGhlM/F2P/pj5CH85hbIOF4LsE5gZ3
McEVsFanurCyA6LqWQ1bVwgPeid1PYb5GZkNqUmoEKhRnZzo7aCAYCw3pJtwcizc9sURLAJbCaQ+
4G+IaqMoK1lvnB1N/aj660hvXALYs/zDJEVq/T8U4iJW23GeZjXTfGvl85OCaIad8AVKlFcEUAAS
ZiDdFOlWHe+u+7K39yhNlPcBTnTqeBMRNL5E2DPg81OdANlL2IVe8czyT1zGN9UeDGzLZbSWV10u
zFpoJ3Hxjb+ZBLQxxR7xVQud0L6it607USDf+5hc20hIuVGkqn7iiIY9/DS0HpWq3dB+zZNEk0a4
iDeEUmQonxznDTWTdZdRlsb1aIV8J+YOjjrTrJLVSa+szOD9/yUR04XNCFvRo5u9Sz+r0XB2N4QJ
NBr19aN/8Js1Vr0zJbxGo34oLlEnZaMjHpsHcPLbtaE7RSBMoQk/lyQgrIbB2ws+uptidIvicgcY
ZOm5mmnEPlUA+esEKa4nvcj0cj0DQxPL9JD+YPx5RFlJ/ViVAP+l4hJjF2nVf414XJpgsLpyLigH
DV9MQHwpLTSwNRNoGo1hzerRZqzFOC/6cbfFjcd/K8Z46uoH7U5QZKPKaJYqGSfuR/L1gVPu2EC2
5gfyYmDUqN1IHW+4H3r3Wlhb1cSqrpn9oqCBp5ATrwo/zBi4YkOevPy4EGXtMAFvntAJqmguNm70
atw9jvyc7g3g1GMZ47j9IoBMuYz9hiPTuLcqiKjs4+MnfYp8e0G7FfmVhMb9W4arRWj5bj8aLbuq
urWhGNx9+fkOLDgdVxAvsXYpD9lH289swqYIeGtz9dCmsD8oPyPqjg9AesLto+TFxp1Z8P6m/OcU
v2xNkqa2WqmxwzIVZBXmznvoqS9zGvO/8oAFIL6gs80wbEgPQ5rvl1mBy0aQxvS9ULW8WpjLyCQ7
LOK7Oxsw93T5DvTdgG5zw7e6D1WxMeWvuvLQ4JrR0TuMHxRHIJE0DAKFvivk/QOgy8kP4D+xzghV
m160EmX8cBKr5CVaJ91ACKY0Z9HPjwGAn+Wb1MPZm2ToR2ee80ErpMh9HSII659E8PHAUyt/2eJ7
OpaVlLvoSfnawm5VMpe+WoV/2C6G4ci5JBF6FUeqpEH0ECjAocT0DuyPbDEezNxXy5TeloNjusqq
jndGTlmRYa5nj/HWnff7uetciUrc+OIekUHIWUbzVdCj7AhZlArB8Pz5OU/WyeC3PWWrwC8PuIoB
e4bSCV/iz1MDfDQ9KzWOJLDSZSNVnu3oQiQbGalIb4uiSH3MVc2q/7MkO1veqwPV/U+GYeRZ5ERp
tmIjmA+z+gZ2xhqDji+IT/2+7N2iLbUGk6Dq9/fTMCvGkp59Nqv+yb0TdKCmnqUkp+g+85GMy2Lt
G2u03x2Zax5Ht1W1YILKwu2tGnLOp2ap49tVUH6LLZP8NNSvZSiDJyjc2TjHocV6TnHXKsUw103d
PH/ePRdtAm/A1/SEZXg2RtWp9GqslciTVdLf5e+PBuun5SRy4o1wTdnhoPzqgRndYvO5StCD4oSL
VTgzkTHNoEkoVWhu+2o4YKbXSH92fZydoMCWvct8vC41qYJ0YnzBGg3r6tis48XuySdr41j6Q2i5
iot4o2CJLmMLT3xzehAioOgyPmV/ZdfVyUEtNOo0547jY23jkl+aZJOG7Z2JBODMbcyvvHtxoU2w
kWuMuhbBfU+66KQcejM4CyUfhF4gbLSPrLz15lpfBaSWrBmRL9obXGU4OZVmpw9+s98UKkzDB5/f
kRSXDw82BjHtOZXe94C65RrESfH1Ccyk3RR7x0Ril1Pq8o/wRXGZBra/LrSe/e9W3jvdVYWXE7TM
eZ0wyqwJcht298xEVco3rnvg4mpFMULZvBen4/+NGcwfBlfWoWUKLq0pzRiFxtXHMjCtSVCh3mCh
byQHoVIajxPYiZbg4/dkibxVCOCA+yy0zn8NBkAVujATkQp9G5nqWgO3oHyFgRQ0UGidoHlirgUn
3D4ny3rfO0FPsjMFrGurkPeZH/QK+nZOwcfUhwNz9fkpwpQj27vj8+yaPwfEhxS25jwIs5TWCwc5
/VEXefS0rxS1th+Q09NMH5OwtubZo1hhAttEJOAFR5oRUGebqHYS3oYGoNuviGnQW4gtKvGVZlB4
dv2idniK+wOy4AJlTifxNdCNb0ZmHRHt56UaybtgjNmAKrMAqb7SPt5uVdGakF/q7S+DGJtsRNUT
/q5/Ts83RENTf122j6ExSuOKSzbpPbN5JB3GORbz7kldU7RbFTuhCBLn5HoESeRQQ/4PT++QkK0g
eYmBKJcJFn+dYrSm6Vx7qqgSvQbelwwHfUj2vbxzBz3P6/PjfwLD/T0kr8aHdGDvRxGY9DeOtxEQ
51hhISCkGMnyFynGuKmKegQE8LEP35AMeBSKTiUhGXbgXcTrE0v0s8P56/JOR9nzLl2loycNOYBb
/dQalMJLDD5qfU3TQQHOmYwULYlrcXnpxQCmyqLItzMVg8hJYJnStN+1UQXmdhN1L82Pv53uA1P9
ZoRE5djWqmsfgF+tV8dD74LVgfwX6DAMdhkRO7b4ZopRE6qZAXdPoyas3oBO/LoPRyPl+Xzn7kr7
5G4Vg1uokxpk6nGtMh2bDwcBB3sD+Ee/SXGXANAq9DtFVHjcMHw1mciFAlH/Qf3wIdq2UZwKwm9t
/60BXme5YfzV47zL5ZtRSccgC3ZUMpF0iX27hhMafZu9KKbBffaNMvY/u5fSWUX1BhE0JEDFSJt7
aMb6n4tvpDOEHEbXhbmoqw9muYt1sgH+DCvJpZCJDfvMkXcKOe8NRh71b8UVAXKtLcmk9oCg7/j1
PJOmZnKqv21DRqQ8bKT8ib6sQ5BGM4SNIMMYaOTtsNI9QRbdD+UUkSDQTS1pvlh3+CphRwHv1Fa6
tGnOzbg7iOnM4wmjvB8UU6KC3jRYHPcQYeeJqsp2eOPVprcoeWitnJNSshvbMO5gnCa3kyF1Dkb4
laKpRWYOsorv+Mb3wSkO+io97gkC6saYRIb6X6jB8Mz/vn7AA8jJzP+EDoAiW7pYlDbRSULve5+x
HJbI4/ZacbzFdnXGYM/34i/jCiTXWaouoSOGvCM3qNNYLCR84NXqMfOu8boMYtAXAW5AJjAjSVRA
S4YAAlJi63Z8jLK+EYNoGHB9er9T/TWtcT3CgKZI5kAdDNAJs9PwSF57tZ0lJv8Zvmi6VKfpkunt
H5iNg/Vq+zHM8ZtHltvDxLm6s2qKEebq923wXUBpr9HQS01dshybpsfLU6SsfGVlhHzwGQrtX3iM
V0JIQjU1jYHegqzgwtUdLxzRXIgiTWyLp59oWnEyNFCU8palwsTbuyhSKRNmwELuSPRPv+VDVQbt
PMJ57f4dV82BYgO0lagQSCCinjzgHoOMsCcqg0cJPnesSMzWR2cKBTOdNjKxWqMi4mbPSiqrb/z5
xHEve3JKQeUOvF1QznwIcsT2Av3oULskl0xjAAH1MlajQhVErCJeWv7WBc9xv0NXAj6bZ5vJn3RU
iycKoP8H7T1UgT/sZ8O8UncRtbPQVNAeR6bH1e3F13nuY5GEQd86GvDLRwGC5Q8qTm7QFQks6vbo
b/ECF9NqCOrTZ2r3/IXAkJ9cqaQ1mlYfDtqRcrLNS1a15Q6JwM5rtIIOLLlai5ykwI65OJfqMg4f
JElz4r1PGdhexE84sPM7jFHFMnDvWwi8b0Hn3d4IT5roKAmdjxDQ+VYUovxkcSN/DbIdHIG0ta9D
/XgQISBGxKFcfcirA25SbqcvVxozi+IYGSaoLNbl83HT4EPrWTn2rQesvQhEFLosHnihwNLX57Bs
lNvSiFVYBu8C7YZRIxykJVNrBSuSBp737KKvjzvfGb5oqVicbFiw/HhxXjj++W4g3OQ1NUiTJlZ2
1XtpC2H4ByFDzf7TPAsFUxUSMrPdSi2oh77NtSKHlgaAMIOAcf+iUw3bC+2ojyNT3dVFnOsqD0nS
6g4KdXnnq2LlQPHGcMcarVdMSYvia3QwM97boyGrmb78qWnFOR3TldWUYIGqdZmNB8hdeQpmqpEU
obFM4nxoFw5Q+6jdTBNQeXW4dXQXRbxR/aMvIzeyd6k4p0x6upBEQQosGt3eReKHn0/Wn3WkrhrP
2yPm1XDrWxbd2c6Vgzc9ky2YV8ZiAahTUlosGsEjOxS85ZHVOGHymeQ1q9XVbaR2tX4wsuNFakqu
0KayMIJ8gknABT57RLPmD2O8uEMmJDeCHfSeji0p/LF8wcXNmIdup43Mmg0HjuRJ6nAoSH+dHils
O8TAQbV/WoS+Tr3pDdI7DsL9fD7jrmgAMG8T6W5JL3fUWQ0+d58GxP6CNfGXD4hrkeSVUsesIkWV
gmJb4s0+UBj1isLGIF1GiFQ7C6Yzy1WI2hpMdp0mgrgocKxTSVNAYGfI6pdQC/RwRJhn3+xlsUOb
n8KpyksKjohx6WYd4+wSlFC7ax8HLk3Zm5nyrLxsYR5L5aIiy25HrdFBX4jt+ozeRoJo9faDbCxs
OKxD+YCZQD+NHfhw6Y2BW5sYcIn3bsf/K3WTrYOew515AU1EraQkBrIL8bBG5GvxID7Kxp5MiokH
YQHk2ATztW30Afr1tuKLUKYHssj9nA/sqClF8aFRL0MY7iu7qIdF/0gxumIBTWLVjdeoNH6nINtk
30RtL36ejuPJSUU9jVC1jBghOa8uOzrfUeKf8+zZBHA6AfC3Y1zzx5Ge1zXyw2G7AOztOI4N62I8
OWWv7q1NKC2+V2buXICHCXGSaoTs05MB+DjiedZiK9d6TzIxFMlcl137inVtCDWBUBCbkvQ0gt8N
WBQjlSGGjYHNYQTctz+MxIIH9LBzGVHWK+LjVhrHgvXWOaB2CE+blmFjwyGLJ280zea/osblIQmc
tsK36x4GqDe/JaQep8YBZJ1JJAI3gSPi58PwUH14aRHk0C0AhCZt43IBO+AhmGbtjrBM3E8iUAUi
WDUQal6UZC+Nr+h66GAXGeBgGJmOUlolJV0Y78AELcDWghZsn5ERO6h/ctM5qmfYeoPsxCQrQ4gb
ocmbCtOt7RKH+y4sLNO6iJhlusar1bIeYNCqyVsfcH4sak56jQ2wDEBQVdXeg8U7dhph1iDz+99/
wyndQjfOimEHgthCexfx/HkmdD1c1bEJUMibAkrKI+P/0Rk0Hm3jgwcbuBM/CxyX4eeoUKIWqm4/
DBTPuq8ZwzHoS73w9XFgvoFm5nJz4WNdjdDWqTGi1bvWHTjRMxr6ZBTJXmT6vwhAb9Ll4KkcJv+y
98Yy7e2ocGN22z9TpXriPj7gFJ8GDvZCLV+H0bsDzKTYtzxdcKvM69WRuX8DJi1WDggsxk9FS2r/
teY7pz3zSJgJgQTYwwyfwdJQG6mXs5Mp3mHoVJxXTf26/qcLm73xr0QGBEP7C9DtQcsg/CUPfJuS
MWvN+/5SoxLCF9KKlW8hHbyBBs629bfRQOZtL5CHfvzG6yE3qvKuZiM2LHRVJdgaZSGBVJXs+y5U
ffMY5ijOjnyqkIBSX0OTdFWSHy55w9QKGZN1G+iL56d3inuvkhCF+JIJeFQqvxPIg3EWWhGt9wYu
Bhs6MCrkWhA5pycGgNMCuvHizlNHDMi92LlWsRcHrS+L28Ifk0+YZXPdNy/FzbeTqwniQMN6k19w
U2WsLv1MdLpAaXiviLy9KAMvLCUHnxmpdUtB8y/0XdOzFAVQjPGEHeWRivDJvF/SX8xURwovOLqK
EgnXTr83MG83j669mREPKHU7jFQ00XwCaxPBcGxnBzB32zOp47zaKbhhDJ0npe2+csvWWpcHvq0a
lqM3VyPLbPylDi33q+Wv4F8DZNcUKjfhLIwAeWqvFHQEslnOd/N1DkXwlWouZxfB8loFkfWeh2VK
X8vgz/osCBI4okEe/PLAnAhmk1Z1ij6IlxaTdMlOJy2O30ZKXsPaclA2kZXfm29rAqblKjnF2gJk
bmwzSqVtwq8rH/yZqVdfkrhUQBTgVII5W6N3QbjSCusHuxG1joneatKO33FP+WFfkeuvuha3p/io
B1UlCHbeoN1/ZuZZr1G0WY5InnpDdFcK9XZpL4ikYN1oQx1Ut9gHjiZRcBnYdpcEckDf1WVbog7+
z5SG8+GF4stSen7jSd/5Ya7mAuG0cxAxi1M1Wy5WjJgJpVDK5lOWe4ZPzkIA9CZiEX1zP41Magz+
MbE01DZ/qEfHzfBefRFl4brfY6x8UrGX0hjiE51gJSnYea5+rk4W5FY8uyqX32r7hav/kkU6ZT7L
7RE199Ov2v5B++zTV003VWLi5ppU6hRFd1FQZ1xtUYnfrlL3/B3n6K58n8mZxavpaTWQ/PDj/T/j
O5QAWPD7WT9Sq8G6AiW0URcIGf1u+eWbD8Vaa7HRKm08q4sUmKfn3m/Jsvhxlhido4DhW0x2pV3y
15otzl+dK8ieiTSy3bNuH5m6JbpTXZyxcW7+emWhhpIQaila3uRpiYU5iXt8krWTSpsRjA/cdKJB
sTYiXQG24UgemV2WVFqhNr+3ra6lUD0zANI914vITKcpIjn1cbd5NfSyydN2iQvVgDi2S8qn5IEt
RV8yQFM28YRVn+iOIgtcVjOiWIs1liQLMj9sM/2R4z17Z4qQod/VGAMAl04kn03Vtz1RxpHoE9xd
2Q1ZzkCQo7viDT7Q8l9nMUvZLKXVhDKNbqEXebjA0QQhtyQFWYgt4FHq7BlyglbVX7olu1wYE60Y
76oAparCQFpMZnK4y5MIyi4KLL0wCFuRrGZYz7i4+edio6+b4vYH31pqq0cejte1ubkPQt3yJU4E
z9bEc3rw8/XhLD8Bnvam2z0EXU8RkXXtK+GR8uu2QLTu9RcFNcHcbe/D5l4kQ2qdDngAkj69nQL/
vaXcUQbN0U1lGTI7/iMo2qozLYCyXweuNHDayr9v9kVao8rFAz5rl8WkfQzKhyMfJchRag5gPHVd
k7/HvJcZgeinv0mhLLQ/zx/w36xT0VuYLB8qBSqkNvnyivPQzShbtOt3SIcXMA76b1wlj8j/tkyl
resT4HIuJci1o+8S105yoI+LB0yGoFsx0sP28pn4yn3aOoqh2GvpoAXnSmz03dcM5OLRwRlW9/Gk
mEK1yOJmrTEAyzbmwJvDzESJLL+QAtDIlOlAxP531S5aGficwN0S4UbrdperhgbBsdWWCkIIab+l
BWE1EAKzoTR0XHP/5O674A4DihPshRLgIFdB4ZOLO2YFNBpjrK8u0qVoucrL4/NJl4O98yvgiFKI
i3hCqcVyr2eCB7s2zKB6zQasX19yd+deCeAcTrYYjrTHFu5DyO/f3t6J3l3Tv6mQM0gJ7FtgWXzp
XTQ1CMHFJiGBc/d2IhLW8sUazR99Af3aE/EJpt8RdeDLoKmsIA8BaHH6/zc0chpb6lxpQLJvjpUb
B1SK1Z0gjS0w0OvvWsGQEuCddFh517U0Yew52UYX5ca3k9R6eCCYdfU9ZKMwVAH5adUXCFIldCtv
zjhTKAnuLqDicgRfPMMCLVqKytHhPOc4rFWsYgKLDZgsXbwLNP9f8CyAgVqwvO22jHzdDhVjWzMw
CGe39/J5PVzOxtgrCGS7dq6BVEacbyLqxy4693G6uG3F+CaRMLVI7MWZ9GvJ2FDF25+sj/iT8k70
L7YSce3jU7qh+Uomnxe9rfdRHLtzKLo+5j6khxL/QzsTH9St6wbxlaMoBxunAmM8vfv7t7KeRBZy
geMCQMgKG4T62FOl4gjzqBjfd894YLPl/bNrPJTjUecwGxnWvOHrVyp31c/wVIbUiS2N7TBeUVCI
Fb6WOweT2y25Br7Bbcr2te8xL0EDZXQF6na2vMpwzS3XbYL9uS2hFLahMOvuosSBM8u/kA6oaV3r
tQxFN3410u2PkqwzTfJbf5sGnPoZ/G3rDlbl3ldj6uhPqdBTh7Yi/m/njr9j5Etr88Zc1taJKMLw
J8j6havtmLFi0Fb1sM83H1xam0+UZ+3juCvnNqsgYkz8ORf7a5P7Youent0mQbJJJSb/MC1lMWEP
r6iRJSKAROcsVI+AIrFuAOMLAxGmuE+fW7veWLuI8sMBCzz+M0HC2kRyQvr8R2KMXUMr0hrTLAoT
xqP4vJJGTpXI25kv5Ae3Gw9tvssGMoalG5thLyW5GSfkYw4gHRsDmhF8XpfaV+D6tbGxnGSeZbMQ
zS5xTYRg35pZAwrVNxVuCfjH8aGqLRVlHd8V3g7NLeX87kP4qCoDmbXWLKoi89eZcAa8OnscSxhn
W/Rx07R6oL5U3atFNZkl6cNjTuxlmycqbTi50cm36rpUM4+XDElxAEOKw/il1/u1bi67GL7eacOo
GrCc+KC+gOQK09M9k3yHz5xKlT6hmYfeyGzV7V2bY7lQW2Dq0NNFA5jx4SkjVcaLBGztlCR7t4VQ
r/94sbDwqc/VF34yhjc4an264y7FVJ87edFpCReYN5KOPBGhHcNrbZu4vke1cm6Cg1CMtMVTwagE
zl2NVN5R0W2mgHu8KXUsUQAtaSHfLUDFGkGyPmsKRucC6j2Yi/xumPbVRzMw1Lgra1kBb6nEcEOt
Ia7kKQE+rULmyJDdeUnRhhDcm4NA1qYd1Yu9QGaQRqMqCRNTptftsMm89ECc9KDnLQDNn0sgxp1o
SfI7usDPYFMKIFDJ0XaIN43bXFeRT1P9q79T8Sbi6DaYEQMjKsaMV2W+kGayDESafh9jPturolDW
aVphg8uDNZ+CDAYjsLStrkSpUvkz4L/6DpsSdqM6Q1fV0xGV3G0WuDNpKuptt8d6NMHtwsbljKq2
ra6+mlW+mYPn0KxkvAnrjW/URIJX/8KXkagVqkG2s3BBYHa9aGn3owunfbDjXn1T1UQcxm3Gote8
BA0LaDKwkK7QMcPWV9RGltlCxPuUc72F22gOXik/WYoYqwTxdDuf/hNtQTAzxrzl9jbWNAYnLA2L
vjv/Vx4H8znW7Sx4Wv9mKVAiWHg5hhl0rvzJsHAyw3tHa0peVVwXgFli4fZOwuRJD4CXb6HqWEIE
sXdXslPFOW7ZWTuJufw+/UQioaPEC46ctDLzl+siNw0h2e2MV06Kbu5apKjIidrM9IFfkeNBbxGs
dx5tqNZo9YSNW16p61leWY0GMKulWbH2FhmqvgSgYD98t64sPaj0T+COTQ5RvftJOx1Wc1i8rdWf
RitwPO9ob5KuFzUf47kvWYoxWS6Cg6xWWOEw8KVBiVLCS411Rb13636VP0LE2f0RLf77wePxTgrL
QdlpWC5dMP58yfQS/sslzj6gUzKo9AZhO15YaITt8Z+5hqGk6eyjVws76xlisiqEMP6UyyF8Eun7
uunFKbuxSxdmeFUZj/C3aBIh/lMVnL3tWA4CeXFVbaxB7T+q1/vHNajF/kJkvyAnK6var/JXVzmn
kkfEY/v1r/Rk2jA3a1TIZhHd7yp4FunhBnxc7W269N1N1w4mfqrKmXymzqSnXlL+2tL9UI7uYudi
UXGhROnKrh80rNPGPYnXU1SLXO2nJy+jtFLJ37BmA6rKFOEgHJDqBc/VqRAKUjUVcZ/vsR4ScGQH
ICVkFiOho7Sfpq1FOjPcaiVty+1p/haHQSxq6u73YXi7WTjQ/TK6vRmL++Q1YO/sjDmv48hk+cwW
apSa8FyWhInPnCor2jpp0rzojQ6gvlaNGzzJHpCGXGAJQTOUSSgPJzWXcweQjLOPaZgJGtg/WzRe
M7AL6af/e4y4clahx8f6ipuF0JOUgTScCi5Kk5mkGUFCHAZwAJXItcNaFLjQmiduEvkU7K3ow4n+
2PBYxySDVpAuIPPIb9YhTLkjIuM3oI0bw75sU/iquYx0pXokdfq4auDGW8yn1+lONPO9ZZcOilgR
B1Y3kTFpr4Lu8WRSvOJyITfLMu6xcS2O665Cbyh88HqRCPRP75190Xi/eJxlw+ivZGNZ/QuC5oLq
X7Hjqpix/C8YlCJvAIJwg+rf9T77zCkG+PCxdTMsTZTHDhYtjqKoDM1VWnIEXyGjRV3fKp4hp+zA
YCIX4Eb2c2XLGZVKMJHT9L5vSJZUAa77c9tv0uVJm4gZv3fEiVplKTt+Vd8eUoVB6vFmksYD3Rxd
UQIzD0wWIvBitKg+BVsKuJLlVAY+XC2h+DNuLiMK1maqrPrp8XHIPUYIJJPVkXGOhSSS6wF4m760
bsfJXeJprCmu9Jb7JZmGtKFLOhlfIXK5jbvBxR6mBUjLoRYSSQ7Ziw8ZHBLflihJ7dFM+Aadu89J
uJFWBpwYGu9pp8/nicoDFPImRqeR/n12IyL+yMiggPRSP2m9FRjnHoeedNMBoXQwb+q5agw6bnGa
mGqvhpIm7j22fFugKe9HCW5TMtYmIP9UqnOO3lL7trpEwnw8xBHtxRocat1hrZznvwDY3uofzr+u
pvbn27lEdLrrPBFFzbvXZDfN+Ydp+tCJqRAKqTSsuLOk/eikQ9KNW103cms33owRfMM6Bj6emK4D
v6EmbJT7cEoTW2IIjU/APuZGPYt9WVWGf1GMVGvQ4fxN8/N51eQp7fvEXKwStEXfYrDFNMiGa1OR
9vz5kUEcaZmsKXm9bPMYER23Biu8MZZCkkOReZG2A7j509bqzYN/O/KV7/xK5nljXS3IfmmohxAP
6FX2R15svF0GhTdQ92UB5VJRjDBl/ZAzRVhpISmmgYTVBXTpK2mGQqUy1KvPYGjMvVsgVRmPqfrK
URUJk8w1FCiryA8Wj2Jr7fFoi8QqTLCHwf6PRQA0HjK9cBOHb1dX584uzRMjawR1W24VDWTy1ZoY
Qu+vDZfGnd7UkXASKXRneThqpt876knqQ4/bZ6lM9sJ5CbV9wRFH67h796A6warDw+HbqRAGzBxk
kqbUnkEMYnVRS2wqWnWMltYnIT+/NxgQDOS04+BjuA5rdwHu044Ls9nWqbiBqvkNWPZu209sR+mW
NhOQlEo5OL3Odvh5G/DEHRybK/u1haJNnCK0F/KXCQCofuR7Wp8zKRy6pAgm9KDY2I4F2WnVK5XH
T1oVpeMlsSHzwH1AdBhsQMNfGG8i9He15Rr+dH8qjdO3v+5qeNo7WUSCZW+iq0w2KBODr8TgCjcM
pTj6sae9BhfBwmQN/KJ3VXHuWP9kMdIpO2IssRfaPdGc6R1eVYLSBMaZCDCeOCKFFrLLthMhY+2q
xz8yAY8CgnehHU0AnsOGgadYGpoPAWUUgVTgHMR01aIEOlKHEWmRwMtBxKeIYozLkl8mm5dBjfMz
4oL5XBbdDNBGn/47uMffKhU1ZinZlKO14aQ4mXcsWFR+nZYyiRfmtrWJFWWgkJ3Y374RmVTz3tfe
LjWK2ZIDhp9gujXnhkplmtr/kbYOCSvN2n1eAfuuEDb5cZZiuxtf2rZfpOGpoYGen2q2X6sKiDCz
GZZ8NtBBr/EYYLPn3h+Od4cnMlRqcdn9XnqLrYXKFJg/NLMaImpbxW8fbEWKZqtQbbJg0NUjl/8V
WFYbPTJfW2gh5slnMY2NCYLJRnEaGsQBkWmjcSmhezyzJIA3liQUNccB2spHL5jgrbQwlqMRIEJI
MyQEfJDhDXidQFk9BgHDKAg77Q6QUE+equSjKNY+1atA+DB29hhG6JSPU1oA106tblFj91PhpOIL
ea5kCOU7FogJaPJS4vtlhpwATMBDqmc+OUnSIODeGkjMXRwB0d67zkTsBF8iGZU9s7CJJQv2nrlt
QdX4EQJwkDpBfenLf1XTVkTsa+1e+Bc2OWqrsvae2XMhgM86KhzNUnbbavNsBxETsdsgjtB4ae6o
J+UAjd7i37tiqNZOalZt3+K1GR7zKiVCs1/AIlVLo5Pr2Uh7pa1wCwga3PxXqX3pi5wEsAOutMyp
x/igwRnfJe1ow6VLVhMRl5lrEWd13p73e+fa1VEzCHL85c37Akd/vFqC23RYOFMlSffvaNDHYC5L
D+PBUQ/3fHYfXUuVH6VNwm6YxcUyN9MYWBh+IlM40i9Ip8VcCuGGrXfB/6dVJlAOxVMUdRFJlJch
8oaxxx0UiFg6GY+fqyYM6xIyx0P5RGUXW4I27DrawuVLYyyu5S2PoTYsq5dT0h/tW60skTCz6PgX
EM9frx/i67D1uyrvCQzPDDh/lQbETFm9cJ71ksd3gipt8u5knVIfUyrJUCovIhTT5YO7ZmaI0JoY
JbdPGXnvJ2Px8/tYHXf/XWFkYmpabJmXF3k1UVwH7cT3dw26m5UlW+qnA1BcFWPkcgk0xr8y/uNE
3imfrXenYQzLVr8yhUaooCSUKyDvilxovT9u70UvTMF8rG8nOH2NmZFPyuRwLLDsDjzfphTPCbJI
+ktzOyPVSydMlpFDagCpKlpov8OnqWooGesI2GubfNpYFlBzz9y78+HTRi/zXR53OnRCBTb8e5nr
IwIkWIRlbZg2joA+VYsetkqNsyTXdzlpMafiJfSqWlye8kqNo3YNirDtAUCYMRbzWwiKf8gNB4YF
NUi59hI+prCdYwfzWT7veZfRhdlHDKT1YnWwlCOiuquqL3hS5SFEadwNxOpaOuJt1rfJ/8QmQXae
tIv6tBTdG23rdokdcNag9Lunb6uiZB6YtRWa4ze9wMdREgF3kaliqHdt/O/4KqcmLk8ufoSvaUuA
DolnNG5Nd0Tg9v25XNNtZAXL+fKKZ8v24hpW5cErRyFHb3Lt/00KOhRAo4GSTcDKxlXxEtgn1UNe
X2rPXbe78k7Fzuf2oWmpCaPKW874rhmHe6WypLxtuzL3pXECJ5u71Ck3VZBQFfyP/7MdDft2hiH/
wuHh+UooA82/8b+2sIQjO5gEp2iC6v+nHVO2NJVXKhQPdOdEH05m1F5/qjTLBrJxqCAXfLzsM913
LJEi+qUXsS7jLfQU1TYiigpFG0bIIeZN7p1jCPRAe9qS5SegzIEzgpyT6ZhZWPDaTaaHVrA1FYRJ
LrdwFLCcVeryJORmQ0oHCn5Uw2jI29umwtJO5OTlxfqjZYhwsRaw62ivO7DKEa9R5r0+rvsHb+QK
M0Sq9/IZXIyjO+T8TaBeftgK5oPdpnB/vHu0cjtmVXQyWECj7Cb/w/9pmnh0KRoc1FX1XseSDEZG
EhsAbWnkK6rkUANU8c2h5YxqyKW0x7MpZeAOzLn6D9YGTzmXJU88u/a1QtfXIJDc5kWQqLnPf3aO
oelvcCBnhbBzPjxnidzZJf5Jh72lCkTbQVOgNlwR76kdzHd3eb99dtaI2bgR9ONuxVyjwnNGmrEZ
Wakg4YyzPVYTHBG5TjJr9J2hOWMlsYJ7ibNRVJZV67t43wdx0gRHNd1/eNWJtWj6rG6RWMHdmUGC
53fsIztulTpr6AltO/YAt/CScgT3zFe7+mI+RX8Pg4M2DXVTl67GiAzLwsi4MDZqmszvonA/wp1X
hyNsgU3bE5StH5i0j06gjZfGaGYmb26jQkV6d+HP483M+yCTiXkRLAlzO+w0W88sDds4Gd0j5DSY
Cyv4PcC/7vXXtFVllkkVOdVBlU9s84Ue+9Li6V6BfF/Qu6GCrpAhCMjl8LdxpFgjaTga/HCvyPCE
xCnkSmC1MAVmMKhY0uH+PqdhTLJvtxpQvFgH0Q4T1CqZ+BhlCqIU9vO+WLsAeHZysoD41mb1VGlk
nWS/f5NSi9d0Kf88Vv4UrLyh2bamFoFLI7UiSQ+Myt4TJoiSbOis16W5jcutXwTaDPH/yG4bsAL1
CS9JTtcTWJqXpS5L5E6eTQQGi+zdLxX6R1ZrcxSWMvwIl9DjdOsaXlwj7/z8DI/etdorepyDqZ0z
4o+tpwBCwsz7jUMjXckeIrQVjwk/VLBj0i1eeJlaCKn0VFean4ufs1yqOFt4gNF6C6fj5FUeSxko
Gj1Isfx9apEKwODE0TaT5yP2hQ9lea8SJg/3IUiOOrMMvVqo5gftFBuK/9iHZUnxFVrXSjzVz00Z
ETi8803ha0riDpomL5+asjA8LyGP1zBRGLglg4Cqq0oCA4NXOLYsvZ8DNRrAChaHjyeYqrSzPKVz
qdmmuYMvPxLDiA52WoSKJaBkFF10vz/PL2+hrZEvS4jnYyWSqgbfpdxZci1Xcr97qErgaLwA5hf3
5TdUPF0XpvWVdRkiuo6TJOMG2DJWnCW5ILX4mFD/KxYR0D1X7g7zzV0cNAVun8pwWYb4CxggG1jl
ZuHrvLyg94o3Gs4YmiqMi+tddXKknf8ceuqd5DaDMVXh+m+Rx/bC3ub6NYb+2OabLn0Lo94NuQyf
oe4NBGsU+SWNEa7DTjN53Q5tBLPielma7/ZLWRUujXofk8ffL11ZnUYas09pAbAcNY7m79gSsyTS
N40yzmvMaA4yayD5pYTqCwfFCg9aYXx7pGndZTLYOZZ9lb/jyw/yEXFqjK87RrvfktT4Rfo2mit4
qwyH/rA38Di0UbXYa73wfEapKUOBQUnbVPkXwgS2Ed2LpKZQSEmX5pkKpuiATMkjIi3jMHbSWQnR
bWS0cKuCr7oVF2Qq03skgpdCO6Vxqx8uDttb0u/IabXTD2+BVqEZ8yJsFIecOtLZy9o/TXVx56hd
EsXoWwqur0O2mlJ9uqTEud9x22u1PwltHRwPRBxGpxL7z4Sr1NF3rmdHhHzu1fyVvxOUR9ip11EL
qNKl+X6N7CgD3nYSRY89FBbGqjauDBGxYavvXULNQsYkZB/PczOYbhEl8J1NTgpDZfOwjO7Wqe7e
Nh/UjCm/3ZowIIzqMH5z7U0SSejZWtfdyiZUTiSu5oAXH3V/ZakWGlv6pLvIFtujnv+TJsBTCqR8
OZt0TkGsRLWq7eugsQ+8ssM+iu1L6buRAplAV7McW1fQAv7lMYhnBE4IvraA/48TGg8URp8Tzs1I
hyYuxb8gGrIlCb5cRh8kXHZycnyKOPDWBS0imG/YPakPccrZ+dbj7WsmBDiSsEpu0grAxa7MlvuG
eWXKSwcEP/bh2mdoEDaRXAPp98oggQ2QDj2N9bM9LD6530OzsCf/R+Kk4JzpR5D07EXU/SDemH7P
mAo6QM9O1npj6VUU+u0mihLd5V/o7YZHSpy08CWFiWJY8SG7OIy6Cc2hrswVkuINSPsY7395Bccv
ABX50R7amvsAawBcAFayVAEmLyNQ2+/5Hg5Cn8mGHu2a/Xr4EEMIO8qV3drIix7T+qVhwXVh+zHv
l9g0aM5MiFdyTEFdBCAHHBbMMP5HX4xXlFskOcYwGd6vGPt/dsxX3QaYy08KkkMmpSbJUAtZPpwA
sO3AwK1PM8/IrizxnA8elJH4JzYDbtA4hoWiPrRwsGf34KiqkUjqbo2u4DsHYDX6inPuuxxakJE5
Lm0F6oZyi/3YpCGA9vvpDY7g+A1Dy7MhX2d8F3XVrG3bAc0jzyf1CsAZtCAuOXhXgNKxT6RhXz1u
l+6T9nDhFWwLkbvQxeLZWDgQxa3wLRMH2O6rtTgHxaeX+uYn4liHGrZF3+CDLVh2/51LHXxu3VSX
nNdbWcQ8jFOzXyVYaoVZ/SxJuCLEBKKL4+8CAfg5COmRcI34P6oAwommuHthIzFPkXCAgZNSJV5/
gPuI7h7UGTVdH/ggASAKVOI8U/Fb40wOkZC+TRxB3pllH3zMXwqHvcbz18qPcsvMJ4WHNuWBdszw
fiU5ankJ8Afolqk0+WD0R7yOA6DP8Skl5B2taClQ8vzWXZUWbMy761FOBeCgGZ1IPvmRRi1W2fFU
MZviIKJSPXBXtZ5oI1XsVdGUI4gIcyqxrhCrYGQCEXxJ7yEZWq/UGAduIz5gthsfBhdA7WhhUAsO
L/4iBsUDsSPYI/W1OTq0gvWeo8nQL5FyFdKJK+x2Izi9uWi3ejS55+N52CRbj0bPKebl3Zt0d3RW
If0tu4x6Kv87is8RLuaarz0SkwHjtuXxSDKiPF4tPZPHi5lFqFwp61iNj6lpKfLTTzbnHjAKfVrC
Wk7vuEz2B8teilnfsK2yAORJFcPJDR01J/vSSsF3HWNgK+eKuQAmwafzEQkOv1CiaC+myHtKW1Hg
Y81XJSL+aQEecNO7VHL3RazSmKhqljzbAxdjj5Y359Bl9hJKpZ9nBRebCh74J+pikyXFN/BG98Ng
XlQiG9Umy6HRi7giE4R5ScndbdmgXS7Khds0+IyZsjOVOMIEDwTquPvfuwIACyWDgFOPEwO0QuEp
3vSIwhO8kbz9znBe9NpCgcQUfCimWAtiuFwfxIsqrMLOgxBBShvmoRJI0rLxjpMqUI6Ul9UBRRmy
PcQD9drObkRi73IdJ7jIKyw4WrWG29xnrBSg+2GyAgAAEPPrpJ1O4q5TTk8BIgQVEa/14aUSrHSg
rthsuM+oRkMIRl93LC0uRpmGaYB4IgO4iokkH/8LU+oZcnQDIxyKjrZ0YA84vW9MnAnfBHIJCI7B
nCHiU93UYFUCqezy4HaFWyTKjEJXq/FnCyb3W5Md0a9KmkaJ0N8lMMVEniGbMrSYg1Ewqd4bmTA7
NS+6fShNztQyJNtCTX2eoAdFHKTFrFl7ucUurPHCZtOnLXQGx9aC6XryXCxwLkkmU6ZakKTx4NNX
n2GZlDEqga+vWUbDF5aDjsavwfSyse7l3SSqL/zzj2kxGcGeonZsZrrzoA1qqn3O6cHnb6DEyT1n
J0mmdv1SVdnkCo2lK65LY5je0yoIXsHMVpUkIT0dC120OocSg0aByycIOIB9EXJ6J3i5l8WgeGHU
5xXSAUYwL1AabgCP5f/l+uaDrIeCz1mS8G1zoUEEW4wnb9LNM0j0uQuM9UW1z+TzKZzrKsUGfz0w
ix2KxZGEJfVM5cD+MNaVTZxPjI8gr6QGGabXrA6X5Rcx0uD2RxQUiiNqyOSewFFXhNmuPWO/reVh
vlzUUGCbh1E1Ege8GzXiP8O6ag5BSfazc4yTBdrZA32EylKV6vjWQfqXboE4qTj4AWTumuZIjsVq
95Z/vuHC6K8ZMJe29bw5tFpGDAXxxEyvW7Q4Bqv2H95nH8Sc8ZcJjwV+NNMx7SdUw1xfm5+gew87
7/38ckwXq44JbKMLsIHfS4jcIqPFJM/JQu1K67cA8E+7k48bTMo7sOL/Cf1/qMcmYiHiZKB/P5HC
XftSAAYcKZmBZZoNQdlSBr4yxwZlnGWk97Y3rtELoIGEJe1VtDVkSzApClF9fOxGYDrP9xFmKQyn
azTct1LLhHpl2NF5UvRLrg10dzjK3svNEnYfYaX9aOnl1prvb0z6+m28vPhq8xOCPkeixejgXidO
Uqq0d+EUh6BdoxcZwXmWMDgz9A/2yMjMOvh2tWZDiVSA/jOJYJ2BNwGMpOCj1icQ1BxYuePOlxIT
5ZeXOmRnCKoSayhymubWgqFBsTNIMYNl3F7KSXQQaoUFUPHp3kd1Dx0uK2g8ByfkSW++iXVSmA1x
FcEDqfLGQruHouXhYUuhmsZb4O4Ka8cYw86k2qnCPgf62f3Orzx2/5JN8MucLcwt2FDsD+MWuvgC
TSslNAxHOKMo1lZ8b+OFnliYwWUM/5pFSUov1qljq9ZNi0MrNY73Rg6Ui49gcVE9n6zG2qQMxD4O
GOXutHlfgxZzIge7OmhDV891RBwsG61NRcFLi057HzfAhahkuVxJm5gaburKshz1/khDz/rGCq8g
U0TxDfUkVjnNmGF+rVI2yCe3BItcfqn9ff8L5JDhyUQV61vqE0r8zSWYchc32GFBvaBSWRKCLNhN
Ze05oXNGKlgUohSjwKSC14mUTxTKs/KQNL8KgeMzZAiDpHl0rMxkxwnamNLje8cvWhRTpFeEIw/t
6zWRTSN9zbkpUQlktG+G6jEKwolCgRpaYpyvyma+IgpAa4U1pU9qoCPJtdZFfzBYM7iy38DFE6Hq
/x5JhPOuVD1+XGzEYA855IEGp74oAsRtPt21I+SSgqvKl6k2TvsOMLfn8MCXQQWvJvgr93GdQ8IO
jcHn6dFB8pCz8tZyWYKkjMknSljLP0K6zGKVOctKi7hW1f0137mCfuJJQDQIqaHb3kMkH2Gr038X
OuBDSDIAHdsumKaXebgjqBdSqK1OvuHQr8czMHa1XLGKTddH64S3ts13+MCfpt4Qq72XNrPoZmnn
yOiqWo9WfsPfQv1ZC59swTTQ9vW+UniljpYii+CDxVRDjSq4lC0W+gsqLyd08XtX7UnQ3JlrH1iN
90i4EmC7tza9IYhcV6SMVgKWi6iALmLop3MS57nmeqfYwaj68nSW0w+huTCeFW6CvcJRBtXFAfHX
3/sX2t3FqPaXv4/tSh/iwyWoP3F4WQSm7Bnc/ShQBft/OksfmtbbHlPNwjrGzoa2YMs/MCRY5OeS
FPdYRNQASdI1VOSG/oxDxzPeNO/p50pvigE4Jk9aQ+xGYjdSTMFeboXnXIqqsUFQMHXuoRg09WkS
JdMai0dxAq/eEwIu7rbEt5LGNfslYQCXv/JbauX/CIuLCOEV3965SDNXMUeiZ4K/8SJlb0K0PREa
EBKhmA5t/vm7xk1wtKMejTQyZxGsyC8r6tH/SFrC2g/J8k+yCDToeVPRs2dIesAlNkfq02aF0cc9
Se00Ihd6fu0HJgBCGHPWnvoX/AnP3dJGf5HoOiQvBagUNDpS4ooajIDUHrUvY8mz9xUCLnvdu20b
SZWj5kU5wVfrahVage0iC7/UPCgL0CCsxcmkLenYXQCQDXtuVyTr4nPOCHTCPZK1EsgnBLX3WneP
BrE/dpacGO2EjS7J5JkEBOwLM4J0LLicvkOCwOM5FnneFXgKNuKo16gy21934IoJPq2OXixF9zcv
PPj2hb+kWJkejWVoGKM9MoycxCYJjfki9g8r7W9mIRgo8GpMQRQ8HQBQm5275YKmMIiEEiZsrCLm
F3CcIPeT41EYcDGg+2jIjUfHKE++NfygPyiA/l5AzA6ZdlD00wRkRsRwQreweBkP0pLvuMPIzvcH
X4X9YXVHohZj3aC87gBPGxhYTK1acSxKcxDOrS+pLR8maRKghR0IXkzOlIFP5WOzWNo9tHHeSfNW
W1P0NfFRNqa/WWi60uQVFGlHvSObPfaYb5kDeBFS57Hp+Mi6IFpB4qQr2h2LhOnqa9YfSKlk4Jif
A3gD8TahDfregZ0Y0lK8tAtC5g7NHfpWgnC5D6GE7zthIuULTLXUNefHj4+6Hdotb1GSCSoIvVRi
y1uOgZzXnR0vUhgLq2FrCKya9YPr+LKK7yc4eZA59GRNt/N8DPA2ILX6WS86HxiJKIynNiJKKTpb
B6ueUqKzgHfTeZI0Wh6cD01QimZMtC77Jup3mgcVNPIN16Y70qXWhLSJzw9Lk3kqIwZYDXGZiUD3
9R3CAaBGXWmA+9WQtam5o7UhCamjJlQ8DgqZFyYPAEADxUiunqhU6UJ1nyemodi9nfw6TEzsIkCK
WSCaj+6vZm7yCbzcX/hjRx9wyxe4hWLnT3ngEP5oe90vwHheXEJ3Z4AuM+QIQ7HyFF3xUsmusNk1
BYCTdfdR0hoHXeWwZxlin80GErFVaOpHQZmoL4DhpQ7sBJR7tvwttEfF06lRAf9xb7QmpDuJPFz5
z+enLtAIb7Z5JBwGJbDhRdfvFlzVqgeqJekkeDQUbnzFtyzCjma4CM2lKUJiJf5Dr8DuXEDU+rPS
Fw9Jz+QLu4UAq2kGon7b80tcgKVWnWOzKuoAB5Q1z2utyN2kLRC3HK+8Nzg0VEVXWM0Zv9bRGwaM
3EweEof/ZAi5EVZjlS/FczHiRaWbvNMwDNx8vwOBduKGGzmd9F5IkxspXDf4n9WaCZuvd4+AkRgE
ef7h5Gft/KbuRkBfheE5f/bnOz6fQnnNwJakdTu1pmKfuQFagA2dT9hz81VEySN4WcnhErHsNw4X
AiCh7IlCP30qK8moApNtZT4QfzAgsRaXXllXf4FJ9Ox4lFF7uC1zSFfno7vHHGQKYxpzrY03lku6
4bFkzqNiif2dVoItWFsZZXUV9/vhKFCafFWkRfuse8kHcwnbNv69aavB0nyTmlcU7qBb6X/YPu3X
3E/9NZ1DHfNJLTubE/jTiKa6ILneLejUYJwY3l+TXKrHV1i3Sv7Uit1kH4CmxAxv4aRaiCLTbZf9
6F+WjuZ+2/dXG7yCoMQjBPqe/0jc3y9UkBbtj+cW+hRKcdbN8RwJYcH0RSUD6U4aowNKNC/ovsoV
4XSKfmyuakee1tlBRZnVdc8wRTD0isymRFv0S/XT3cSa2fPc9jcWQ69RWs/7hj6D1mvM7L85Xux1
rlMANeTnf3+REtJfji15GAxo2AnqRgkTSbY0qvOCyVxzqDZk6IF+IpwcyTOSU4e+xW1dtPqK2N4w
nbOLeAhdGwYlw9I+zn/HsgfOERcpsZIogcB8DJNH5BYcByFHi7t2mA6KFhbU4Ue6tu9KI7aSye2P
m2o3s0NQvjQd8Hm9zdcdoZ+gzpReQzGGawx2tAndax9JN2ShJItQKGXcpMi/02JDSb905RR+Vv2F
ty4WX7AvMWJnZLBXgFVMFwS1GEvBPVetoN3MEPzuKOsDbnuZDSzbftjdEIPxDWHCH+DXZTAbmXBd
cXhNc2NptG2TYYc1fPNAtKu6pbfNgjf88UU+derURRryojmgv/8gq/PwaXejbYDB2z93WrLl/ZCR
gsnghUGJLB3+WnSBczln4nNegyQegRL7wBh4MJBUlup2aYYxqCHkVtfp/2O6ztHp2R3vG83x0QrB
eM2WxUZOHIRM1HZMR4NWk9/Hu40+bOSbGKdE7n4xMZRnqv5U2mVa38nAfVv4AX4bn7FVAE/1Be8t
XIivEwjFO7qCM6RW2PPy9Bu0wtmmzUegb2BkHWsALE2PED3Dl6dQkfWQ+Q5S8jfSvwa1Y5zC+L5W
AHSdlyK3HPM29hS/dl3e+bqrzO48/e1qIR0nExz2lpi4Av5HMyqhMx2WtSIawlThZiNJCMLQV3mH
8AJfca2qFiexd3+9GR0NMsHcSbp918s3O9LjkCdJbHrFpOVbCOYkzKBNIwt/hSqm0XE40wJHivCM
Tvh0AXdxT+yUeQb9QozsrnAdELSKNmLxvOwb6bMbvJn9cIwKtBfK+Ol+W5ZgwD+ZhGNlquZ30Yf9
RCkDP9xD4yNkA1WEgmL78OhktnIQBK6hYvgtJip30ceNnrJh+inilD0bQqkatibfST10RY7/Of6H
wVzPM7du8hicnXVqc+RaUiBOmyLAXn99ynBK1uSr9FW80zPbC6kHHY6fuvTvX9AS3xPmDjDjSzd+
TmGI8dtVAClZ5qxbt8hLPAnOvjZAjOBtZ6W+84S5nsS44Riz0Puu7g0CBWvYPy0+gNsrkUkY9cz9
Amd4QfJyS5QaujiHO/3Q/bP+gI2K6xPQLEKE4/K8uOQbHeYtPqyD709nhrfF82XloZvIznaX3INs
Ie2U7kBpe336wZudA066pEt1xIlevcLLO1p13maZHI7MxIPYFrbTCaJuTdo+5ahSIcqFaHT4s60j
8jorgBqLbKOJpTdVcYPgDzuPaYeuFqjiQmodQM02JxbWcnOX6/CYqeHv/OgWvEeTmWQP2+dRbhFX
uuevMoOazyLFQx2gJdrIiDwQAENiHGXt1Ws/+HHCXXvbwRDols8MgRy2AMboilvWYLxiQwKOf11K
8jkpyanxq6LNQuEWNuoEyCVSuDsWfnJef3iGDKpBTMDXyiwzVFZF6BzPsE4tAa4CHyLf3cF5D/kk
i8GFKYgCU+8ntFYiIYoRkAKNq95QOSk9xClx68L5RZ6vw/1NMBC08dMgiZmPqlpuiCipAIdh6jkG
IrtUT2qFJpKX+wfFPcMna52rxWC0Dk04ufkOH6u2ZzEedUODnPLAnqOrMB5cEYKo8PV6eBSbUrAS
4LZVmFOGuuuiujpRj3ENnaxXYHJEoaZWsAOKfujcyYyVHEWPOsLpLDLT9rYv0iuA6MNJ6t5smqaf
6mqTiyK+ZRjdIipZU1iFfm+AuYD3T4P70bWJBidU0hudNmI/QkbtFFftdOzvIyuKhIv7CxXa4Mk2
ESeiOPFqVxddzBJOFnz5vHkfxx2wdywS3JFSXWZP6MLTwaCQLmc7ejkQ+rHlkiDdMRFAewDz/8k/
BVkfEgiP3kebTuma2OpSFwbbcAAoEl7ItgHh04QNngHcsc9tvA8cQeVUnr7umfRuF8KojnWzJfac
YABmx0Q65nWuoHGQ8u0b09aNvTlsL4QtNmZaMr1I8Jr7EjtvaNK+/3XUNqmBAZJab78q8xvvp/Em
6AardjmYYPQ6huigCeUKBKBvsNseIMuE5rsxDb6hZVShdDYlO45wME1acsk30wnQgc6faDjdSLS0
p0IK+nEJWiGd//sZ5m+XubQfLpFAo5KXo5PpU/sEikWf7odL1UJqW3MmSoWMX7KusKznt/+neh4d
zYDOPpKiEod443T2vrOLClPs1S3y6lsgk8ojckJnrr7a2BEA+KEA0VmIOrKgaumzODEN4ht+x4pZ
T5FvBROTbMNPMpaLNyHKIsJYrl2Zc3OuXQi13mZaKc5cnLG+62gCtwiOUe6dN+Zkqw2ndbstQ9/9
aN+k9kcUhqVcueHp52pYxdI4u5b54/kMdxe2gfc35WeQ63NTlaytpOu3x4mz0MV98BBAGufmYO6T
g5NUrT03BEMjH7C30JXtTUAiCKy7pI4qgFmSFWXIPYbmtXpP2cIUQ+5W0DmzNYIERJntZoqFXULp
5uyVO/S9C5xG8+CEx2rzBgg8Qo9oL1JRUswI+zY0YV+WeVIGRMGLuIypB6vW+214pvXHJxHuBb3X
V3aUrIXG+Ej6iHA0vuuR7wB3cKgxiNU3McB8nXswO6a10KbbnOWwmpzIlS7h8rCmikEnRo/dAWIv
K2y874J+sRqxPjOQHrGwysLKHGFvaAZ+uD7qAXBuwFe02LMx5SscsYjBPui2Gr4ICRc2v9qk/oY8
ZKVNK720G0n2YgYlr5HmkmcgzLPEqe0BNEOcmmHjTbx1RpB7nHHleWgxu+W6GUIu4WM75UWfl0WC
sBer6XqhaS8HU5NGC+OYxCs6E43Yyjn7Dd6bB/8b68I3dw5/MNHrDeKOJazxrtTuaxagvy/xjsDF
P1EdPzoGPk6mk/IRAIZqVs8aWoSkdfaJgu7eNM4P85C1jlcODqqX8floisdFNkHJJaTcqYFIRR9C
6nWpuFx9YDY98AX8PuRPvFYBPlj3Aks0CLpmyr6RuI8jEUjcdouU0raNbTWh850vqWp4+xhrFt2r
QnY4eZcOHPH13Plg4jHoF5pp4IvelI8Nh1mH1NX7cFWJr+LQLumvBw4g3avhQX12R6UHzmW5pVzh
NRvKPN/5mU/Y3vIs+vz/5r3kZsWsqgnejDWEbRCR9x5nHDd7gp2kPOVzxc5EVTBMdC1xTaPG/q12
wzPgGYgfCuBQ92pJKN/VCurES7yG+Fs+YkxgwWS872qu5krsVA5yyyOgOOmder1Byxz+P4CXKhPz
A2Nj201DLsWm3Kv1Smub7fSmx3dFe7uNcbwbwK/ldQCFFo3tTUfTORy3grbGu9KgTwI1zdZ0y2Jc
yzWnO0RrvLEG2XbHnXfQYlfgjxdKDGUTSP3hMHXu9xs++BeufJa5G6/gKQLNRme3Fe9e580nNBjq
1sdEhWic1QnXAEE8A7OUKO5n1CPgM+UDRZHM6P3V3Qn0SWy2INyRowIe6we1kPipr5vm/H+/b6Hu
LHH3wYNQAH0jzUc3Ao9dSDXtSWgFijoxYs41Rtem2E94Ik2XIVDQb9e2TaOblZRocKvnNCQzlJsf
X0lfQ55X4tln0U31wYRdMxH4QlYooCFzE6Kv6CjQutWXf8t44LUbYR2Z1ai4iZfIw+iK55xKl5cF
vLSHkZ/BAPB4gOMUJtANAm5wXcSK/WlkLTr9kficSFEgjxJW88wLG3ZEz4PcH32FvFueoePnyDZt
9u+orsDcyVEYXmy22Mdbkuayl5TcvKNK/v+RDnEWL6Aov21RUmhid+9RqXDEc8CCEVIZ51O6T8Qr
9egrar77idPb5U+hGvWYLQ3MiJNvLvEpKW3NtSlcTqqaOGgSwc6EI1FDtszUM7/txNgBk+EEEwqY
NCuVcol32V/qwF+6philpRsYPtqFyHsJnZVTp552yTfOOH0Po5Tyl5jzD5jA7zAjk7CBGMDHSXDJ
HqGAuMrRiN2vn49mMkgHAtvW2ZusYufdoicpgmNcArwQD3F6MIKHKyNdzJfFTdHrbHviSXpW+pYC
5CQDS68RPR+VjWpndxTI5ffSBGgm2TkrEzBiQNmh8YrxT5m7vysKHIZoxxQjGaju7ZAI2svph1tc
lUFYKSKPFJWi/g8Sv+Cy2T8TwjmXDY+qnxIGegnPleAPRURQk3dtSvy/F4jq2y87e2NWPHxkEfPC
dMjSvTIVlfLcQbjDzxDYNhJKmYz9HkWLiBwgzfGvscqnOsyRgGE3lEsRWbaxliTSPkbAZNIaPHxE
q3nY1SRfyNakpcm06Es8tDqs178ydZ234cYHLsvr88e3UzkIssjFONJI2V9h3mdiIzqBALzDNjVp
GsFkISTE6IsK5Vjo5K3ZWJDuKEwLvzgowhO6T9YLFSvCvwxE9Fl0+H8vqX0CG4CeqGUyvjDdw1q+
4Cxun8exhyORDu3zLpU6NlxbYpIXCJ5Dh+emmrmO/jCV9zv7z7gQhGaC5G/u2SE5APIJjyqJLPlQ
fWK4RDh4Ig4RnLwX7r/qwb0WcnvTw8sEdrc1cbQuZQBGGBrUPwZBhERf3IdFOc15tVcwD1YG11iv
J0pVAnJLVJbVuoPdSYZS/jvSe8kahzf1mLdfppPxFQtxxaUB8U7OjYt2vcCzAXzHevuZLIC7OV0K
9v7mq9MlkNVJW2m2J2Sz40vN+TbOq9AGuaYX1HEjAqZD7FtZEzdxsmogMAFxJCm5MbbERrW8Lcix
Op2XMZY4YPKvnd81BYH7MhTO3R5ssUJTmeztQ+T4v1MWA83DMCCfuLxrhRrjLYCSygFrXWcHuPGD
IKHAv6rSi9SfPRrZu+qjXjMN4o8QODGelnLl558PUgFUz6OHjg7eUEUL+lQHVYJefgsFXzpmgcJh
mPWY1B7xTjoy1+T1L9rYIuYTCEwwytnPkRWd60UV1rD4I39lNZnZdHywQEQnhe9JXmTsSuE/5u+U
6OpFn2Aleqwdas6cObqTxDf5lDPFgcT0kmiZQMofc0IGjX9Yd1RVlnukMO5Wmt9ErrA3WDnfMzpg
LCY8XjJzyWxQOf/qGAhsSXcgUeQZsVp/pn5IL0uEorZ2uQkJtYAqf7IXQ2h7HNnKS81u2bwc/v1F
WEhkHxkoWaZi/EmAKEnWI0dO171RbzuLRXQZPvj7lZMCkL41m0efTo3wabY33yRPDydBVrhgGDne
vHIThNG/yrB5LyQK2z7QXTLKyUh4s35apaNZ+bjZ8Rm8gpgTrJtv422MDuNX9tI5NDZmkHRq8Hin
kitM/FPkYv+0bqX6fDFM/IGOu0VFPoFySb0CFsbm90Od0Kzv6a6onqo8DnsQz7vfdkG6LKhiAvzG
aUDMRd19Dl9sEtj5hWFdHL9xrPJ/aG1RM1dJ9cyEyoDtPMlI2CsG7UwPKTPSPKBL8QeiTbLo09Ad
nRUFNEPzbwk3d8aZPul14BrO1RHA0TqW/Msg7FmAq0tGrQOt3MlgIOVMkCrj+MYzacRTRw0KTJ0w
UIfLmXEos1eizFITGlF3tzMQx2CfpgXAvgNtet9hd1cx+ABDitph+kNayaFzJxX7p20LUaCF9mZl
vrXRWzjckvMJyAjsE6rZi344eJaQNc7G9KDgrfeZ7oh7/pixeYpYKxtqnPQPi2f1GwU3Fcn8X61A
DLKGOGn0l8NMvlaNl9G7ia+K5IkkyyMNPqENu28j8Z4IzhPwGgCIXlMTqC3aRR9DLr+l9/UKQpNL
vaI5fSSjIVjWOgqfDaPHtB7x1YUOXNqogh8wu0U2KT+y+y9YoR9siPg+LXb2GPiwb5Tqk9PhGybf
wsT5kfOccR7NqFkXEpXfNLIMCKEh7TmjVwiXx+KLsH53N25IDLEWfv3RvCezpcxaKq+CuqVuxrqj
hkvOJbrw3KAXudxgGk3Gqecq8Nj3PLHjUJal2x9RfODu7bv9okTIhFJi3U0NOFjc8NwwFDDt8cUs
hcclvMPN75PPS7VhrHUfhrK7+l6HOX1xUFbxjFOUyJAPyQActfii0W4QSobeccnNt86OkAzkHKOX
OxpN0pnfxoMEZfoA0E/OekTtzCr1YY+GMQnhlBorFgBViNHyXSxsaBKCgHwP8oW63+4D+C5dK7sm
053bVSE0GCTy72UPvP9tYf30cvad0CcSVqpqLV9BJ4qKfXD7w8BroY//NgzWYf97tjDH3PldLi1p
0K3+POSo3mHwlXb+m51O6SNkxLaBTVnCU7i3c3Kc93tIaltRv7iDIbrTW6qTaqbnIngrQeMA7TJO
AhjFKGfW7eeCuu5OyPmJ+xiXyXM6kXAVXGcOk6A/7Wk1ytYTnTnLGxNP52y8V4focAD7SQED1ePu
2mgcmYmzFKUIiukpCo9oHXA78bVhdukZzRtzC0A+4ILvohNsfvlZN683aw9rpbJGXuHWa2ln9+4r
DwwwNRV7doHz/C3HRsW1sAH8MRm5AhmCBLQEZUCE26MmDgGCSBpbLJBcqOd4plgilyuMrt1VJETx
5s82ytKpOwi7U73EC1Ygmt09qoCQ6Ym1nYIZMvWNI/xoyHv2u46Wys8pj1gLEAMfWjPG1lryLOUT
WWb6Ps/8gPtlN1WAaxwFm3S3MbqP8StUZJTWG07yIt8maC3LLkorlLY3cbL+VSFoI1DgTzc9Qcd6
8A7hoCZ8CpKlvz/yilZ3+FqSm3kze1gmcJij9Quop6Pv3LSVqQ1smWh3nsqfPtSpZ9o42AWhxuOO
k8nOe+XjzSrLrv97DVEmodpZf5EsNUGCgkgm0GiCCnmCcSZCh04T7/4u7hiofVhvXq0YSLDjGNtl
srMNrdiBfwq1VoIjdCizqRiHdVhulcy3uNK7sRL8REjItXyu41RCo6sP6ok3GnOeFMwG3jUbWE2A
isRMKBmE5uL0xenBJIOV6EU6oT4YQr8HoIZ5JjXAh6Ks4mZSGm59jB0AFfYxI/MYksmMXmjArQTX
1pzDNDvQ9c0Kcw6Pd80z24VDzX8le6HkveSIKUcZQrPXcV6WJHclfiN6Pk8dWbpQh7x+/B2m2b3B
02tlRa9dBLc0f181c1c4oH1nhzyxZ6iUCIVxOYaXQMjSwYaVFdkhQbEe5CJkY1I+FPEX2W9LV4wN
z+ki7sjwefVOQ6+LheA7R7Vcj2xdg3tQ4/GnB5fHqa2A+tYLdJ++KkN4TobFwhAoBIz2ODENQeLM
2S4i4SRAkfCofDhPN1kClKQfHBdDLt6oo/F/a90RiaTq6aRue54Hcb82bVRvDRDQZ6RCLMbmPZY+
WZdFNgMaGbustuwfDoxZVfh1RiB8QBTTWKtQTiX2h0qRpzNekt9Og/7QDFqb0iEx0TC8okdrE6kI
UcRb+/qDt7zG2cTRaFFSito9j3i/j/X634bWnf6kDPH0Lbq1TPcpMFAKV5QRqtZ+MWMzISEQeKnt
10If6NYjUp0d+mgmOb+U7x7AKNPwc3e/LU7bsINH5/wGPTuc9kRFBXEwy8FY+dDZM6wH7ePE2R5m
+yQCrBY6R2zOu2q4fL0JqPsdngymVdpNNAfkWsDBjlJEnQ+HMirg7fhjIrmuQqvtISrv2kZ8AMMO
bKspnfIcB/2/PbiNOzrO2KOyyapeodxg4kzq2eSDE3ifOJpHnntla8xrLDIZBMk9rDhgvzZOg2YI
dODdnBkgOXdqcC6JjgS/fSe+hCNE90ByCcvKHjyFbbHwGsG5YKOWk+U/nyVvNa9BiqzUv/OnpOHY
PZg/iiCV6csEw3GYDGpz+e+mtHJiysgZpgAvJ2MaoB4A41rb4wuBeysqyXdCsOjOMGXMHZ0nSNJL
onKB/EbI8bTn8++hGrKmmIa1Wqj7VhWdW4V1FVJF7muqE91O+zImZA6aoTphX6XzYENAxLnxgAxi
17PA7n6I39VmCPI7DPy3d1huOxOv36H0k3TLo3WdCqFFA/I5cC/z/lMepdbhleXdLJEOmaRNAKa0
JocQcl3TXCxLeV3f2Uw9FoMhgQYqS48tNq3yJRjzGEHNHQEelqul9i27ogXDi5VJKnbqQFa7fNeE
U5kbvVEhEKvef+ZUaCzKMrPp1FR3wbykoAlruIQwR8E4yF1XZuWjHN1p6EiEdnxvaeoa3mtEnFna
Yuz+lUHZLNYXZ+68jOsCQzU68K5lfk9CMq7ckUvZkyLodg2c5xAw91XQ7MS1UEaXHf/o3ffUawW4
ABoYyZaoRETj747NzCtpM5YAb4yn4M1OoeauhnTGq2QJWBLYLTzsSZlYN+g70KbVuX6dP7X0jjMa
PR5xmTnvP8ck9c98HzAMnd3uQS/ptONO3fA1EWfcG+EqUULcY2seZDCqQNOfQksCLXvHHxQ/6QRY
31LH3GyNHLjT9yUsAPolJ/DAU4rk5DtVlz3Iy6q8lfVpLesFc6uwjAOxi1d3hvrhyqyp/mdxuNs7
YUK+14TDSMktYSmLq3TngS/O9Q5V57X/PYc6P8Lb4AnIl4PTNz0tGXjV0yk5ALWi7TGMa9oEDcX1
X8lO53kmdxjt7fjuongQYA8eMdHVLgLjR97bOoDTT9xkphLmJalHiwNrzL4vBQtoWQcqm4hheIlz
LqORdItAakmEYfsXwluKtLJqc6fIO1Dgr4a2NMn5EDoeT2YZfIv6rKD1O4z7dyj1FPuUDcCjFlj4
BM6KR8NEVGwYpeO3+CNUT3NU9lM11ixe1TD7C8f3TDxf+Ow0PHJ4TLktPqf/WOsI8HNyz0zUe+4b
CliU0oGNAQyz+ziIcdPv/Xazjk8/u3Zqs12klopExVQKZb+I/bBJNz2AbcXuuQnSPH+h3y0cHrHz
p7vmMoN/ugpfE8AeajEb1e3sYsB/QR0DCDJ9H/Azhmj668FpugCczwZeKzDqfVZ2b+3YTGzlA3Ce
4hgiFyV2P1ZiY/Ri3SRcERVnaQwtzRrrUWITExMvU/3lufUXJXqn2TR0hcpY1FJbB3PvEfCwD0jK
FwBhrTmmJJK2+x7HvtByI8b8hUy7Q7au+5HoEnch7ZxaFxsk+rH+OGR9c5REP3+irhyr71jfM/GD
x95/IH8OaHVyevnc5ytsXfI3mper8hLHk5JlhqKLvHrvMeM17FUDUvFuwZnIyxKiu+1fWA/Bbif2
q+FrawAciJk3I+vRfTmpNhZ4XyavKi76UJQqXI6YMVLeZd9IXqNbxiiSyV284H0FtLFhrgqVS0Zn
xjYKl5+DFMYhwE55EkHwLznAE/+0HfUf4W67d85MWdlmjIJx2O3FNvObRlQazyWhPtF8nqJYPWtX
V2mP0de02bFCq0UuaJd4hEVL1IESFHcl0VDrGtmpVphwqiRwwQOf14MbSd342ByFlN/T1OOo6Plv
4078JR3IAZnqyuNh77adEPMlwphqzeCJdp0Lx0/nd8f9f7nXezXxLdhCVTkG7ynNnGPsxiacoxx4
UiAVRkENggsUD3/ct2HbmqNf4dwOt9L6+Dko4NZpm6a4lH8ByIoPRVvtmB3zWRLfbxNanxN2qa1U
eBmwtTnAfCiF1+wX0Kwcrh4ZhXSmlancJRt+05ZD6Jq4Cdu9+2ujxk4x7yIaOvBQrq2NR+PlXObj
qstDn+IdCtDPyra9peIudB5gF9efr+TmYTk5R4ZWxEb6CCTmrGZweJ9VPsEKYAXB/GU48u+O6oL+
4O8DH8QfZ1GrBGSb0B1GY6PbrEnfdh0WHAMqbKBTLG8xAgnyUgre/sKW0gXC0iA4ZQ19vi8FJaeo
q5PgDM44YcUP6H/4uJZLuallSdDZzkfztdRlTOGvZqn7tLfNB1xugFGl1PlU69Izz2pXTXtJzyFi
SKWtoKy96mr3ZQLO3ibBSIZvT/8V2lx/K1B7adss8eLQLUMfPQAHl4QnvfvX/JR9182hz1cdpjkD
94OzCAINjUAUhDqKugLiTYM9p/rWREbw2SADgaK6TVbjttMee9qYMCw8AjDeFKPUcqQYXNbSpwh7
9UuCq/5m1IIfnntQk+RGjEri9/yRDB0hWGI7D9Vb29FsoQD5T1w/N3qRuH+WAx8gPT/ucYNgsrbK
FloGIdPN9IpIdOQKM29iBqOQLkDFOBmJiYQnPWkS6pjr571+rDWBuaZ3MiB0oXb+UuKnDTI+G6t2
TzYNG5N8QBE+zEkNgNk+huLdxsZX1HWYLFiOjCCWfwqcL6N+D01WGa03hLSqW+OF4S1tt83tqUWC
4UmCV3takcFo8mFQeFlq1Y/JM1nGBy3HXO/3xHAWbL6jClB6OlAJf2/cogKLp/mci35Th1T+zd5y
rHGguakpvv7tvOV/3pmuJIjKufEPXTxTsZd0hGXtnDOa3OP0jOTyvq3NjI2ljzw+5OfsbmFyT3pI
3Ji/3y5vOTlMdmNfQ6dOdsuEnGxilhCNfqGNn4T2tO71zVXhQ2ZfoboWDvIvvYlmqtqf+QwXe0l+
7RsY2NW5/10AKzoMXCai2jTo1IfGfbBp6Dp/3geaa2UWdCyA73cIxRLHyfaNQG8M6vRU7QUYOz1M
60KtcQtj79DIBM3OBXbxO2DA8bTOqWmTEM2HSb6DaNcTJSDjBAmsT+V25A+5pjJH3eD4FUNHmPPc
L8A6QAA+tN4N2a0Lzab43zo8bRI7QBKlLFqF+SONkRKtNy1vZrtXKbA4DwtXnsuC3N+E3ezYsy+y
4X6NiMWIDHAB7u+Uk0uRxhmIOu2HXS7ta8EGT73KSSR51eOjtVc2AkDy7lvuUWn706t3fKpNQVOF
Xu14e3BhdkkOPxgM2uksaA6bgYhCoMaQEYF8h9dWJdmjDA31b/fG4bAKlTGV/SvqK0U/omlSIsfm
aEhM+pCh8e1PsaSKSkoohe3tP1jruYAR7cfN0Vo0aSckXyKlQa6QT7hJCG8zLGQ4Fnm7DcnxggEn
GL7Lx1BddueP27BzNx0wvTG3XzDEEYnBBGdC8fYgV+r3+vJQFr/w9ME7DkmwJT5bnrio/QipvP0B
LuD0z4m63JPiJ3GLpkmH+4k8VcI2/DjduTJ5D64KnilFSVUgFe7O2AOvnAsNu9Yl7+PZhddL7Oej
ykeM1SYNjN20W0hxwE3AgwjMvWqSSwuIgkkTDWeH2wH6+cw9DZvR5mmqrIzwdqlzpRVsUPqJu4XM
lVmWJFw6D0h4ROxWSmNE7ctrpycrG9ujBVBg1wvg1RssICc9KA5Kq3PaSuhSvVJw24tv1vF6sJc2
5PgQI3azzpmpK5Niph6kyUGdU9tTvL7ft78rja1guORq0+78WLfKmha/x3EjyKn+VSIV/EQswgln
nfIwPXfo6Sm3/18WiToJTi+EMeXaTr3A5m77s/Hs6t1CjziaPFGwQ5HJoJsloHMQz//NE9W85Mtl
YiCA1a7HqWFIPymdjPd1Eq+aoXU6k2hZRkzNm0aMFtX9Znq0e07nTmeLL3u4H/qI9wpHLG30YjDq
420u7pf7i4r9497x6yCr3I86WOKNarGV4Oc5pbfTANmk/UyPss+pGF0U20aeHF65YTIbwFikMQy/
Jq4MywlyTpB2im08hecsN/chJemjd8SFuzMKU/ivP516AOYRMuuh5Ix+xbbxzSjabBescn9OMn/0
lTW9JQsIJv6guBuBoztreaQEPI3DGkQAOrK4qrEgoTFTQODYysEjDi2PIseMPOqvXbjJ0nSt30L1
BekXt0Dh5AxT8X4nW/3T+Y7li4O8n3VKiMeeufOIV5C8GLAIE+8ie4qDepfYE9cMdGjAdOBhcZtX
+XE6c7C17TJrlCb1DpGEpVUUjrIKYl0V+E2mrTB4OqpCcC+d8c+kUOZk/LOHzHS8ZUPWEJJZG89w
h4fzgn373STpcWZf43VPxkVK0DW3uN17nDChKW7noe6VYhGcIwgTKpuqiF7JtkecDsUNyz3yqcf4
sQUMZRTtfGb9VGt/FLIdS4DFhuqUwC7d7H/iMFcK5CktVMGFuwo+KmXfwYDxvzC7+R1yAaWrhBMV
+YTQkB+AWY6ni49xAbdpVsDgdfMS1K1hjei5JIvkuXaAPWYMIrciiL7De4xOO2Nq4udDl7InKKkV
uOWOJ8Ga9DQ8kILUjbC/51Da+1/pX5Rlq8md6bCIpzBLTnOqL4T9rvr/bhQKxzsLOyLGwU5FsYj0
95gHX+o1pIGfa+umTceZcMsxA/LIidZe99535m1oCgsrTCOzXBu1QBLSCxuiJaLhU4T483asR7Sa
48sqMRWNfTMAA6drrd85tl7Iwuw7K/QTx5/Lept4JFseiOKxJa7NuyMRbVDXFfnP8TLrvJKaC4SA
C8GAVHfDR4yu0JWMLyuDaSU0vah3gmy08DYS0wWHMeAC42gC/SOTkFhlLZ2bDH9Xahv1to2li+am
A3A3ie4T7UeBML0w05QSKx0rZl9flNBgJdpux+YHXp7wvc0A4DKmAHNxpYTxZBo/7/YJEtxMjLbS
WAibbvTSovqUsIN/KRNPtLEgmVROQvVIjfE9hcNmeGTqzzjWRG+vtZoTba4lHji40GYjzI5HZvc0
vzWg4taRteim7L9j4MZqPwF7LoDs2fKJycnS0cSazlvj8GiYgV+sXx7mQImC5NxHcChGcZlDx/Qz
YkTngu8FqQTqdTz4jOo3YdzaD8HlFbKlYLI6lpMcQFxynWmiJUpGYU/vCEZK3Bt1uhCSwe/Gszlm
w+uNEKGdcJdOL+ngIbiayaSmbv8z6nG4u8krg4ndJOuwIpZEo882TsH9S+D/+hYTxMnh2pUQORY4
rDQmjzWuBVPH6SqYko6VTueUixBoap4zl3WWr53Yae85VO+ibfKAlsBPLn2JOjxpZ7E2GU/CIoB5
GFpw4srW8AcpUMbR1Vy6VAad1SrDPpZ2Ik4USLC+bKNmcxoOIi6rgAGI52mXjH7clNXb55a5ukWI
TKLSlnoQnvQVVEV9gUkahci7r3WVzlvd8TMSkTlqn2G/lnj5rWpNsM8cpBYpVsciCw7tHtkt9SrM
/cEXrbzP3wbGaDPcWpB7wAVK7OtaVI563OqOHMOMTq5fUfgt8vmUNmrd6f+t3c42d64yf3jhLRpX
JyL8xTyJaHp1Y1rXnhCr1grmIYHaKBBNNcTvVH2vORmL7tJjp7BypUW5L2Peipi5lpk13pyjjvtx
JPfXI6m4SW7sOpg2jWLyuRRlXNmoyifXYXGNnriCSp4VNPwM/6Ae4jG7M3aaid3wLKa4C5ODuZYs
ryMMqtORMHIZITLFoX8now4ys2xmKUhQeq3miTmw1Z5CdcfUZMf9WdBdf5KVa6YzjXw2AIqmd4L9
PkO1+jInQxTXKy4x/Piwp97QFW8iMwWkOHfSqCbSuAqlxx4HXRdNhFm1+EwQibbUW1+IVTeYDauL
+hvs0LuyQMnN/DipbmcE8BE7NYSbCF85DPybtIjzEFWEaddVrL9UmzAiyRbGoSJTFj+cCua5qm05
pqh/KEkRfZqdAGhfjowl72A+CiRIP30Wggw5ZzC9yjf/Ct5nHeY/agV7IxxaxgxECpFxmltDFq3J
N1KIjYpMh1E3LnsZOKtikoJjs5wiZoEVVH3wzDdXVObyKYVSHkrUDuhNsMThqi8bSHxNJWmVOs36
ozgpDQj5XS9nzIAHdJcfUz1q2syGZm0xq6q91xRpERApXHH459eD+yrFJKLT5zhJPwXPBU+G/q8D
sqwwKII43YA4Es1tUUPF4A2bUJoPYCil1plt+6TDtYCOXGO+cFYFrIiWy6oQfelPfwuVWhB3gXQq
1epOCz1p7aQidtrPDLuvN++bYanAeUm/D8FwnP8oibQ/FfWb3ccTuRilg42ZSOZbe90OCD2f3Vgn
A+SkgmU8fPxl756nLJakUDgnHWTEq9owpozt8ClCHm/YhbgdRj14deDVmzvtp2ecSiaLoltpEi9I
m44xH5e8n3tO1PrpxCV18BAy2DNFTk+AX3Jmc30N/xY3fSTodYUjVDBOf5fDd1dVXrRg4sc1VNbn
I9bYG1nvKysJygOmNIYGFapGJjXsheTW2arfDdVyRp7objNC5Pbq+RZHuzGl/pBc556ZOFM92Q2T
1KdEt1w6zZ5vktAiJV/0IsbQjkRYHaDyWhkYCIQNJqKQpEmkLJ4gtJeluJCY1OrZfbqvuXmyO0Kb
7DUkgV+Flnjvx91D2z0zl9z7a/oMtemKPxo5aqc2bB7jcyfYgO4cZWvXH4gAhVhHsIztZasB5Prx
L5ScyquX7fVtITgUedmwcV5qQAc39+lvPogf/zmuRbzrEUYDy1mirpB/D3Vb+qwfjlfF8YFVSw/3
2jV49vB/9/0qIIMAZ9N95sXiIwu48KVHvvB63xcnXVxIE2SbLxSANB3STo0H0UvaqGlNMEZBaV2v
yiiJwJMs2xR9iIsXE+cVN8agLNiQ5gsPkRRpO6F/muUw2dgtQzpj3kxZ67JFwmdohb5ava6qWX5U
9kcjjg141gauQL/FJLrT62WxbZtNkfKo6OHAKWRBpLwNqNOJ8SUyCQeaONKtbPrrIvg2tyNKI3WA
tXJbl8fgJZvdjlfMYyYT5DKLKyIG2k/v1KWUQBnNxc1mbVFYNpdObMRP0qcTWqijqDOfTa75kAHT
O0GQNjFVPYUD7Z77AeI07ca0slbOqDnDD+yKGkUfYWYoJvm62Ft3q0EdOcz78KQFRBAVO1KfMu0K
QRY72NwuBXvlpT1LGPHr6wRpohUt5yn64QuAgUJMr6T3YOIiAFrk2OqwcYZDEt7G1rqhardK1Fte
pxR5war6QGdXVrBqjtQEwc0rSx5JT3nTFi8X5zU8kNz+3PUAenLRI5Ed99HHgfP5ieth68If5kSd
idVuBun0Bkdo1GN/fYNU9DqioeQRKLcgQkm0HkzE5aENwCqj9p4BmUQHByHNZBnxklQg6Vfnq5W2
U36uTeWk0UqNhJZ4N5zz64TE0YBZxbdjdeBIbaU05cA/jOfcqWc6qYrln7W2EPrk52a9iN5IIHAF
CocwMKLt18rXzI3Yv1akJjEuiyS3+qfasPg/232GNT0zYjMGYVWOplQ0xrkU6dAM2oeSuskIiK9v
+BBlfZzv1hPZ+3L4qSO9QFe714ywwhoI0aQxJZPStL8zrwcSWRSVUZoPEQZAG7DzpTss55mDTTL6
6JNR2vjrg+wvLnnhIVDD2j+uBqLf7pTI+9NOEPD7ibi/ldQcm2/SdnAr7xQtLakU0/u23q94ELk2
bvwg4ctBRe3vJPRIEJPRGGKlKi7soyvTArKLd/NODbLqhtYrMcXMs7LbjTp9RVuZpvA7xPsiswei
bqhL1Rq89Lhb3mOn9BOIsBLXMzRKtGMq6Q0fZ8EXAlbdqMppS24fcLRnNYsIKCYMeqlfvRTcQHzY
9jFgtylOIq7b2asVnUHSQnNrD++bkLFU2r2rU8LVNBteGNM6hHjufD9EJe+2pL7lBO5YuIHOXMTi
DrSbitqlRUODpQt8vGFDQa68VaIRje1Srf6y3vt+Cw84kUj0j0YtL9Vg0FaTHSRup0YGHlXamJd9
tckow/8XY2hT8y/UjN/xpI4MzznpFVz2v1IZsJKhm9+1vfK1lmOFxhpIlmhfOYzpHlgEaWHi8BG3
6T+rJwFlU2skx4GbW60ynV0UAAONEs5/eRJyjDb8HoK8kMkAY0VTO4vwEy2rxn1kxGzVybXijpbY
M3STetKOjHx9TJSh3Bco4noPqpcZ6JBzNm8XANsuzTD1hI2EEbUEzmBahT20LVTMqM1H0DPJcWN7
UjjFZ7OWjUgdBSsNj/wCEnN/JHDI2WWMsG7yl50mylz8nJfCIc/CiQphcPQ2quj7KW9EzBOIkP4Y
Fna8Kju+zHBHNBZsY7OWNeDLWUEkwIo0mZRN838DgbLUlJ25llua8QckvgbxDeJjDc17j1cofa8f
Coxvslny4dx6YRACopct9cfJEs1fl9nzZubhTUX8q273sJc3KXwLjz0eLugTtNsSQzMSW6bLjns9
cWPKHFbmzYUdbK2AbD4ZIWJJrQHR8drI9KD5IJK0jPYb0Fs3RxxzPq5lb9LSlExbgDqvm0g+2+yT
JviKAelP1MPhN5MgLQFi2Gk5b3aYdfbt6evJU/O2DYYf1r6PBXPNTZMRnC9E8xOmSZeA3WCnDsrG
F+HQOkf/bkmAShPOxmfS61cMLcy0QvzuClTQ/zJzizo7tKmu/iordwET57SPDXjGi9XxePQ8uRA+
cGIMaCPmXZt/jUkctu9RLXnu240AKtdSaHSv9IXmxJzCpOeB++lD1HgkigHXahzun9R3/RVFVQU1
sPyUNrviWPiPg+Sr+Y3/V3CtDkX6OSabSQtl3UMxaXMX5BthxjxEKUPLtavDY/lmDjLNwM5CDQql
Anr5JwKoNRZ62DKHmHOpBxmUChj4UpJP0yeZNd0URJqKTaFD1pLxtSfBYRFWYSxenObPI6kaoyes
aK65Z3/ssmH45cJn4VVIPjFYCgz3MDTdjNwfc71F2KzPN4EyjBgPeyIllNKUpWjbpv+U048xJ7RC
jCOaiaFVWsuN27/kiQgkPyZZw5C0NLr5ttFHwf7VTGJHBSVI4BV7ckeXniKGhhglr3f/CJeUVEUw
a3bEZV4CB+x14iPYcm6DwGhVhcaPkciRMSc9F+HXTjAR2Dpc42+mQjdugAFRw6QapDy6xUpVAoHx
N+3zaq4I4hYNgKBVjhCX/LOemxm7+jJeFazC4q6yYpkTodlwVmAJVbYTrvDbHFys2riY84lhmspm
EuwG/RyT+/dwZoyt1qKo9JPJsxo9njY7yi1GJtY5QItkQ5AM6BOx6lfOvXYLWyOf0NBh9pEeok1v
KYqz8z1ZIzNZzNd5S6idPG4MA8KTUW/6brCuupRZhVakxY5c4byt4ZhbL4Wl2jpq9Gt08XiI8fxf
zc+54PTaU2S3H86QDkV68oPS0p5EBkhi1mLs98sB9fcBDFctrM4l7GFz/sGphAMFzTNfOSjfV8kB
n2XefVbfsDgchmFMdoZPcrI6WHBDVa66gcpIcWnrGAsJSMNwaInewtaMAwixQfzRVdkpTT5FPMaf
RjdXUxNVgoiH3ag8qMuRj7HomEOCkAmWz78I4yWSAeaZIv7iN8bfpHaTmZeY19KuUhIoPykG/7tW
aQ6CxrLG9KphFDKuF5NevyPwFjvCwKBokCtogN6xjy+JI43cEl3zvnJE6LzoWzvxz7Mpx5IOuBtY
eYRgs/zAZcCfz52/dbulsZ6xXMbNZRf21NpSO1lfyWksBThvQp+W+Pu9qD570H5Kl9ORs1UkVhmy
05YgAIRKcTeolpPPWPr3sAbXH0E/nvu9PKUpsRsjb0euqcsnQVx7Fgc4mrm050hCGcBo4y/LEMtK
1NIaighSxeg6W88paHTetWm3Tdq23KGuintN9rs6+3+Sy7SJ2k3vcciI6Ww+d0q+Lpv0HgBPYamq
AXiPsVZ/JN7YIk0Ld+3V6jPxnGEL+CF30uCN/Eh9WXO42ao+l7+Wzq7tlPsTOyFdsuCPRtp81tPx
pwwgO9nqk6e7xU3DbnlJvONktsjZBFCbzbL1hpl04cIAzntg4ztXc0465SX0B61gHZbX0ICo6R5f
oMxinwX8VnrQBCwTKtRNAzmSMKwJaHpVXG1efi0/I1L5yHZFY7wO5C9i6rx7ZIyN2TkiwNm7R7UI
UYceLsA6dByNhr4o3yTrKfeZKwrrlheyO3NT4/Afpu5TqDEtx6B1AKQIMIpCyouAR3OMbzXPc89B
ttFaQEhg93Y28PtwY6omI8iVBhXBFUbLXaL5M/nQKaGDLyKJiZRyAjYHJ3xeKftZSJxVXi2aPnfX
ll1gLkEE3vwV+QJ0OPaVnGm+ycXx2HHW8o2/60PAlBlE5uV2yp29DXrazDd91rxA5QO9pPt/CpB/
fGCOxYR1dvCEOssHT5JxEJBIUqvkjhiQanIng/XWf1PmUJQZ051oIDDdTRoqoADB1XXM2ayAAIsR
tqbVSzfccDtS8Vy7UJ+Drj28Ln81egVAR6/vDOabdO83wc7UFQz0Z8Sm0WLKibLLu1Fz1b/X7hYL
VhM03kGEJvCRdoGGept87zaBk94sSlDXr6a+uPR1Dc14AvWDwslcQ+mxGYDbNXbcpOMCWvPLh1EB
xHitekdlVKaZIlg64NYUmdRrHrS2cvuNTMc7BgDiI00fRDzCrAif+Gd/hlnFJMVDL4q80Co9v+AA
9CuZczxig9NhID72Ava89xkim+FUTrJ/bLn4qNVTrgUOzqh7FAng0cy/y4R9+tICatkgs3oTSk2h
so+kVzPLnqdCHTPYny+8QfdU6RStvdXDQ6L78q51nTDjx4sAPFnvkEL6XPaICI3Vds7tMc/EZB/L
XHOYcQwnW1p/1KKBlj6IEe4fD3Ee3WnfQJEsgpaSbovCeU/u0eqk2LnZeNzquCPOM3CFcKQaplf+
CfDOc0Vryt26L0U9NNV6wBsLWHzv0Ge3WB1pqcx8pK+YQRZxe1c9TLP7G/HIdwIHDFSB82J7WCoj
dExXOM1xhT3NuhOYBGDTdRLQFthSGJ09GRIn745nctB0ZPACD7+FQUiFG69IWE0mG349H5uR9V1S
Z79xaDoNojkO6mwY2mMkjaQdUTBd8s/p+KFvZIuR8JSvyUWogN9aZXBe/33yx7921qF+bTwLsebf
bmTcs+wwpt8Q0B/dSw3PYysyzvRrGVX7HARjj6DyKhwcjJd/X4+sdNeNSLS4UvedXNq7fI4oNzs6
mpBNC0A6wuVsw03Y/w5cMeM82UeJsjTUUjvR73MWhHAtCY7FcMod4wHMHxiHQIe8XNnbjkcibh41
sFOJx/IN5Q5Yo96bI5/seXfUoLzWi1sdwBvXnweCuSB7L4CHptAvTxZr4Kh3H1uqat5doIiJ3r8T
QNXJ/2RjrqHSjehKClc06IgKRVVAYR6K5s4QUMSRQikH+NDJJM1w1xKfHDVpboD22+TgWiw1A58f
mWF88Nl6QhTi+Yu3nrjuU3NiyVOtt76kks8MA8PPVKwhEbwOlpFY2O7y0SM//48c2u4w7VEh5SbN
THEbhQ9cZP4j74M4PS6PmvkyRhvVamxsfg3AgOhJhuIJsHjUcs0KQbVDtk3TzU0h4pSCHo8B8NT6
EYXGCgaL0T17PikQUZysCM4cnP4nl5GSiW7e9muJbQGYLEelJ9dV8HNsLz3/RFYLmGnWqgCBdx3o
6PRpdAPyOmkkXiRTO7sQKRzKmYanlyRyv0ekWaaRgEiHZwKM9uATUJ32jozkJw828wdp/y2O+pBD
xVsAUHs2s55FoIjo6I61TsWYTiX8/b2Y+/G8uleevefS70sYEexc3nGeTOx2g3J+59Hm8rBXwo7l
TeD98SKfkcLWV3rToVQEStsgecmH49Ixqsw8bFQUZfbTs50qxDzx7Ejls20u4rIPfVpAql/dhcjP
P8zg9wp95uQW4A0VHbIm+m2KUJ7dhia1SazSdAJuIIahYwpMW4uEIGWcICOlT2Iy4iH7HBIA+tni
25Y/Wbq9vkox4EHM2V2wIg6x5xsWUBLgC2SCqquqA/t+fcEBcOYbInyuh+OnBmtUxLmlNIwo/EAS
GqaBge6n4LNN3JbNAE55rCXEj3PITULYdM9cahFn2PEypAZlzOIiaimSTltGYiAq6HYaWgQIA3Gh
shUbJ+T0P8OX0wiuPV5uMK/X/emM9lfV73aLPGE1vDucTao9q4cizF2AxgudKjoRlFGYLgqVqTwo
6X0zBIS9TXlB/eFtG0R3yrwuSNMFaiO+CtV+egLOTZ3rN18gzNxPHnpkbNG+3nn1MPCTq/tZGf66
BRDmK6OxuIC6v0pILeWFyGV38PNBw2TdFjhQmxHLWoVPLLUcHTMWFdMJte6fwpLX7fitVF3nFmNI
1i1yoq5F+RmWx0dDEOkPbwSHO+ktc/wuADTIjDevfdyP5COUm/I9gj+T8RejBQtB6R/C6Ay4LiWw
h4kP5drwG/Mp0Adiy70n5GlMdrNHnOzqWzfoIIIGaF1Js+alI3K+RsaFomsvSNtfVQyMcPChfWIO
pS4ZzF8opNy6fFjdnxKO05HHD+0fBPaaYBUIjLyBP3aA3mlAFq1leq3zXM1lS/XPjjiLyE7jTGll
kSZBfW8FIKaIZKYT632+qLo5oJ+7ocMUtPNExVsf34hSFGYXKWp05aoGiVezVCQIzUsJXWrOSJZE
VB3DPnDp3qpeRrES1T70JycY/5PS1MlYSYoK908r72q1OzXQxTzKqtfIMW9eGlUoKUI1UheWg47m
3kvhrrwhYULb+35zs6DqM4q12ZVtUQ3WIptK+RF5om0iujFkjnINhbw/RH6PD2ClN98JkQK31pZS
uIZ+SC/GRLBh4UUhXN2c9HhBCexBc7mvQTdHlIxJDl01F+1A6qgYzX92pYMWslp0igNLgH2gvzYB
kBWSnYiQITouzc9GFDzYLAcDB+TCzalOrysS+GynOlpGZGv+c4T1iral5BrsDNwb7vor90v5sUoc
tL5zcjYBiuo6LHQU+G9h+fMEKsydt0TTqrAYyoapK4lw7EJTI+Yoi2MnO4ShBQGpE2tSP9xwu/Ai
rWzLkoHBQuIdrNcwIosKEa/zi7iBtkiYFsntJLPKKW0vw1qPrt2BMISzntc4WyiO0SPNxfT6zbpm
qVRBy3m9y9ZEvlqylyPtmlhCrmN9L1Xr6Mc7W4ETzD1WHM4z1/8+4OgsW/M6foNXzs8AEjspPGXW
4WwVYO7ZZykUSiY4HobhOJk7c9XDezpCHQAVMjmeDV1ZthzcPyAPLwg50P23dK66IxdirYMlX4Ve
nzKBkJOokZ1Zuzv1rOgZea4+9k1f5RHW7KbLEejgbx8P48RNvkOyq2lSVTB2PMKhaZvmtfvoT+Yx
hHxlQ++FaSZVXlVQmImc3CjiqTXxI0R4ppK/dHx9wMqrnSUxsGexyvp43GaqenCax35T6QnKxGMS
nwyzOQIlgltaCuRZUxuvBCbWJ8FwqVNBduobs1/i61WmsJnhqhvgorNMyZQGi/yY6XP/8xaEK1Y2
FmaWDk/Wy+MqkU+orlfw/d1b0Uj5BlfJ1o/iM/DhZYNy4UL8H8JTUMP1iIKoFZyzAOtNLKNtqkxI
MgWP3sbNXJknrTAb0gUa/dWE0TpzUHClyg6lhAAsmeph5uwqyiqTPwD2RjRg9WNk1yOYq1nA3/7R
pLI4Ut9+Pl/An/jcPA86iJBomJ/k3Jw6CZjEdeoo3sduJvk1+0cQuusJq65xhc2rWgm0FM/BEjAY
AoKED8rRP8haRwhn1VQ9LzZvYygRvnuIjySvu4dVZ6GkQnuiakaGXeTu4mHKG92vDeSBNcaR2478
EdpX0ydzVDvb/Y84CVxXLKs8MbLPrYcfk15TLp4AZSdBnxInDWtoeOhLYNgEZkEyZFWlz8hkOMVe
QKDPMBDGehNoXrzrqeYEmnMgblVYoISkqb+NSqnU/IrbNaaq7JJPhY15cpfrvO8Ntx8pZKcs6KxG
PBmTJV3kLJdglZCmI1G8zuPNaNQW/OwMSd1R2tovcAnA91lHKj6TGJiAyYiQA+DUclqv5HBsf5xo
28YbYJ0lDQTeJAd4c+38/08uFV9eJ5mAyvec8WJEe62hHHC7p0lVoGauijxPWOZI7/CQ6zVb1qf/
wUGNZCzm9uOTpO/MOVgPGIiDw6zFuVZGbgs1IylfTdqUaBVELx5iFdHp5QFpd8KxPttc8swhowXu
T20JOO2MnM3Q+E2wZCtx82hS5DdEsx8BkFVNjKYsjqsdradTZX+tKOTsOjvCtrNAe76TqHk9lIjA
m8uespNJXLoqPqTZHTFdsuyGhWlq5AmAWVZKZ1yHmP6rSlj+rCeDI6/sqGOUvCTGnK0wN4ob6sLG
k2OHuBQXSorO5CXzD7f/QK3SGFMQITmttrHMFmaeRKkuOucTNZ1VVJBovNeQ+tOs260kLM30bdKt
cC52o7zZ4iI6PzXhJ3EUcMhp+dZQrG5Dvo1KhFLEMDRCePzYW9xDWsVnfyL74SYjlvWdyFfArAVU
rOFjdrgc6XXXvYQp10kdMzOfGqJk3WmqvqAG/e7IutZn2O3XlzBzYnowg2L9S56Ev33dX3j+gukk
YwHHjni7Vs0y+BeBq0uBmKCNbDw30FmBhMaxKeOSJTfEMKd2t1THqwqPDLWAFjwceoE664Umqyao
xIm07N4lZ7eOilNg7q7VrcWueQBS82uO2NOaT3mxR42bxvih7zmWO7DWT3tLEMH4+z80pNQ/foFc
ZuYD0m2DlOO/1DShJ+cc0FJxLlxEEbgLFufWc64mzYe6ymiVxlOikbwy7Yuq3azyvHU/uYr6Vf/P
ck7w9fHfLSsDirDlllnUO0xPphPKHey/3d1OYXgYw1FdDbPQNZmOsn1iQSlK/BWXjuhM6q1av9JU
YMLcdbVY0ywFhd+72yv10eaxUtNVWYWWrrLTi7/QbDb5jwPFjQ5T3rOOLX4Z7258h2489+XEzdnG
64kIR7TQ+vUNZkU6BwQXBZGB0kwhAw+jhGB5xIdJBKxskggRTh/EY73EkfjSx0M8LJdqddMDoZK0
/B8r+4TaMwvVoHtKuJt/9OHHjsIllkP+FamvqNAVQ/fpxEnWJ2FViJM6YZn4HSZCJUp31RtLYGwU
OHp2ASVd22pLO0fJxXJ04ROB0pXmaEbgv/UyPBZwoeWPA55M8NjCHsCqg+oolbjrjpTayXrqPgTQ
kfdYJNkJ5/h+uqyEj32xFBCpi4fBCIZna/ln8oyMd7Dn6SwnYxajJgGvWvWuV1096ZrAKWi4E1+l
oTOth6UN/R78GfUBPs4k5kxQrLH6c49elcKmkk0Hj4Pi+ioDUAk046GFqh3mav8RsBt6pQV9g6h7
to2rvSZ8RQXyn8gS2yhIq00GUgE8Q2J/arwcBPazL4ZURCaWX8fy5sHSUrm/29k3wIwSASl8ykVo
4rz7JSssuRAlxPLRrWEedejXMZPD2c4DMzEtLTNY084qdCjc2gjBciMmoafAy6AQiQzrcFKbCSBF
+8eCoD9Tqt1P18UFxrp14BU67ux2Qt7h287Mz1jEzlDXc1PlG4Lh76HJLXxMi+/wHAorClWOBLlB
h1G5lu55L9XY0Uqt/GQgfEMJcBkRyzcs7C7xjGRAO83cy2NHAQUM9HuD6Dn7YiUZid1ILRKIEioa
fqiOX6EzxGHT0zaaCBYJUYJvZW6LVRnIIqzlPOwrpRU9uTzAB16/1xNZfG5IXagKduIhWrhBc3Np
JIbCTzp/MYvOdx6YlfRUYLzrQGdEMECkIppIYnqkskvD9lmZHxAGHgv9cJZhKwuEQVV0WmUKd+XO
V0FDAY1m0wu74Ye6BrQKWGRuVQMty9oJ4XJagd0HkTOfK/0IEyKa7OY0CTugRNO+XpAepRn6LjXp
tQnJgO98vwWNgnpfUsLoL1J8BpWLZFJaLKfUAaA3YqZq6EFQekztnlm5sTiw9DeoPdsdwRkSA6BP
VkBVW9O+KDtKLfLo7FSTzJQkCgwrFn2nLxonwr6eZge2/pGVOaIubnE/GHoTWTRJOmRdGClBEgxM
ye/ZbMQrAybQQnWWb98zGyLzIeXQMV3zXxAKNZ8TNn9lqoNS++rlBTlY4J0qB74anzgAc3iq5LDD
NFVizdwnXowlbhTDVbU3E0z6D0ngmvfsjuClOy7wapun1sBh2LnQDaB26fCjEabdYhFNlr3rrnWa
mxBKse9MS6DzBJVSpl9pJAmyxtj7gvg5uEzGEzkbdyAzQXCrkIFW4YOEgRi3kj9/0Wd/qgTl5RBU
GBdM/QsRK21T0NjbDmj5eZMzNiZm9oOTJ1TwPVefThcUQv4NdlPqlpZNZ0256ku+VvOqbr38dnLa
kNCXUnZRcubSDSj8XAjec0L3nAFieifA8rUMSt9BPL2bVTuXVbqiV+ZMbqUOadVDgl6+ax05dROE
kzdd8kQNBjQF/HCDPr3Xw3MG16g8y1K5OpIoxD+iNa8a5nt4zvSZJg0CPUtIL9QhB4eU6v5ndYdS
JLzS4IlYDWe6QOlWi+reFYyspXip2BHk73FyutZf/Nm3Nvo9F7/T058KUPeJ0fdK/mC/YKB/uuNU
DH9fSCWXqrIEiXBMXwf1DmZYjG1hOeaYVeOXQStFUTQBFwq84Mlz8VyMcf+uW1LGMqkLe9Rad+Mn
sOhG/3oQa+HuFboXS79Ktejr3xbV1sfD39fOKsJN1ppjODKzlibC7KFBjsXHT9rpmVfUsvlHSS2B
2TKJm49DdlzgyCTVEx4QQes2I9ZGfWzIy+RcxLFPvircz0m79h9ElCXjVi4Ws0BV7lPuSBRThS4z
AyNzhRzqEwZgZZs1KbEbAJg0TfnwpVV5mU2ZQyY/RrLOWCfPFMcAR71TENx+tgx0xp9TvkCWwlpI
gim8wzo7V3paCRDiHJZ4pDUlYce3cchDEupPzSc27GQ47vUhCcWDHmmvZEJ3eevaKtcEEn216Fkg
Jnn8RPU1rusnQ41UWl1ztBa1QxbgifGUDmlPM9ZXIBF6s+1C/tyLw1W28Jmjg3cf2vbMPlg/rRDW
ticFz2e/Q//gr31KBC/YxrlPNPbTBzosx9PxVmMWPvzYamLi75TG8pZI/GeECPCPraO6W2lsRCeq
ezGUEwCoz3d5/f++4yWNJKQiTQh+ez1GCHDVEUh19o8SxKBo5ByKckJMUFjmKiXUiD9ASj2dZQFV
p1VH1UuihPEImf7IQjN/UkxdZ4XAXWPPVE9bVQGXfNWO4hq3h2CzUIXm8l93GWfDepxRc56YwWU0
gQfIOB7sgNIST7gzLPWNZeO98vT47Dv66EGuUPN/P/b5nrKEA3V/60/MmoqHMd//sXgup8Ds4t3s
RrfrjObxk5KfNHo4Gd58+nhgVIW1F34TvKqd7txggD4+gZDOWM9XNjkecxYCN2zheStRL/rQofC8
6qo/46vCANxvP5mhz2MTq2PGEjaBsonk/ZMAcT5sTIKTvhEVWtjWdFAasQGEgfLCJLOl50Xdp/aD
2RvFAeVoWLl+CpmQTs7asBQ1tc6O+aK7NNW2gmaq/bo55YnvCpjBUfDRmNQWjeAwLbDbAG3fLYPW
6FJSm+a4/K3Olvppv+GMYW7TDpaPSIUfoZ66UzKFzPLq3Dht3pc3ZmA55HSMP4bU+kDTWIWK28ka
u9WNXF5MSANTK7GujdKhyXK82e3niFyyQglrzj9LxCLjOt69QdYWNcIQxHUxEkWVSdIBsswai0eq
3y+pd58T9nOrGAuwEUKT5W5Pct5R1OM3Cm27ojpPziqcrclh/kHqpNN4ccxgoGmVVuNqMeKMF2vQ
bR13/dCvpfA3+dON1NX1Xbq9iCO5oPB+xpdqBz56K4jHo9YiT7R//7ET6DsA4Vc0Sy6eJkdVddoh
Wz366pGnURqgKwnwp9gOIZVPM8Mq+8HlRh05d0ugE7rsYmcQCPoDv1U6D4SjkuyNZ1tdzR8AIlUW
yaykgLIYb6oizUdicCMmM6rPkQhIzjoKejRRgjCxJWG2NLzBYRsakXYfbiC4Ny6Gw84TF8/LFJIB
sXZu8DCtKh2vF6MyrVynuOs7xLiY+fE3dH3DpJqku60RFO4OrVGJvrnikDLnoeaSFM7BpEi3FF3u
Oy4RlaJ2oCvx5u3IeEX7Y3nUzPyA6sE+eEi8PdikgXzYIN8gP+13F9LqUoTS7fzpq1GmeA4hAjds
i1m5kqvVI9C9Yu8UcXT32hwjZAEM2/YjgG7iNPq82YalDHK0Q6k2lsAnuJYHw6w33VuCjWacGqYF
oKh+CYqGE5GG8rlFINys1bnhn6zmI3povicyoIDSVqJhqgvlj9/UOVGsoTHymdJADSdr0kSYFKwB
n9ROD0caLffGdEMwndjZFJaWtLQIamC4SSDox9WW9InPATBDygVJHoG4hXgiBxGXptWVDZvojFZY
bQOXGmMSXPn+72YCZdilvrL0V4XhjK9Yfzg4+BkDia1S7aiCn45F/oipt7bKi2hPSTCi0wZF4332
KLRjcxS1VuSvPAJ5MIE2zlPTPbdURsLySsidmaHADglDHrXtMTHESoHFZEndsd2z1jKzZqWfak/p
yBc2e6QCKGZVlLpwdG4k8IEND5VgkAaoNFKg6gmXw8CC++2VPyhL9H0Dq7GvUFWjP31/s7poIl/D
4qyQQT1T/zn8EcWKtIQyVFZKj9S8wOCcV5CqA909AyDcRWjG7iv4IPR8HqX+uwk8iUXjaMXO9Xt5
NF1woHuH+wooHCY7aBfeHZ+ZIjK6CfK1G9qTm8olSdf4+NnLYrf5GRIEnfn7LuhhPxTJap0EOI2j
YMZVs1Ip7wMRq5nRrC6liJZZTdhb369Or577LAlrccJuPCPs4POF+b31JJKecZ/QjsM/+1hzTb46
hp1GUkxPo/bXssgE7Ix2KuYZt5CMbdnN+dM5F9ENQT0hveCUmCFDsCn+Mju3f88BVRbAUfSifARf
GHfemt7BwLPXFhfDzxXKuyiAS5GXfbGjIQL4nhStRd4ywvvWP1WT6eIjWSEkiUOshEYoqHcKlzq4
ZpwN1BrbZQ0+Cc52rDXDudpXiFFgDrrnoVHdU2gjYF8JswaO/eAwN7dhRih9trAbMH3jaXnssp2U
Cf83rRGZTvIqliK9uC3N7o0+rm+4KeDgD8ZJTAZLAxraLEUnbwltoiBjEGcHS+SY+AKdbc/U3YrQ
b9cAFgH4RK+S6xfrdmwN1/lPuh+DkdNoLdKGn45NlHrJR5god/Q+Kb1PioVzsz3jjk3CpjhoFnAx
bGdEuI8JZ1q6p5T+g9oqIv0rp/rk5g5dyEZZtEv39px3ZepGwbkC9Mo5LFxI1u7F7HC+IqH/0PBQ
ZXBvDZDN1WxoNcG4j1GECHpvgrQn/Kj++JxobkrWpE4qY0vRq4if5hO+Ngu9my/U9p7sV/HNn5nd
+lz8UADqzT9lDtSI3VkSZe9//sPtZW8jEiZVJuiraR/kKaSYviar4Mp/VdCqE3tlSU1NWiQAkvWL
5D55ZcaJWRQFakJomY3+C72whTP1Rm/AyQkfSk1NrwFqTFAoqCvRjBAv2ghBXUGOkQH1sX/Oe+Kh
mvd5BdkBaVWUvuQGBr+2LL7Nx9190SP5xEjplvdycW/5N9+j+Cd0k0IVFQxxvbS9DZZlBJs1qbR4
ALC5nJtdq0mPztBMftIJmM5MCJTwRP7bo8obmVpQ0prxR94v/3Z8Qi3yv1g9x6uzGsiR2yVVXV2w
XkGdopEaNhFp2YdvjTV9VgYEPP7SVSMnRPwVDrg3o/FCHJq+iuiSxZA1oT/aJ4hJJxpSD+4Kpgxv
9gtkUMk1aePyOBGkmu91c1wZEk2saQWlEev9Wh7L7P4zMxm+vVBjidsqIV0T4sNKTwRGLr9V5+IY
WYG0jnVKvlBlHsiYy54TYoPkfIrKo9bb0G/AvIgHLPy1gK1u2MRotZ/nf3WLAUGnOft/z4Gda+8+
ddxqARidStr1m84iijsHbqyxvMeRZ1m6zAkRVHUkg2hlkckxvUOcpoPQi4EsG8Di+7ZV2uEF8eMY
90oFERZ6jToa1+cBVfJneKI0Tpfb1A49+kx72eu3SYNy4yP/jrjd5ANQm7GBudnPLP1cmS4HM1jg
Adanwj4dm7jiBL2bj95sLJgdGNqoGu2EYufvyB7lPi46aU7hOFkLaWpb7Fbm2heDEiV5qRNnhl2d
sGmm10GHLtXhM3oVW4IYBjaFxPJuTTTl6Bsz5li4dUuQNQuwn5uD6hFeiY+Rp0YmJY461/t6EszH
Z+oT5DAVFWEStIVFrZ1BgM2rkFA5iBLlHJFY/DTffMd5u3sEl67c/9legZKSKUUYsuHup5o+eAUQ
4WpHZOJQSHu9UfU2WKsEDC1kdbLH+O1Xph1vlKSrb7lip5dWgEM7cjGv1Rb0mL0bVQ5VV3futZop
kqHHGUgu1N8aa2LJDI7SfVUhG9T5RM/YrEH4gV7GlBuVKF8fdbp3hprGre8xSn6C41E3ai9N9lZ4
KFuXyoUzxPkyoeF6FzyaWeHUmskRbbqAMld/XOBoxX6b1HItAEAFX3ZUiZ5RD00BlwXynng+mqnT
coFIbTQ6JWe4gmDc8kigix6iqtvspPTpY/+2/kear6npk5Gm0zok52KPxTqICj/SLS3PXcgZrf7X
TG3GdAiIPOnqadjAzJRLOQb0BHI5a39Quh4BMAhXXigZVSq/LqN9yyj96z1JwE9byFfTD3ucG7YC
xn8EO1D9TgVMBmY1V8X7oMP8evFZ176cx836T4pGIhqTKEWexxRnrNDEQVU1Bzkq7ryGpDxN7+Hm
EQ7CQsYKjrj5DVF3WNbobQ9QRcbGemgE4avtdSbPpUQ/Q0I+1J1CqeJdQwS53bErmyLVdoc1dvS7
Ci6TI4ieOa8ltAF+3TTwHUagzdyz08oiZEc4eYkcSTSou4rm1tcnLNBpYYE/X6VVpW47da4Z/KTk
FPHqOMSc94QgoLyL+zPzsin47xMsRIUPYJL4OcRwE6nSfRnX/nx5e3tA1lSpIDhvz8hBbwmFoXpj
MCORNhF04rUASSt7AylNuEza2kBEL5CaoSUmPjFp5/20Dpj8YFyuAhoLIRD84uV0uqETsS/PF6vE
qeicvYcuLiYvo2XeXffmismi+33KkX9OVUBBV15+9/SUq+0nBb+zEJKoMb3Hwjih2JTqw7h5X81A
VRHYNmQBRHnjSfHIkgFNZWu70wCeF9kJBqRPqbx3qUi/J7LIFUNdL59tHFy+wP7YzKv5/23fOuHM
ojjtOHUpWPzwzFPYWekCDCWVU65Eea1HPuJwfz32tMbDUeQX9Da3pvH35bivIRKxDfz3Ra4WM9nx
2XIlEbEDGuhDCAD2EBOXfS0vWlR8BKM2ffwR0AvQSRW3VResCLP3ICHJWhkef/ebf3IWEdZqojjN
S/97drbwL7WaM3PioGApLFqMQre4hQqH1Fr3JdfShG2hJBkd5FckffPkKulbdi0J4Aq/zQLpz/K3
T11Mog+ZPBNzoe4jwZsNsBF9OurPx0VNLH6x1Ese16ukYxD7qsUzK4P7VdgvZ9g61mrFT8Ar6UFZ
a+Bpp07pUQMBKZM0kCRMRSY2ItWmr02h9GpOFX/sqTgL7fhQdc41cCB/w/v5cLiJnrDAkyoWTBdG
rpfJJYXD9DQlPH4mdh29Csa1aJAcCzDB7sfHngWaTop1bR0VJtszRSzKqVZC8jzPUrwG+d8mOrh2
ffH3oiNZ1TmKPRBQvmVvcZSTNzOhI9XiUg/agdJA9h9DozPUiDS4IEFj4gul2AMAug7qGRVgV83i
P+40nRb/Hf5OQ+zX33Pu+Lkj1SmS12ZcOfnxMugxayp/GB38mnfW66ieuhVuQhNvEqvgd1XkJPML
dFi82wnHalf3TOwgyFIOuurQC/QzGY+p7pSuPho5QVJx04CpnF6KcCqiVqKGa4hD/0H4DelNxuqK
fkcIzk8nh+Nwpo/wW+OVEjzlszHzYmdz7+zcc9EQndMtpCXvIV0hhGLVUoDYhAbLkjdhBdbOGF4U
TT4Q3u7sN3Li3/z+5gP8Yu3qVgXcNOhvDZOyvRb6tXi0GoJdS2XUBdOmw0twjhUWaf/gar+RGNBM
2SGmPgW69bTHeN0viq96EsBHuIiIWaWSYSAZnKLTuOHS9mxgOzkJyiJ3w+SGYVVuLFCGnG/mhvLn
84sZlkcfvCtNN2eb+5QT6lokUgPzYxwf7qscnD+VB44sgHr9VoadfRtt1EfLn35gR0GTc1uWDXEd
A09jgnZDYhfn2qhUthniMYdQhktZgvcLvTwzzUFioj3PtGmUaLWLumrDSeBSL6z57o2oyJwGl3Dw
leR0+rIlJS/OvcrXmBRIm0pBxWKeTPtLtxAUr657zHjILbhiADsDA3gKQvRKphvs/3/cncXnE1Y1
ukN+NEYLnmp1l8GV9moAdWdwJxBUYZ0KqY0SVvwOAT92RWUcLBvsss1Foq6lSu0Zx71trdkOiCkH
eSgJLe4Kut3aJNOZjgnOFhOt2aR8KC39mzDRBQKTw0oVCFJpfdv+740QP9UzVVHusUDms7nQMa3J
PyeLBkOTkGkKeOT5/cRH63mdLFiU8NXAoE1VZ1hOM8C+QTcQw00vX2bC/fhanDqKm5XeJ8POQ1NN
Ayzhn/VVLjn2X2y7//x6XEJL6WuqumfqQxVcdqKvR2uxPADXXlSUsKUzKQ3meMa+xMe7iPP9MtVm
ilaQNIbBPTMX4YmQ2Eh8rxyxj0UKYR+S8MZSYE0HqPWKKz/THkHWWxjaFZWKtD94cE+7WtYyJUNr
3jsIcbVRtZ2SNvj+NakNw9KSuUsIX8TnHRMvPrZuM1J2qPH1zTmsNubHxwNpBknUG0/4TR+Kz4be
qYqOh34Vgs+Qtx8f/JR6Bw2hVAAIJYSG/Z0Cce/XQ9cu+VXznNieuF0UjqjzMeMLDPxLC/PYSC6i
RrrPOgqSTkgtH7I4CmQtJVv1aT85mJ3h8SWkXWu6JE6vCsa6Be00VfZCq9wVR3FV4iHgOtdrRM7t
HnGgcsUn2dfiHOT+Lb54LfupQ4NqMs1aqv7q9yT16gllnkJbhtWDlEYrmVkQjghag4rqUFgYbBGU
TjyCQAjDVZRhPTXWd4kOpMvp/r8xjV5L2H9rmpXOCWybTgCCOJVOLR4pyUZjpfZGx94tDvUjHyOy
FZxXI5UXd0rlLC32zLJ1dgi2VvLl7JceX9mCC0sJ+EI4noznczNDHZ01y05bIN43lQjxxE+N0RIn
SibKJb/jOBw1wt06LOekQGNv3bkXdPaoa5U9GTHfhdTlTPUPohWD8Ne55WGowLXAPKVy3UvhYhW+
XVqYDP+zBXA3bQvMcOg0L5ygRSbgjz+QZ1G4l1gDgh+K5HCULQYyRHKhccnxiRY4RTCmpjQhbw/X
nv28u0ku+lOHO1C2cfJuze5svcIpRVPoD6y01m4VwpMjfM1tYv9Sj3JiP3bWxc/czkl4kSFlN8zl
LDnnT7GSJhrohOzdasR2FtEJ0jEgXeUggf8gARFUL50FOW8VO+CRKIyEHZVqVoNt1UsS1CELAGRJ
7mHw7l46o2asmzBCJi+7q5lOr4jNe/oOF18kLR+OuXSD94LxpJDKmHF+H6sZnnKeAoYBpmOpK+wq
bq40/zJmshhb+vKGlIV/LoqUJhbf1EfSZkbjHobgoAfg2BJrnkiUk6p6z4wR8tiOzb7kMWo0A3HS
/L9+dCdHpsz6tCOxnnJaqJ1pktMCDO06HaOlJaFT9gMhJY7co8eJjX9GL17n1CqX5Iem0+q8OAC2
+94Ouq2n3XjbRUt9p4fa0EhM/vFISMaVCrm5fOLxOAOEO67XziCLIuO0xP9mN/eNz7moH6FX4wF0
Xm7S5k92lNth7qS1b/rB7bSAEasSKQXZaNyCd30Hw0jeWAIuHIRMXp8xyDGXzRvvEq4H9qUG0scr
+3TWe5RoJx6ERxQwC6ELFtmpq3rRzp7MAGh+7qnG9AL4bIIbrjutbihd8/Nh1Djks89k8QwsUZ1Y
oI4RNCVgru8BAj8ZQQvKt7/vATZegQQlFoHqxQ3/oh/L3Kqmuv5Nsmd7f6FS5YDGAKNQx5COrlCL
eK1zz/3791RTrsn6L2MBCaZ2crg5rZQtGOukbM0qX1Ux8GdMuZ4wOOR5eBxS4LNY2cAvt4VUDjAQ
AFz/3VaZ+SUOTQH2vt/XvpjqkFdVaBynYB5e5H4IxjFZ4Yl+S65e4GgywOcd8mTBge+3MI6xHJXi
2KTWfKfB/6j3g6gaXxn1pZHHFme1ngbf/H1ptimXxRDqR51MaQxb0dy6DWS1ySy92ieIhJMen/jN
DDkhGL7BYpItDAxGISQomZEpqHQhT7b8+hfpLYSXjasAzIFb3BK6Bp15KhbAFpigRvH6JYv9+MZY
T5IcEldysM6KCRNUAsragBGaK4YBSvTk+5zMWt0zw+YnuI2EcIPWRpXhum7MiLCUPVPV7YC7D6nY
5cMsZa/jKXCtKTjhlNnvWPjj9X7+rNy74jWYX56vkMnbm01ZqXYdViinT3kADNYIdEQX94vdm4iC
SAU41d/xvf/0Whv9pXGOEVxNFVeuw14oU9BPRoI17eaQo0uDwUQ+tNjxeQOa1q/4WC9wN0LfUsRX
tNScBCtjtIUPYvKKQnF/3BhX+7cCUxFLtA1qt1p2XkIqmJGtd9OTu52TOLEnhM5CcQ/SQFoYd9Wg
1SMsv2UXOVl5yHKjG4N5TQ/fxt6Nc4KbItEM6pQ0XymR872OU98E/tnaU4y8NDCVn7UmfIrV5Zzs
kKAEO4CU3Mkpx9LxFh86D3b3Fg1k53HdCZphv/6T2xtx0sOWFeoZyXB8bVEXgWUm19lLkHM+ntPm
nvdChMgmJ2QxMvENacEm8WTj+nYuamdAJQpF9zYGT1qgY5jF07A+mgT1ENb+kRg4dTy/Ea0oqlXW
hqmtsRXMZRL8FFwWu6BcxQhEC9p44InVuVc4jvybJKJZjLPQ5XSMSUm96KiU1Vqbcgju3wmdShBD
A8gOS/UbRKc0tLkOHeURk9Kk/Ix3Z9uwf29uWKAyDSL4ZU3rIzUqABZAfnTnon4UcoCmGGOuY2sL
mmIqFfHb8RrgRRF35zTe1iy38fNVM2/TwnxoFTcXI/6QNEfWPJbQaKaERCjBD0Cu0PjrdzGWbDzs
9OwIGHVk84yE5JwXtpWvQQVb5nNhIfaiGbqTS60kQVeNID9OuySfJumqcRcy8NAtFht4J0Zq1/Zw
XXQPR3ZIY7eZWQx+IOsQuBmCbjbR4NzwWpDnRqlRiLD0CV05yqKc4K4ihrDq+5EPGokSQHfBRXYh
LiDD354jZYq7t7EJggEqqr9Uta1l8xyoYrMGUx8e88/znSFgqcvpxtOvfi9irJyGFNkbrT44S2OY
AMUntEOeahoUsbd4KNZ7pZwl73LcXZvf8QwiWf0nzet6BdX2G96rK9o29KMtjjjjQGKsihjrr+Y+
voNL0Y/hDg0Pb7LSiTOSpNhTYBJos8V/NoThcBY2tbadzQrwwDuwAMLkKXYgklgKjEOPgRvZnh/r
GEsC4Wvc8qemCV9hNuAatavdgerfLR/Wh3mfr11qkOTtLcSr9DE1v5BWUrYjRGXmwNQRGpOVVTV4
vUspr6EUEMntsYFq76LVPMrDe9UdGJ8ntZoE+HdaurF3j7qxXLRFHv1Sv5T4ICLhAdwUHyaTdMmk
VyHGjGa5k+zTOFg1p2qRsy1K7U6sy+tXyIjiH2n7VE/zlq75rS6tphutsThQTgVr02en76ByC2h0
dSvbR4LeQN7j9QD7xoWK8T4vEK+EnohOxvZaLdDMtMZrC9qBXseGw25NT+PzX6dx5bfBaiCNMioE
+he/KRFQTEGvg/UsjHTCrVZC3vT3NErSSSSIucS/tCEAsWyNyS9WztpCosiIQ9fPvozNYwtWTTsP
MjY4doUoc1/E14gjcU3a2oBgz0yDfE9wIFCwD5Iuq42K61Cbca6VXfDpY299nzBiirYMWUUTb60q
eU4OtVePbs/SobNS9kYCacHItsU8WZcTQSzYcUNsT6+oIwqbEwhQLfPUL8Q02yqJVL6iuQjDDjF8
fraaAxZ1yg5hEZ4g3c0UtMNFzP4J1iGS3OJfUMdjgIYcX0mxdtKJM59j9RdWWPCgPGoYuiUJSU+7
LVilyAaHTWA3Y/hubbvZg63UH7z45dIalG5S20uwikJHQZopQX8WN7YjSs3U0bBnNbp/6ZEe8WPn
J/XRCU8uqLglppt4+m6Mk+hw1/61MnVeo7YfTKwn3QHFuz6TejQUf5zK/hieVpUAuZeDVJrlyPVJ
5rn3SYc9yKpeSDN6AHSjK6UnU+K3xY1ipS5PMxBjGHox2VVObAjiU/n9QCt1xGPnOmDsLnvNx/RJ
U1TpjUHfRVSMsyRpFfuC8fYvAmlPgWYrpVgtAUyPdUhi37ofHW2K0udN0/j6U1TCAF6beVct8aDG
pPMClZRdqYN5VbD29jnWNqK1wd2pVNhcUxAauxOEdvu3ZyWCqQN9xtLMov228ZOk+JwIh7SOAwkt
OjJ22viCXF5j7ihfevHr6SpkU1Ug1OyDB+vp8bM/zw8o5ICjxMjwuBHOKCvgR/Xw7PqN2YKjF1AS
LEP57+WAy20s8br2SS46DkhS5Q8XQI3CctvjAbe/4ZU9MqA3BMmVKZTULOLDzpLPQSUH2LwW23wp
dkeClJ5lvz3uVcSnSA9uqyIAvjLIMde5Oy/ALNfwrGM+mm/PljtD9YdeYoz4kQ5UMNVPKq8GRGBC
/13wtkysBkD/DC/PAtkaNHoucqDFMjaXB7HVslWJAKzMQSj0eGO0c6P3vXz+CbqmpFjPF7M1x/jU
T4p8RCmC+UL/6JXnQpkIIGwU9Y6lc3lEINKEbYPOwsMt5utmyhFolVBmQ2XeiBnvM1jjwQf90/wA
amxZQy4SoeU6UQGNcoflc+4Ea+aAPVjXNyK/n9WPoI3CY4Mj7q7H64Qtm/IwQ6dFMDYX8bLcag+P
6OD9oDVwQ81i/4GYgUxtIyvzS8eBiQK4L5Mce11qVJ2lmPcfYwQvQ67Bp48+mAAmrmwB1t/kt/pY
0GEUuHV7gW6tZ+Pv9nkrp2dEMd6/Srn1Gpbzj/ySUE5ndXoChZ0TK27xHX2+LnQGO6kp5axFscCz
f7UnsedD9mUHmGdCu2ejeKG2KGCG4UHugY4/enwYfSlTFIK2Vv8viOnw3mImeQPlqhUyV27Y16zI
qI0UZuc0rKpcoL+DJxZ9UOB3cTPK1NXpguLFWWNwEMeJY3hPV3eGEiGVcabMFWngPjiaSl2KEhA0
OhZhx30P92r8CKhzjXxPlqEk7TNmz0rvizplJs4B3X6EJyZK3Q8OWxviTHIA3FOvwN2axxOw4hVG
joWNlElZBJ8nb4NciBmUbASMILUTQB8tFx2GdAXCEwN/7H33l6UwivqZzRRjSyA+AQV77rchJygM
4q3jucd51JzJM2VGN/NZewceAa4vmDZXQTQkyzxJCtkKkA7oH+Qjuv0+gIBWs3yeKvCKBQvaoKWn
nqUkad0wb7jrm4Babjd022PjTG1f8TBcCfURBpShTDi+9nJY5Ahu5K4R6c6K4ERHaJON52wfaoPU
M15UjN6qUCV5VY7mqLDiIsw3Y8D0yhzJ+9DaWL3w7ln779BUHipJoTkEYsMPcqWDZslJDqLaAab/
8vIIqOQkYh3zNIY4CbPrzSlA0WbAd2kIqcy5xzfLI4WeyHdz8Diqv1ZKCVcvEKZSjhGyQ01kweLt
qoLhrx24QdckHki0MvZOQRAXgMH53zCVi8U1xjqZMhEET/JTlkQv3nJd30ANiOf7a6pjGYLNk4ET
8nzR57kX7ri/0XXX/DGodtyq2lpg6oIrgl4QCkXzjYNJft/VQlKuSPf8KkY/6AvKtmwTsNgfXQSk
ajPeL1ZlEnYRTsRmmw++Kpgvc7XeVQ+F4XUARsjy+xBgKy3kC9L7In2eCzhRWW9MezSumt1gkPri
y+hPyOzMP95L/9N3t2NY3sizydgvCwQqbVftQEqxnAeZ/Pd9ooFfjEzF+77OVGmAtYqCT3bVbPOR
m78HkmXkuahQrWzcBS5/O51Qk/J4LKDZSHP5zIGXPdyZjsmZNt4CuV8IUAeJ/RJ6ZF84wW/gzur5
g5bzqrDu0bd7AJg5xFr62ziQhmhXNp/v6+HMDFVI+saa+Fj4v1JjqMRCl0aO652HzQnhWguUOAt+
1vkNeEmhxIwXRI9cQh/QXmdc1T/KoBXzcfR6te9BAX6MZxdlqkNH6L/21Fm60p6nc4rRku7yzaH8
5XjTmqKGwirLrFldsfJDJeO/mXDOhO1WFqto/Mee/bw36qTCzb5dyeN95I5pygBxVWap0FAMxRDC
OJZoGxhj5dg89m79S9+NKxbdQDQIH5OZH2gxBSyUnQ5irtT64s7hlELZ93VcFPTJ0EU2gQIHa5iC
OncqtZwWSwQltaCVMRawQsgdWI3rT7kv73Yxy7lI6JWMaWmWjFuUWQQUJvm6pHB2ZbbOSPo4QNWe
shqIiYA/LuxwV2fY2t5yXWeLJB8pRdZG2jEyvQ1+Z5Yu2dVHMLTeX18UGohRQwpxpuwpAF/sPKNT
QZDs/m5+Lew9H+q7aiXz3RIvJbGD9AH/WZRnMZegCUbxbpbncVjFyssOKPDg+chFTRcPTIn2n+7T
1ktt3Wu7UYVEqXehiAnLv6oHtgrU8l0UCCIHWfRC9FENA16YGy6JdlRs1yiU0BBc0+A8eAk9GEq/
OS6OqOnJ8KZ5B//cenYtGodsEAau3QnLqHXRvfuGDWlU9RoMZkuDGVp3vcoyHjqYakpf8yQMUg3m
AikAWka/ER1h15/FISBsyLFpZu5uugD4UtEco26uh1nl2pv0USamw4eSFYLRAN40bUgWuM3RDnqX
aNboyIpJqJF6l3LKRQrCzKLyQpK5j5HVsD3PMKxt3EDuiE2T1CjAVvFpboA5THjjq/Ii8zQDLo+v
SSZH6Vyn2XxFk+ZqzHbcbZa/Yvru3GkN1Dfor0Za8gvEsDvurkLUTtW6c8hFoCu2Yqi5hc7w0DOD
mIvXTUykUDoISJ2+gjPcCVMr5I1KMVzpIW+TEWqFcgF2C93H3gXiAyHmQDhWjITLd5dBF/lNDNHv
7WAcYphgtGlteGJCazKihGNZgk5MsQpetlPqSldbQOdvCtpKqnmXQiRjyZb46Cg5n9PDzkpMVjUE
n/djZb/dMOSlN+htfaFk5lk+1CvtB4hKt39SBU/pA8km4L0nu+YtVcl8eG65/c5IanmP/ddZTBxx
/++5VmK1XYwAVeJd3/csP/4E91f83+vKOqc8vDfL7q4w0oPV2kBGmJ9qMVC0mJ8krJxUTbhj1VtS
k9gKNPVPRRC6dumvq10569N56E6RFa++rayYaZboGvTWMzfiYYvgw5pHI0oBwa7IZAgGWrZ2PT+3
uic3mmjfaxXns3BzzE65Ozj1aLa29OIvQ0AP6thDSYMA0PxjUXtH1hLAHMHr64ud16lwnsz6HG68
czFTLUHpw5wK0iRMyqWp/AC3Zrn7sy3GC+ON0wWTfXhih8agrnEl/2u8YypRibO/ikGgCePQ1Fcv
Btp8QWUlnfWnXr6ml6YjNDk3PaZCX+zLtI6icYd6LW6tzL2LTJogeQe/T/T4/VGSAjzvObtkvMOd
JrizTxvspdKC3p5uM9TA1dAudnstQvP8jT3V2mSdhS1giDlqMkw0jZk353+DESEBdhojXVi5FVGL
O//7H5Q2BhdGdjF1kMjRkrZ7eB1ee12xoyPTnLWajaXYgUdoMpe3zspJ2Y0nXUeqVOPIsJzwjmFV
NF2pbY5NWx7Ixz9y8/5c+f1h4vlyeyuCmeEwnd9t79TfQRXX+kqaTL4ZdoaGcz1CFfKCieG02yGb
hKFBSVj97wNt21RdBaIw90YDuMiKj9Sk80Eh337C4gEoXbTphmyKf858NbUBlfS/wQQ2Y4dmH9eO
JjE+hGSHDtlMx4K3Wid0LPtV0EdnFEPwhw5PgV0/DAi+u+kQKAWEg9Q0B1+aw6vvfiE5Mq/YW1KE
KUoJ5xBUy7+W1u8HTJJGAACsYw7JcXIyY47RwRahxmCehLCzW023E63gm/lRc/kIfHLd4VrDCvEO
DkVzmZMwyfMj2zyUY7c3fb/3JN1dadtub45r26LNtEoqvi/eopNwPtwyVl/8ybGhmIcmNJJsXPK4
3p+BsabJIOxQi/7f60iqj4ZHbMxnooiHBoxDT7MpIcp4D+wZzMBJCG26D4CM2Nyc6+CesK+yk+b3
2+S1z0zggEGDD2AHNwiFJWZeMy4mAZYziieYZ6GT8mqVcwgsuhYyoozZ0a70ZRiuDDVkb2JoksuY
eEMf3N3hwzEMCNvLcTYUZM/a4tgNNntx+pHIsYZZi8uHXv/q0PIYyn5WR/uCLy+KE0ImoIPwrOYH
EtthsPusHPpoR7v9O2OX2qsKpJ6eH8XTeoGrgRVR35zpL9HarXW9hdoWhE1XhZkqs1Zm48uNNJo8
9KfWpQc+VCOUWiaC00RigGTaamaNXYWwDN6YKpl7lskPAiqT94/Uv69tlCIbJjzPZldtSk8+7R4S
Cxrip3km7Lap5gDUHQSgBUTKuG17NlSCAly/ObSt3N3dHp6dhPxnPawMbJX1tqlaxU6gQ4r0oUCv
e7EvNapMl8jKchRPiWjbFaAY6Alw2EM4GM5DrqxXFb+f6aBrXFep+f9QPEmCayLgW3HoTmgOaENJ
OErl3JaPu1gVV9IpKNBM3fOBodYgHoB05Pn876KQqeYeqm2XPPGlOjBuENG47mTnl17J2hcNQTeC
y9GcaPPkmxwj2Cbc5qfdsHC2EZfupLCmAGO+NjLr6ohK487jXb0vPHGVAizh+5v3GTdlzeck/G/W
EZrtN/lduLg0fbF3ppbeNxDNmtf9R0V1Pex7cVPx/baBF8K+4BID00N7qc9v4+hL7WO7HDxGSAmD
8G0onkFBO0EXND3gwPLg3Se/YEct5HAxnezhfx6KDye3Jg1Er9VADakePzRwk8UJE6NC92U0a5XP
s8lcJMwRMMkx/5/mV5fv7CwGL3/hVbAOsACpvWNa2dLRH34i7DTYFiuyjnzeZoVuYnuXd6XmK2n6
Rmj8XqVneSRjOIiocaXOHqazbiyM2OGYZPFX7zoBBLZcR69SEvFQKzmICp24zh4pKeBazUZHbEf9
MPVTgbVVk2hlusonr7T7QVX2h6QDvGeqBmEnOOdzLLVsIoj5wYoqBvSIMZE3UfwcYE09L0VqQ36Y
5PxzFLoGGY1Wtyd3TGZ1nzvbTQX5VPqLBOlYqq25EWeKxhH9WLbouZAxX1G4fBHU2WA7dL17Kj8R
PW9EzbAVDevwV8eWYIR/E0W1meFCzF6C4q1cNSGB192+9hHFbsUGgf0bF8ylO9lim8RshXs+Kz/D
lXDIda5+8S0cWmEvAmlxCjLcazjjeQus8yJjrixwJSS5NoIYn7qb1FbIQPqpAZpj7UAWv5uv/7to
qvvxo/W++QIfuBxykxpOnhNgOS/Cifud5cvOrJHR/4yHcafrGGCagbqpncgfqRdA5GED7Q7onc5k
awBGMMQXUAVHSVQTbDyIyQWKsd9D0FtUDDJR6zbZf4dfuxX0Yw/ZO4SawIsxjgcqg3uA9I0NmGAC
WxSxK7yN/8Sgprq/bQVvEchS9MXkr6E+ikmSa7nB05AZD2OIdFCn5/NIbRA9lQO4risqaaj4EssI
ltBhAJj7ddWQ+LFzfGTr+dgQCi9ZL1FpErjX9bTbcpFLC09xi3bk8iyOnTe5UME1AoOusjgmkgHp
o1breoPMpWbQ3dDX8EDnz9Qim7vyNaEJj03x/u+O0Tw13WvGu7DUVX0dn3Rs0HgmbIzqZOhe1Ieo
1QvQxY2/YIRlezI11BAWjVMFWzos7sU00IESK1WBnYEHV5HocHkD7ggkI4eygEaM7y3N1hY2Y2PQ
eHWzwAv4oh0yysydiZS9gKKE1eBD8kyxnuRyY5PZCcDqWS3T4vdasval5CFf+7hae2vJHZF/kp7K
35XWdXOoVPoUtkdiOjIg2tpq2sbbYYUUda2v7hcR9En4BUCxrKxKPFYiKtJpFRseGCb2mXRl0jtn
kIeeKWnsJ8guO7nS2IMpoQgLXfNZvPzSJx5xWIqS6TainFsGq4OqRZpPP3R0Lokdwnl6zG76h/v2
sDo4Cr1/2l+9eX/sYoxX1LM+MHQcrlvxObd9Z34otlppKwIAvgCTNNH4mmqRLlnel34tScUiJTrd
gLTEVdqVEcaMqZgOi5Hrk6JtrYEIyDAJXa7rk6+X0joNy4p2PkcA0iMW2HJX+ZmG5jsQnVjt6CxO
PLFfaPhxvaoKYKgc/ZMYi+jHLrt5CnPm4DVWGo3AJ0LK25Zg2VTxplSvvunbINoZbNPJq1FyJIOz
r8kD34yYpRRr+pY8DL8rrzfPMM13bs08YYzAfPJtx1kYwDmzTon4xt33vrTace51lt/6R8fk1RoH
+gAEbENQz1DsPowdffFWJcuTjN4xfWqEzIwE3dOr3Wz1ooaSJFvMUN42Hl700wDNrCdSKLrJ+HvP
n6WAJ6gSyHyLXliPV5sIiooi1Sr4EJ3pdd2+LHkm6C79ct6AJbFyMOCXRwOMDzzyL8R8NRiHzhLN
8Ayg810H98ZA04kPDn/V82ztPuKaN/8dmfk0mWk9BrF9UNkusYIkH3aS/AMdpvvbmCw69ELXSDKs
5so25wxTqycIy4jCHQD86/7DtBXvEAcbTXywIuyvJX3T3d41D6b81H/uiThniNrrTnQ7yE6BwIWs
4pISC4IdEzsLJ9v86yDVlHdi+MW08G8zOmTUu38OADegfhtDciYNxiQNMPKKatqXviDOJQV21Xnj
dow17Oi0U0G6cjYysyl8uX5GRhIxAiEKWWEyifXcT5VFnUk3jBhSVLWWFSh5egyhIhII5fAfLnFw
QZM0s/YoiA1OTUoi3tfsP+EnuD3oVHpBVuOFG3S7hsoGBeSunNfGRCry2SMx1rFiHCx8jC5iFfV9
GvOgAHK+2jAhRmwrPDWmZD1evJM5UVzWgApTCTz/u3zjBFQg017a6I2NcX2o26g5xfxiohHDT0Pb
30Z6IX5B6uhqCrRdILX2nC3rE3CmqHNsD0DA0RmwmsRNAeL/u3VRbl56sP8xl0HOTt8rNTwJYRBm
fVL0rfMS8EGyMP6PYGuPjkZuAKHpoxgT3B0IXukL8zjPurjuB5wWccWO4dLyjWVTchCXacHeSvoK
1CKx1Df7Xf414wX/JRTSfoSaM5afGMVjiQvAIwKkg7janD58B7EXniHuLSNR13wkH2JTW+a9pw9r
xkvProf9o6V0XbpETNWz3oqXv19ZKmUciZCoFB6Qc3PPq26b6rs/DBbEwK/WU2MleR0+k5mblWMk
hoQeilhmMQcn42Nz4UXWbxJddXQX5uG9fB1lCKxPLyKc+BruUUqDAgM9R2kHobxFn58IRBDLgTTz
W789867fbqsmi1hi0/959vFve8W4OmcIIF+n6vAUDSMXhfpN4DWZ7BKVyuRa0aNwVPekodL9DF7f
uxh8BbjU0LVB1o/iXpOvhYCB/HeFQsp3Wa8JWzHJDPoqRXRzKOLHxKsrqiikubjyLlFRDIE3RGnM
2jcv5sYR+Q8T9NrJw2a4tg+1VniUe5CSUcrDsizEuVPxmXXztu6zwb8p98AJ5vnEbGHlgyq/nOY5
QdECDx5s/2om7WQZqYajg6t1rlsW89KSYus31AIoIcXUmMnzVlKZA3azg+Nr9zzy21F9chsm7Dq7
F2xY0NF5N1yNVgBsG6sbsK1zk5Wovu+PqmmJXe5AskaLJiOwtn0bOqExU2hLbXXhvzjltwxlYrQO
PSHeN7t8nUnFz6+7w+FPUvZfFFpHyGz5AiPA8R8/tDiTwyYI6bJSwhRziGL6qUwBwUgTF5Szy7MI
i+gNGFCC/e3xNUDpHFydigEx4j0E9VSMGpX2yDisp1c3y3epTxXmr374ZzlOS29wWbHVBb0wtLFw
UE0XXzTy58KnpDNyDV3rzvV0F54UbyF6DFAD8NEfim5iNPmw7GFa5GfVnoZ1Z3Ij9Pa0yOD0RY71
oE4h4DdXlTsJZrG0N0vRF4g1VYrKUNVYQZt8amP2acqfKzAGAQcXaxBMVWUmq8otGzLE+36I2Eb9
wwMdOIXDVImWWy5nHzijb31nlvzS8QV+8zKJCwR9p54HiJrSddN01VgtFVpmfcy/RLUM0QNN4V5p
HyNrpaWAxGvNN46UuS0VbnK0PXGWcgIGWvejJJC6sHsUAc/2DC3Z7h3J1g70qHbe5JT7yD9RVELr
NP9X6318gXWGFA+R2OUeXkTJLJbqKZrbOedwehRqijsh9XIjFu11he3hfg65HQaiStbA91h1pe/P
ERFwPwlApAZeAke0M6SaPr4Wwb5k3KsrZ/917xAGxJbJQmU2HWpW850vwbVa/8jTjigW/sa8uXc2
JYB2B6Hf18OIC8nLpPJTtSk0bXjS9umaCbC+6G7sIXdtMXje43jt9jqlb49YQRZbRsHZwaJJrorM
ssgkiPpHgEbXF3V7qSIqRXHxOGZWquThOGSAbJTlLEQNGudAvK2DvyCPLnNjEpdOtqgvIQZre6i+
ot/eROWYe4avD4k8hjKuSbQQ6qzala40ZTFnBHRqc5dBKiv146yZsNrzp/fQXrOkm0spPi3G8CcZ
Cuqn4SXucw/qLf4rmGKEwl1Xgi35tVEipjc9pNffqcWgDiWhkErDH2oyP+m6NEtXTKt3YcZBS/2C
vUP7hWJzhnd1T1wpTBHWojHofflZSvLlc/6yIP933OEiYRdgOMfB+t4LcQi/abJiMjmhcdSOaafg
oapcam10RtbouITbRpft7/kB3NxjSMXAGokRgbPmLm17Ci5Zs2yaZFg1f7iyGpKuoQSuUy6db7Z/
NqLgEkor9WWZzrSQ/1diimqdty+EFZF+pJpjJYdJTmVUGZq2w5zeJaCe3jiD1BsPmrfEQ94LxrTc
YtcR/TZEm/FkbnybR/WHLlfVyKDI27weyOmCMunpgmh5GyU4P0FBN2w3U8GlwNOJKQxTQxIAT/8x
Ok82IyDvNBjsIinN5vtIH8zQxd6/lY9jFqjaq1LjEJy58KxcxB0+AffWpH/aCBuxUH1zyayHFpaz
bU/6BpW0VeKYMgJfcu2JY747pjrnR5vYqIokTT06Efv4rHRSfjZV7ogof9vroBbTF55krFUq1eu0
kIR0dOnS4ca07gHg19j8GnQ0hABQQDI0/DdHUlOq1zwc4a5xCKGRI5rwDs2XxqerBFQ74P/xTEOF
TB5dlGyESK8TDljI6kLikXiZcp4Z6UQVdC+HmPPjO9huh+YMSGfe4Mo1Pj2svbluMB2OfGQwjuk5
ua6HKjVFDyEHeQR88BwiWrp96Tjy6SZa+7gMHOv+yGAqV7B3+9nQ0dg9TN/XJqxo7/oT123zLxTI
H4kTjckRtnPUHMpAT1S5NnBZNDv52Hr85UudGenpuYa6HxM/dBe4ttwntOS/hq/5lnd4CcpO7VD8
7bNS6ZC6Bbh5I/2Lj1scV7m661WiThCBsL82MYjVx/qG8P47wnGiS6JRFLzLkiXE0n/9rJgd07B7
MC4k8YqyP4jl/CLKg2Y9qPhUplDXmIJ6fEsMhp6v9hMSTjVfzxdPFiVbRpsRXnB6kO75I/k3KU3Y
1JE/9lowUUg1r2Fnxph6hjJUhHKN0tuTze/yohNVSee4UW8Cv7IEkeLGpPl59JChaAgx0DqA6OtK
bnHbdhPgnTmmLRR7eJpUIMLM63q7JaLTrDA/3WKC3ZN9oz6nAwQwdvLCSN1eDofMfuRD2wmjElcx
6zlgp5tHdKWLW/y2cqV8/8gbEuLb7HN5lpkrL7CBFi050ZGcDxWfg1tmYGob1X51NNTFKjzUsFNi
uR5w8t9cCmdQmrtw5kL3Lzwj1mxQaEhlx+RnYnP8Y/ppjTpPuXkSKXzh76YRzl1rG14QK/IgvHwu
XJ19uKZmvMSgKyiEypuBIOjQnFLL/PyqEQGenpJFR3BUkjSlOWdeOseoVrlLp8hqGjm5jPwOxd/D
CNnSGJ48Uaibs42zlLTahUFWyoiHGkX4T5FbxBIK8l9dgnY5xUEh8t/SdgQuGnAszeu7DIh81KAO
6OwMUuDkKzW/tNaA8yM/CaV0e4kG5C63zH98fMtgaeOvCjPF51C8qhZBEp/DCYaqEinmC6xmFGmr
k1704s5+Xz/VWfn9VUIOCCb9HkrpdETvzD/1qLtibdCuxQkWXntpz/fau8tDBsyeQhUFEDNgMBjS
K1FlORibbrSR9EO1oDAsjakZ2V0oK6EKcaV1Dw3qNin10+GLwxUES1tLa6DumI6duKqoQp07riKX
JOjTzF7qDGoyA21YE3qGn07gGT3EpRRUm8KZkgfvp401f4hpN2Z3OPvC/o/FFkow/ijnVSH3SBze
ff0qORXaSRB88AI1JheGGuFP9Zk1Iq1G73nkdfZUOP/jvgUO8eujSQwZ9xU+nWZrJFUvZjA6BahK
GHKw0DLDUgWIaQlfDFbefGlFH93e/pfvCCtDq0BwtxSNQEwnQjDLStiEUK9cRoa969BxAcC0lqaQ
7HqnaeVxJdoMMkOeAmByNq4hyI0c+glzlqiFa0/iwfWCBsF/VmoJYDF8afLV/E9qEJUrrTlXFt5B
S50EZKHcx/eoVArBFZa7Kr57HZqS5tj/k9wq1Fof6Fml2LDnOW/RoVgHd7jv000a1uZV4OzqAq6Y
53uK79qBL55HkkmFJij5A6fCglO6J9lQsIGAC7XUSWhT67Kb5XGRMBhFX3swY8S2mVdCWCRb57bL
yTPmJ7b1lsn/I04Gxo5uxd1vcyJqZSA4m68++sPlnnpB6A8ucbvYl1W+qi35YzqjK+WQ95CUidDD
RaAlIMWXrijPGkhPFOzESZgPwvMoRWlgHO0k9g1V4JbWbGTQFK7Ng3TuAHWEnkC8CSDlsscocJWu
OJokuv7pAE1cLGWqT4jQYy8Z1RkY9lwHdTuTMhei4q9jU5LNygL2BE+/bXsaKU9kT8sFMS7hzNPG
MrPk+rdsPEToBzFLSVjGhMdVwkSWodI4hAsn2micInL7nEJbPkhziRq3cEV7HMaNUsua2bnxTTJg
/2il/VLi0BAuMqzlYPI811xcnROku7VIV3pDqxcf6O5JvcfpJSx94gA7uCGo9DJWnu1/Ge6NYln4
WuNDZ2Tzr/52sK9Zj0tjyiFcAA+/8HSBAAmysc/ZFHjv8huWpUboPt4NVzf5g8tzByAh/F4C8oqv
3ROXebYYV+bejThCPP/VbvnQCl3UbYAjiH9S/zvIwVN7w8PkRAQ0xPqn0f7X6wXxrp5t6NLPlc9g
UFt6JU2R5UU4fkXSpTsSwpE3ffoHcRZFkjFKCXFPPPlFU0mx9D0kpgNxcmWH2OnXWF13KeFbgagN
6KT+8wx80EdrkSQnmuhRlHSLQ7pvj4Vuz1/fcoPpV11b0Mk1qLiW18MReB2f03e5th8l35pI8rxl
U+z9L4yy4quYsfxCWdV1Ei46gk95r9DPkdjCc/ewpXrOcWl4hW/3XrNlI/vqxMB3XoeIp4W7p7bk
2eLMqpDLfRj9Jj14R4fDFZjLsXMC2IGjLnGB2k7eCr5DvW3iX66PNVNN2M+IyMsyAB6jkFIAsnEJ
jIcvN24myHTWH2E0hOUC3iddMs1UiLxIfQtUaylnJHbFh/OKcEoG6MEWwCrKMZ1wS0t0owQ0MPp9
1YEgdhldW8xE755llC1azuztknDXoN8eBrEE6KIBOzDK6gHwD6TPfB3VOhnoncPXgperEc2Q+H0/
ELyC4yDNihVK9YIQqkFRYML8tSNUlTjaXNDpj+4FV5ELnpA6HQMRP1nHy5GuCmRigQHWi7tYCV/f
qybkQP/QqRoO0A1khCU9Vk28c8xJprvI329TCDAvwlhdsbv3fPXDaLFyc5Y6CKNDuAhjk9Dsm5K8
GGQtRLUBbvm1/ky3lN8/w6d5qhr/1My972PwXtnV84Q05Atfxt4JTRBTv131V22/aD6A7wISpzCu
25LzAf9bk8qxADMal7D1omojNHNa4SDWNyaO/SiWklKc6sN6r8GQrPowjZgT4oyH9eNMSd3dkVX9
s8Pq6yClfcbau6zAFHuUMUBM9h8672vA81CTyA78UR329XqPa5t71KPXZaMg951bUr2o01/4qq00
gq6Y4O0W1G2IQRwb4axQR6TBUb6ojnIQcx5cQphophjmPpF3Dl3LZ1CUGRrhFJf34+CWUwT58mjM
YMhIRKuYdbheDVb5iziPYioBBI1MUndeqc187juJfU4Is3DQfu1bgTPPR+igfPZmtI7k+kh8j0O+
xzuGGpDEzDJeeEAhPfjEvvAKs7pRmAXKCIaxB+2Eph6yZAr1SXrPKyyNVshqsHdZrQ0yppW1hHmk
+MnpYxehGp4r0qyWFbhjlU8bhrGakuygCMwopczHm9aWERqgi1PrN0f1c7DAdLK/XRuvtiNE+YFB
Lc905IZpKy1jLqU6Cazn+eInszpWcezBDoKZhnQ0UL9H5sat1K40tWzJYnlxWkKRg8fBk8Fxcjfd
EqTFDoYkfXJDwSVyDMbrIFHXI/q4hrdhHumPK+EAZ+cQvRYd6FUsZ9mhu8We4cz9KflgAQY8MWKC
fg+cIjXVgUr0vRoHLbgQPQPZo41A7QgMcH/C3FKwoBXzNH/v/3U28Qi/RsJP9MXAFyXi61GElNOp
TX7LlzGbdO4DlxcVEax9hdcmSq35QqX+5ahxO00dfWZzvTbu+dXtwO2YboWaGFVOpBQrNmwLAdr9
74dsC5L/SAnTkBMD9YeqVwDchGS3tDtbuFEQzetWDPU5D01pogDhTxb84Ie464jF6Mp7S5P5Oy5q
Y+ZGaW5XDAOvK1C7sWvjle1qLz0tfkhlZJyOK6BcDQ9ATbCxvXK7vARVBmpfUVZzWWiscV4JyvQX
MydcTcVcfnVT6A56Fm7sGIF3/F4Wx2cI8cREIbIjW3AKL6gcjl1WRguyykejYyWqud16ze6nHd/Y
r10nXIQME461ITNC6U7yiQrTM927v3TdELQJMO9KZ9Xq6FHRvj01LguDxZbsfuELWQro4duk/N4k
OOLzrwAntLLi3J9mvTM3W+C4wdDQxv5nP/ODi6/CkJA3b2nbZaOJCF2RciEsfjimbkElmPPnYaRg
9WmTlIbVChJhPNGJ89Jpt3ImAnnwbERPFpBJH8pY9cpXGega1RE7hDEXDtK6iOtAgkzOTt9J01Wc
rIl8yNZl0nANbUt6peqIdNYsD2EBcT/ylXqA1MBpDE3NDnURpjE2X25cq3Vk7UTZDjGBud6si7ar
LDkroNE5885m7F7MRqxOmL5sqjbeC6vgXVP6FUvVJPKAlBHg+EFE0ZCB4d6rtoS+mSZ8zd1ShbTL
PLtdm7cake7WOZcFvwr+zlC1W1zdfPX7kpoWhGEosglcP02hdpdkDAwbn/kboCSKVC4ukWAQu/tW
hu9iCssT5DepmPqTYlhmlvBEBtBjY2CWbfJ0VBO5T1+ha6meHmYmxDCOpRvMuPVPT0rkzgyhpKvW
LWoqzigEK4eNdcxHkUaMCYMI4FLN4Q3KaDASuOJPEX8sNZ6qg9g0cypnRW49FWS8HZLNysTS1b+G
athkzGVHuM8b04CS9+Z6UZjvWtYEu2LDpY//X5pt7HtXaV9ZMflWIDnHaaK2R0vV/R3Hnhznz2VT
09hxPG+e5dCyBwphq2dQve86oofOmbH8X1++Y4vXvsXKqgzEoCHTK9nyq9ZKUNmxRzmiKqOcUiFU
ZpnY8+OjR44LYbkwhDAbP9V5tINlG3AQ8FKmN7LVUT+EaJySUq2hq1QePravDhuexnKgeP0OiBTX
+7TKuF6EHw0UOC4WEOc6sOwHg5lZWAcEVJkygeVJNTQdK3k2lqCLo3GA+pm+BzKadtC6X1FRCu/A
DROJ/XfxNemfR1I8CrqsHM9e5VueOX0suO7cebAwmTHMIBRAX6MC92Pjqcous/mJ2lDoqwFbUrCX
euiriXptLqvhYVVzcISqWE4R8u6Q6KDwMFzxvoondJTLjzmrPqC4v7NzP9cP4QzZ0A6iAwvSZPhP
S4XFs639UZHqsc2ccWADMYUuziBEp+ZzkYeQSqjiCBzgw1V2gCHH2sxDJ4v/ZQRn0DhHZjfapa2K
haauRUsN3NOsUIICP0QScQQ3qRuT4SznszySnTj5SwUcBK60VZXloRP4QobuVTJbOARuEnNp/otu
6XiXzCb6aQKNWOZeAJwrUfK2Njk21+A6S4sZsgeihHkenxNCv23Pvbyns9hfdy5upx+qHHK58yqJ
zi2iO5kBUi5c/OqUZqxF/RSSV/NzJaxHRNX1m+Yb9+C/RHB4/z0cFroWBZ35yh9b7JTu46wsYPnb
62aaLdSpBtOFnMx4IMrsh7XvqRS3zkWEXoLjn3Jq/JV7ax4I2Sgu9mhbjBA+bopBealoy+eyzsgg
Hrtg3LraaLn61VNAXBylMCbYTyAc/yhQpwvpQrblRxe8hfSfJm+pQMce9s31JJgvms4ZZ47gSBQA
j51rrWtKJb9okpZbverb95geWfxnH/NpkZ2HqfjXP4N9LVPVpSjiOFxIaRCN+LhQthNUsf/4tqC/
MFmOKD4gjLxv+tswrFa6yCN/EbkFLjdo9uGKNYr69iQGN8/FGu1M6LBY1auYpwAxzD/4rkeQxPy7
oDwFno6La44Qz3bBCDfBak4hbihgwtmMuJp1t2XmIOiK9i5Eqo0IZI8rRhYEWAJfFsk+iDHmUNtF
X+kJIu4e0ouGQwEky4oM6Nher5HNChmt42V0fEEl9BFzOvP/ghwYfCocjVrWVToSv3K7lQdWLQJH
PMvnDL7we2+88JMRRQ0NDJXO7QRGjpJKUzEzTfdW4GOlBUCpWgdG6hr/T0QFolF1m8g090KolsHS
oARtqZ/y69THnCUl2i73NrcUBvlJ3nqc3cdt0RjW+X9GmIPBpcEIj6f7G7JTcl1Hx5HqusDKiQCm
nSnPFEuOPRJRMkNivhE0dAkSwEG59Qjxr1YTnogFuMxEI8O2U7RIXi6o7LFoZqvfxqTO/vC0OKrV
HjkzGYGqmlD9QVnixlPMj5r9Jq4StY9zRXvmEbN75LmpmvKeEgUwQQ9e2IMiY04lFKXdU/mAXlhJ
t9160SMOAJQD/TgRP6EfcTSeZCRY0HqwoNZLaOnD+K9XUhyAndnSRGIecXPIic/7Kob+fccoN6km
OabM21lnsYfOm/GwD9lb1h4m27IACeHkXVOVbk9o6MfElEDwfVnb9gFKl5atSAtcg/6hD/JFkLW9
LdzI1s7xIV6BvXx3i7nCaakwvMiPzqjsSZRLDIC3s+Xt7DbfkORE1LdJaDZf81VINc5ZaLN+XfwF
RfimLUZDhK4MhGxc4JfipV5oEKQAhAarpzJ++1UKOSdcBomzzRgpHwbdHnG3zABHHbI2jfH9VC2i
4d8ggxyzJRes5BZitt0pC7he30TIE0hL35ybwRUShJkmL9+Mw5Z0k2tqY/SoZce5VaPw8F/P+inq
XkwuCc2IIIb32FXTDVFwC8q1ie08Xv2ZwxZPH58KoEqpmWudHvNF344W+8X+Uz3bqjnhSr/SsBhH
meHxSvvUGYJ9cOaVcox64clV40xtXBwgw/Io5BBNBk2vaHh/zJUwdjK4Mz2pVz1BcrQo42oU8aXn
3rXdMgIiHu8/UjkxjEz08Ht5QCOs9QYFWR++2elmxMQnZsTOUZbP3iebnqBZlBGDsDvT4NT6PTW7
5n8wvg9HH3jcB/9x7zUmOzmlyluAUoYxYtf71UHVIcDnE8OlMOJEfBl5kBNRakThHNyG6GgKLGss
scPICmp42nXeV46Ix1CrLG2cezuje7krk5OEgo5noVEBEGYAPjrcZo7Y5ins7EiIbBxk71IIPMgc
TSlYm/xRVWI6hcd/cl2ZGCsGLfNiUKszOz9v8L6JoGjhcvQxZ7KXe2bWSjNJ6kFUBqGPDgap7t70
+KCiXeEU1p0Or39MQxLPXMILwsWE6bphsnkovp4RFlc7XvhCx6aBHlcK/qBmBEWlsLreIZvmFgTu
LOoVHH0sWF9jL4fbopM/SDWC83+tSkJUeNUUtv/SDl+7AINbxVSWjEXS9WqCwckDuvj99xZ9B+qm
NZtIf0eCuguVX+sO2wUcVma3d/auTZ7dw62IOp3j8TqMkUzKP5TahjzgSszT05KDQg0pZ5DlRihY
bj7wtPB+pcdK1ibXWiGsqzJ8YaMeD1WhG/WHYbxnJJn5QZnpXXbJAcprMWH1WuTANt1lngT0vyHW
t33e8NwkzDH37CZq4f22rTKddnzlB35kCPSVa7L//GhZxw4RKSdHdz5cL9YJiDB6kLXzhdghdv5h
xx6OSNS8xstnZ5KhpaH5qScJc7wAHNny99XsZcLzGm1KSmLIlyw40PViODh7KsJaLY/NCBPaAFmj
NK8SeAuiDKC4ZLwqLnfWpu/Mb3ic9jplpxWlgLHKvvn7mbL2D955O9iKUhc1Mi97Jfk6OW0GtOhM
5XvESDvrD6K3RDpNa1LOP7ZQ3rvlBP5zdUxIpVj5cAf/Od3neEM4QoHP2qEPAZXnbp88wIbnotOv
S/Hi1w7SAZkk7FSZy6GojiOuJr56HZ8k/5oakZUgDUS8GMc0av8IAMq4gV7stO/K4Wyh+m0SRaQe
6zZBF5dQQ3GFQWq1z2uJrzNEoKYCvkr3ab3tgwQo+YLha81TNty9QGxeJYkuXCyJ1g7lvmM7tzIK
P6XdR5qaJKM05IVMI879jPgfZ30Yot+2BJwJLaa2FLQLwLsOLyQGH73CykVLRj/g8ALQIf3qvnrI
1ymmN1aIUkGmMvZIx0R8wl56RB/jEONxg9s8BQtvfl8ZaTrjoC6RbBAjicBouy9qV/r5P1PDIn4t
uHfKKSjsrjdvkvrHdNEh5WVDJabYm2fdyzAzQkJ/NCB8s6U8HMH7ANdWpvqPzgcdquXfxcefIyFE
p+EVEf61KcN1bXaM0688LvgPM2JP2eQtmKa6k/IrtdpxwnQh8MgH+XN2sZ9JFsSw7UVXGm+PeYq8
g0Hc9BVEVv19O46l28Et0tRViD33iBD60XvZWQIBkjMIaDmU59Ej3KANvRn2+t89YUHLT70jZtWx
aBX0D/dids2AC5/KAMJoTGMZEiqm0au7WQuE/e4lk7Tf7CqqtXpn9yk2Ahi0nHtzPFUgc1WKSNdc
WwUZt5KabO+7S5hOfMN49ofNsJxe0YrDK19mlLWni4x/4kfeeERMOAPK3z1fPIZOranHDRG88Diz
frCb2JMNms7X+WIoKTkQos+3tjHA1SEOG8tJqJ1D4IP6rLzb3sPWPkqZ05qqfJQGz4WMa79PhX7I
LOcOfAMS5mlLj7LJ2xSd+S+gebel6i9D/X2SD7ERF0CJbadgluEMJMnho+o6fs4ZF1e2sjdgoTmJ
qwtkT8MBPKorFxfYVxZLKdAi63F4K8GugK93skmSghJ48Y3utMnDyH47enPi2LDc4nqcwrFBtKU2
3BGGxVxKitgEeRhu+zrmrB1Sq4Uaa0J3vm1pG4HYL6UxtZWpduDsWU33GMPHkKN74+rIevVRHhWt
eAYNh2id67qBARPuvkdTvL0eg/+dpRR3Vn41DML3XygVU8Q7bEqIBFj1JW0Sy3u/hSGkaa36BNP4
3OgDt56KX+N3ENI2d401Vm6XhGRImrCrj4aUscWedBbuAqrgd24MePmlZLZm5KCM8FmHLdJ/E73F
tFb+JNZk5uCwPF2WzKVFiuZwH5VXIL9LNuOfjf4lzcztDEi+BUiwNJrU5tJFqOexw4sf4OujKHH6
9pncvVJ+MaiAP+9oF2EPIikk8VLTYZ398kiy9i+QTUusl9NNEoISHqEeZO0kh0JiUnNAtETxHNeG
ZxyuJ3DhBcp/AUmJBabdPQ/zd5UZqo4AyEXRcNhEY/2y06uyXmKW0cfmPVICBEhDDLu2+N68xVxI
v+ECXqEg70gLLlu5KIfkBpMXaLgGOlpPYTgkeHnwkdOKVqyZ4hwtAFiNnVteFB4WltBIpUXqZWnE
0DaP1OGkJNhBfvGOuotyoJeczTszpWzXl6s0NRqhU54KtaikBcNmjwIBSJPsacRzCFHWp9TdsqNd
ILfW/8clPgT6YlyV6Eo/ZrHdP5Cd8yqQlONYR8AikElDeb2lin7gDbheGmfSbd2SlnWPC27O+mXe
G+RWkQHX7OSvSpHDObSBe/rBqTd+SxezAE2fftd/I1rZARC2AlHGXvtjHcHeCEvHFZL5iYenKg6O
WSb3xu/gEJnCoRS96pGJUDkKLqVKe7eC7XN15utuY1NICmCSNa/XGeqFylDdEf411jNU0Z51Nx0d
tiJN6ZlnEuZvuxujVrYqo7BkN6ydqQzwzuw5fa5gCUyfiXux0jjp3aZCzdrVKxKprs9bQHEUshs8
GRXyP9946pWDfImsX+xMBETY/G9Vevea244T8iytVoMylDFIxnLxfEFCI3tQMS2usbqM6tUpdwwJ
DxeDw2A4C8ClGXHwocf6d57pbKw5AeWF4nI47gkd1N2opX1VZ4g/NCk8l+nYeRlKbXoQ60XZnU1L
lCMY8s3aClgwaS30CsKp4RTvCD3CIxXFA6mtNyma1012MW2sJ7OXjBi6fteZwtE4i0H9EK6l8dOR
9dF6GwMJJxxj9dVk28//ifJPs1OTf3PQYO0GJAEmXitHehW2XgqUPjWYkwQkd28E9FSXDi6gqsaR
hjQwiA+fFmBCEEAV66wJCR3hVS8TIwUWVp/CeLo2EKPIUr84ZSYtRUsqRvZKcP4MbZx40aJr9n3c
6lkW2Q1YL2Kc+jeEUt5twtiMnqaWvLZYH1Fr/FZEgxnQwwzsxBhZEqV3+YKc8Fj6lMGdABmjyDwf
V7eqXbIf1YheT91U5JYFfNUuG5ZZaNBTxSEUof2xToDVeNcXYXP4BWZ78a+4rETDWP4rpHfnNm7G
qpjFwoENOKkPhOYJ8Tq2iKM1QqHzaH1mGF7llQLAKU2x6Yt0XJ/jiRR9viBQy9mLVtZTPhpypwjj
ByQxyu0cYMfn7cHra1Kfqmu0MBHdomEtsDVxYluUl4IwFGZ3KDH5r+31GWK8sAODRpn/AIbcsZWO
Sm5Q7M6BFvU6Ctew6EqLF/6YnZBEvbkdBx11+XMJm8x6e4LKhqoMzaV5ergTHYngckDDK61KQMQX
NnAqKjzNrZItHJcXraOm/XKTAiy0nsdqwhm0oqBP6Qgi+3a4skRfT8llGrg09xCM30PJTyvrIT1j
jtUPD/LeCKXkkwFgRvOhUUTJq2W/cAHHrVxazCfrutlFdCbzek1jq26VChP0ZNdjxBfwBrE8cA2S
Dmbf1UXUDJnOAe505uA6wz7FlzzFV6gjujCQRuAUAvkUHeVVBEETBS9dZdniEnuRAWkwnDXRxCr5
zOrzRiBvNQBWxJ+dA0aKqZj5NczJEmJytTBy9OLJh41KRSwID7vIQA/y4ppX7eajssuJwugKZJ7n
jRXKMg0mXlc4NBykGx9wkwR0CyL8wFF3DP/EAW64JZNGq62klyRVzz4BxCdwXwolsVIAsVMndRZP
QODocjfw/gSkb3diYgdXcU9vh/+P0xxItzcHHwq7Pdhj00WWk3WVqxpXHR77p7pn/5LJ3f4msL0Z
KesP1rdXQE7Z86bjuw/F2I9zKblXc/FJA3Ybww/JSYMSCRYwfIB7PL0lXbtR1nHI7thCE0HKs+MJ
vtVf2VvrGdgIQVba7PXg0C11Iy8Dd7Sxy0ePBA141+dsCTaqXKJOxlSA/b1RDhmQ0VPmzrHTFBT4
Ep5KD+SdzzK0rD1mof2fh2UQEQJfctPjQ2OBR5sQIK0HaSqaXm2gzGw8vzJpiFaQg1ujK3+a5qIP
MOPQnFw78D+u8ipW1hrI8CdJK3sXOkX83I6YUtioF6NBHWSf5OZizfPR4mWm4AQtmwT2fiM6Av8Z
HYBsj05qWajuUIxQS3pwDMgkDAdYKUdtRyGJOoi6AJ5PN6x5mUHXrgY5H+yd2KYKxZFHf6omPskl
B66HWBa1XHovzd1r4c9T7fTjZQLCr3QtEY1JobuwlcDLGCcl0Yt6DdjkbP7iIrPLuhwSQtjFzjfi
PrJ/dMzC9Up4ssoROpvUuFMRUwcwu9VfUXmIcUDoYhkjk8kAHu+tHUfLAyOSP2aEkhcLSx71jim9
WYLdDqfvPauELJb8zI8vbzQs2yVkwGMbStZaxhFwvwSOeIi2akxeE7Q55FociVmJvjWrzspFeYXT
V1vMdLOApHoiashLdZvjYljqYPn51C6mWufWdxZMot8V3D+/OhonOW2H9L8PfhmDQ1NohdkFP78j
rp1dN5VJB1OOHQwfVtAmiv3fJPIP2eb9F/Y6XPFN39cRkKVXMEOk/stT4eVFeKBn6UiW+FTLVGWY
rtdL9AsySELVJWOS2d4PJCSYoIDOM5gNtbgdC41G+9feVTYvSSM3JowwZOqjfW0cO1KHbu2j819M
Lb5k/yAhLaE3ndg2ojVFv1Ch5PjnnvJOVTECFFa7w5NYtXe73OY5MFjZbWc64YPBJ83Ukm9BG5le
znHG/C68KBRCLassIpf9wpYdUlymk4nTXjsdTqn7jwz8TmCzV5KiP0sVVHSXsQqpM58bRtqYphiq
zdcaUejfFJPv9yDmek0KKotrZ3upJYB+vxAcnFLkJlDgP/toCxk5fIbHKuXbn41GITPS7t7sBdEg
3bJHtN5aaKD/N/mt9QcIgWnhrsMuWuq1pocAMOkVzZiXfZlArJBTs8PBvXWLDvctdU0hFt7bJlWs
fE2+/SDQk4gg9WVtrKcXzPYKXe/mk76wY4GGzseW18jrnu9OjjM/qS/p2qzVukhDKfmirZuGHaS8
BE0u/8+bjNxqhPzhGa4r/h1Yg3gZ3qlt3OM5FO+GeRF7CqGG59VL/z//g+5OlVknwt7BLxrVbVXU
/Ojn9NjnDPMqQ2jsP10vf06P7hQX33f5vmApZzKaQ3gFwXNzf5ZVrssAEXjhToBs9Y8aUM9ZwO9q
8MRbpsbbT2+gICD6VUxBQCOcRareyeq46A8JGegvir107AjqBRYDsYYmCmkIcYk3V83IBwB5V+HD
XsAgPaaJKPB8bdBcB9uvwZnssJJfZfIYeCCUDu840sevEAMCRcEg5B1M7K6TIfbi1lpp9jRCCYvA
FzR+FOJh5jOv59PhUI+dpC8pKc8lx85i3jIvEx5bEfszRTN6GOMizB9dhkR2skPN5PvYO8uHF7xD
Usja5Y+oCqPYvOvYQiLJL0a6laTj7QvB32F1btGrV9UdwIsYBdfVvSFIec5ryZd2VQrG1hgd0vn+
AXXT3aqCfedZIbaKL3IyRs3cNSCOUQN+I32RGhB7V3AvDmqME7gtDWvWh4Q5nG9hjZ3tvQNjEOa/
p2BqdxmRkk7+86aDuUSxK4zg/mG4FLrXbDf8IB13WOlhwgtKpEt2H+5k1K5jDfRf+aCl6L+B70fp
Mg+HNJUC139BIYHhHJbTUrWk3QGZzinl37ubP+CiciqJ+LjAq6PMh4dYaQ55wbV2evgVyFOw3INo
mjrb8qLwNTQgFKgOwhIRFjxdkxaM+8WOKybytqj0kkoU+iXTSEbztRNw16FTWi/Fdfy2gqVacea2
8aKs//RLJolSN4+BD1Cz8YL9iTXYpiypac9R1UV45jqKNS1LrlqLEmWxBF0QHInt+j/vMpDuUGbx
0V373/rih7K1pZp2IpDAMmYm5fd83r5/ctNi5p+QGfYabcBRhP2qxOLECK9LCmmHRCJLjU/J+jvO
JfpdP6C+RROR8CRax/ba4ZjrI/P5oluw0vxNjmDPj2zraMkUckbX23E1/Ads2BF7RaHJOgbQWgp7
Xk5TnL+yW1PDfcLrwZLh1ucbjGJAQg1VXRlakWB7kCI13BNn8wJDlywhWx+ofhSOSSpBOvLKkJ6S
fN5L4n7i67+iwyULI1ikf5R7jsPXtwhkNEor9vYmLKHgqjA4hzMh1iWwPsLTYUFBpcd4YnXvCgQ/
ZtyHhDqavMrDKjq+G1OiHMQOxUq2O0rFoMKUDnjTjHABllXW+0Eiy2BLX36kF2KIuxciqwPi5NYb
TwEmozEh0fSFwEURlbjVG0RjDtZ4ru7FSJa1JSopxH/07rkaTUlsdIgRtkKmEnfWQOFzm1BnxVi2
OOa0N5X/1oOHc9pItV5XCgDPbNenMbbNnAm6cRMjW3sMm5blpV4YZtC3zQxOz9KM0xEdQI8MhWcz
1887fhg/ZBXa4GHWmqAJx4vurG96xvl4TP1xVaha3xX3HXXvdD/KpBCcheTXIYyiUlYhUy0SIP3J
/tBuMJWjUaWZF5UueynjVTRHQx3qpH4T8aCZQeVpohXJwUPXSQBt5NoxbZhFL2fw5eAxLKRtKLTk
kUpq/5U5DCJiWqpU7AUjXIy3y+BJxqCH9a9esF1ReqZJ3cfbCsIsv5JJBbCY0il22SYWBCCuHW2o
gqY43hcil9dcMk4VJ/cywcX0Kq21tSNBAgn7JVVqGHuTMpflCjgx93uo1RQmLQv1pgAMTMrMFd5R
LlUopro2pm59oeEb/astlGQamJODoark2Sbs2E/c+quOmGnfUPyrIBBxtbvBdQQM6q5fH2Y7XtXE
NF3vLJrw88HDA7fs3PHeZKvDFdxLHsCB4xDAhf4sakZZcUhX0EDoDr26VJtFqqy00BUp1t+FP5f+
aSMP2yaSFlec1ex0THhwmQhg3NgCLW/G2F5+BmmpajAtK1sn6cTzYMhBrR/pGb9mI7qYGTbpUlH5
gpyb+goZaiszPVmxM2Zpeknd9kP3/95vOQPq4kJiFyDwsdArj4CjGWFlfZlNjBWmZvFNFL8z1aZQ
p+t3bKKhcaFj/RTgZIe4aZ8mXvwYbINJEJ98NCoF0GAMiYQ0M3ew48x8ViuubhiSceQxNP7NCfju
iCqv66CIwD4QvOwJzZhc6BXufSnOiiCJpwJuIajzaMA3GotV1QWX7nZE3ge5ZUF9Xk1ZKaRcrNns
aiMKLjW/sdu4TGF/zjz27qkbD3HuZKPKtbdF191cmm2vR3DWikmdg9XYsqv7GDHCtx7NZ3YxrSeM
nQFr3Czpp9qgH5cx/bT0O7N8BBEC1CnorFY1bQtJL/StAWdUc2uXUKjE4O9/QiTyehvpPskH6W9b
nZB4qtrbqhVGdh9KK73lQWefn8XGXRssIZwxwYDvpt7Qi2GaXCi+MOJzLFy5An3eEsLEqDUBvqzj
3XnqUqOCdlOHqArByL0yV5JQKzMw6fyK+tlWelznX9BnfAyAyjXDALLOexTFQn6FFXZpYbo8WXjX
hR55CppDC+alxuuUZehoF36H4jxtz4tOnWQQyb5Elh+ywGlkRD5vUxB0UUeFZtRtC5hJy7NB9cBK
6NlEQoLE4BhsDcu79DF3mL81Ow80QtLZpvCjCJqdXkkJbSzwyzxrl/Ez3o24jas1d7aoVskXjRDz
Uv1yrS+6dV5w+nnx0Z/S9g89s2B2Vwv2q5IXxlGkdjixypKQeZnijQNBlEEM/Opg+E0E4zyZfVq6
aHfmG5KI0KellCgX1G9ZC2y5XNY+2QfMBLmx56eNIVep/h1Eh3es6szzeEQTfwrHh/+u8LpfyLGY
3erdlgmcMSvjn58kyBoZFlYoxTFqPDV0LuSGCxfkP4GqJtWJKM6x9WEQ8sHJtKQUdxmnA94nGLW+
jxdVVnVYZhgfo2WaR1PHHvisQFAA/YR6kZoO1KEziOac21c7So2LZPj0BJKdcXffM1Pzveqg+KNz
cZrraFpiOxmKBWp5ho5D/mg7odttQwHUfbmPFurh0gUR1y+LC9bXz8AHnjJKm3bZuWY2Iujzj0sE
a8XTQgeTBvHrfdyRThVRyLmc/jcyusjvgW/7RWBfO06n8uVZQpcdd1XyLAZqPeme/7IlnB90xix7
1bD0d17p5wj/mLYx6lNzsTED39A85LydTvRRZjRQUi6DHxlYc0FRPgS+GiXBQBnrLOYo0lvcgo+g
9PevKSWfNGusvh9SxCgxiW8PrQC7eYvwIXRuFxQM+RpCmsIBR+1tE5Ua/7PV4k3vESQOHJhwDI/B
6u1wl7jPR3pkqwvzVZLOLLdLwINpMaPw4Sfg9vrp9hp73I3kFq7qCaNqXrX7nZGNdlgSOyRg738d
Q/Ny74Z4fMwbsGTkzcfo33xR3+M9/bzRJYYRzkQe4N6UWWTcVkMgMBfH5uhkOng6g0s+OsEo8W+i
XqRra1pnQRejfIzMbcKiYrsclnnZGWXfJAv9NrbWfvbjTysTblc4x7vgsEhKpVY1n0bc+mizjnO+
lrOmKc/TpsYK6SMVSKfKgKGCcV23ll2O93Kfy/5NO5Yp9arbuxrZjl4rq+oxgZRfMQkZ618i4oXo
DZDtwe2baDnAELb4KEyH3H5ZnZIM9nuOQ91A/NP2DmSqRvTcfYvgOJ7eow9XDd/+zakeItpW3vlu
twJi5poU3Z0XMOg9J/6d8ZwvB2VCWDj3JMG96Z7bKOV/C60Yb3eaxDt4RrGhzn66qzRof6jYxgc/
hsDLiibTcZJEKzvuXGgb3lLW7nmBcF9R3+RYsAfv8Q7TQOEKmSs7jV382vQWL8C088YRNPB2Rx7u
94Q5Zpv7x9KY7I95s9EnDTxuaD6RaQdRUjO0u9/dTLiSAfoUbMITAH4NGcJU6J4A8tvhtKrdXM0q
y8YpcWW+l/aaerc78jFa/WmlkEXKYMIfB29orzf0a3Im9/uQhz35N4VwevtuTbBvR8KxTvcYicKN
LZgrcvZd5P7czhkAaUhWgT0yHcoXPbUfhxWHokqWongFc68lVpvX55+wBqaDSZDJ8qKhajq0BqKO
jjUXHc7fJ/wpMYzs65dHDPqTzdIwYyyR6xuCExRnY0v+KaDA6lI8DDn45k/KTg/bJ9la2GR2LAdr
21NyXfcTxT3BLZoutwwqym+wHvgAkLlP478N0VeB4usvs8PjA4cvscDY7n+BtnP1p2QiMONotfxS
qsH/ae9W/L9QIEvPQj2p6ly1cqTcKRnlCa9gp4yTjhFbH9iAUWvGgF2JCEWvK6AhMPdpwAwnEtsy
FxAnDbCLFB0/jFVs6GHMZ9jzcS9hKFM5tzEOo/Ck9gLSJO2ZbR/cZX0pnqLOOXgHnI5TEhYORqe7
Cp5xW7Wgkqr/0muJnQTiekjCjcamhOcPtmGX0nuom8ZbKutN26eHQpBp8gRnBH/jfGcLXXCC9L4R
6XyX36ru28Rlo6zDyV5795DWQEI091x/JgsK4GuBY6m3piSU0dwvQ9XiYKwGYj+N4JSTu8kmS8eu
wUZSounZmW8o6+hYoyFhM2kXH2sHhX2GUw1U1ax7b3siODYe6s5tbgQAMRpjtMdjoY1KZyuvAH9k
c2JooiwdAe780sa/SUJ6MlzcqUy6GNPqfkho66QH7iAfiOB3pH5PmdGLFjhBlO26KNZnhumYHLuZ
ecp1KtDLFDCJY2fXIDcNQ4SFUTiy/KJIxF/bP5njyi4/kgVHJT/cw+VIX94Wm8XBUZFkG5wGJv7t
ab53TkX8UGH7XyyKenibRzrIyZ2QWhb3OnsJJOakQ46oPLTz79ZLWwEE+y21YTMy/fjy1VcWZaHK
Fnb2+TGJzAcN1bdyYk4RdgiwumIVStc7uZ/P/S8eguV+WbWglzU3ullM0MA2ra2jPmzITrg+FUQ2
n5pkLTNxXenUAKylwjO2Rm1KnCeVBQIJJkpLMuNMVitZ44Y8qkgEv9qObCdhX1qreODlDyVC5LcN
LgxzWmkQIfR/a4zqhBYb3QgSfp0y0a/k6XDvX0s3qOYyaPHnoBqBqbBeHkaTdI0MzpMAU6AhnvjM
0e5hrWIpNlg0C8c37DsDibG7a90YfbvmXu75GZAWc/aba6cVAFnNmyfkV2FE0St0vI/otg0vG8b6
X5UZNDW1LXTzs6Pdolnl7VfJgfxxLU1Gx1vGYRfC30eoc8zAZ//AKsz9euvggn93oB829oaGyyFE
ee9miDEwUYrihjmbTX10q+o+2BHj8qkp19jydfI8mBs8RaM88Gu8V4pPV6wG9Q99n1931Wjhdrwc
mlT0EUErf1yd6WHqTfDyA1k0dxNetklrTGCdBRQDUynfsbApmPjHT1QCmaI73UOMreNnGZUsQfPX
hpgwEwTm7YNowxYHruaBwebrgqhyNvlBPoDbPo+ftIuWuLcTlgFXFsj3Y756ISXTYdgtWFFcPBLm
jnUj207P/SMLmz7js/mpcKRPDVf1j5VfpXTcZxzuBiFOvg4RrkuU/zxmVEvQvn1fVHAuDFXJJQv3
3a2dbsWYz87UmuCpip9tQYPwwauv8K9Bt+RNA8mnDet4BEkNKd9FhDKHBUqCGqHVmCXkpuXrXcQl
p/EX0aUyQY/ZqruawWVvzC+MVTJRmaalgkajqxxM/BGQQjrXNU7q8YCWGHTlyuFUqobyXnJsQwdR
AcdNc+ufb+yMyDhx3kaVYvJVXUQwnXOMzxcDMeG7l4BWwp2kbTOwIa0qA0i/V5N7cBsYNpZV/YV1
PvSsgGXdy5fYiyBUfz1RS/gftcWwC3mMjE5z5+poSyAzmFWlFn2/wC1JzyrgncIV6iu6105ApGqE
rfHzj0wGS4/WrupTh0PFZ2cvuJHJ6mVMFFcJn2s/ocRrwIyn5NfP2aG1s7m+YlL0KOjV/vz3R1SZ
9Fx+XEgSl++FNmCvLh7tHC8ZQEyOiqm9oWnU5HhmsVpjw94roHknC5yNjFbfNP2mBpAIM/Lyn/fh
7aOdNYihzxtSFlqVhUFRfsOq/mLnKmlVXHNWFYavMyLXOM0qSDd/7F1w+UmhXevFPsxeioYU6nMY
0VIshnmgSJUpsUyqOXNs/GKpOxHl8fM4rE4WLUDNE89G35ZWm53chfb/ifoNhAExmJBAVg4+aMO6
/npTVLg5j0tZ0ui/8nI8WOcUe2pfKN5neviQ5DltrXWQB6QxiusV7aAws31ZeP/3sgRzEgbxOUpW
szGxSixNKWLFvVC+ahvYSxmDkiZHW0BjrJ7wsho1qxsC2nJgqfEjT1jlOo9lb6LLkvfxNLonvvvZ
UiQz27kUS7xhUqEypE9Ghk5hpVYHAF2eJTUF8Q6bigNLcKQGEIG7dI0CGU7/0b7rAm7d1gaFNNCX
oCX97PimIwKnGdGg4cKKyrxIYWPLIesExAJcs8DH4nGCvh2EcuLMyJm4diIZtagK5bZIJIODOGQd
TNEncAMSzag5DxTnX4qiby93m4S0T6u67YoRLyJ0kQmd62ybDoSFCmRtG2c6k/8q0aAFIxAnBEkN
QPTwJwipfPEmoTM0qTx0yncvvMDkWY8LTslfPeosJTiXO8hsh3P3E2YoK0H1ULHtcheT5W/ycnVD
IZdHpS+jhHAgYFRGjf3nshC1OzWLn6i0a6PGK/hEIZHPZTTvvCwYZmK+vx5Rvi1eZ+HwldoCM4J6
ITKDizUmAH+fIbv1rXJ2P3pjtjlm+ywFSOmMH7FTaz4cua+AWXCJP5ARfQowOWVJrBb83PEbGTPU
Khzzj8WRhJT0FsVe5e66KqiicAymakKipORwwTfoDYlNZYzLxWWZ+smJuQZ62FB5yCudmvlIzbsT
o2VLdoRfSh4HEKum35cDHftwLcYYsBBrzaAuNKJ2TPOzsc5ftNJi2R5fy8Bvk8ftTZTTwJry3A7P
c5OwGg0tAfZymBufyr4RKVoMhFHZUzk1ke8tMpdjFsIyIlZ07zcRUhdfjTKehTJyrBHiaaVlEkh3
IXVjT2lWAApW4jZOPny1d1xqt1iWVw99Ida8X/E/3DQDaucgEgNvPUn2ZTLjU9x09o0EX5JBAd39
GEgj+Qr72Sn6FLpjmc6FDpelsZ+oLHmYsLZge+Adaq/aZgvibegPNWCJ3XwY8Rj9uXUfFSxM86PF
NEB1YlOKt4R1HCSaZpjOoGY3EcrqGGEhtOwiDHKcBjBWleTRIuJUX+8Cd6ClzecvDbgiuvpWL4TE
oBlVWwX+mMCUh5OVPvUw+A8u8O0Y8rlVbQk1vTWKuoCBr/YZBKWzb8prxr7QaJbvJu4UtM9CkA5K
gsNmegVgF8uEaLUSwFTLxqL4K4LjH6kRQd0F3xuh8aPO99xmJHjRYB2cxsFZqRyYIJrVoSCuT5B0
orEnyN+DugVvxtkaWZgHF80i5e893mZiBLrfLZ6ZznbN4yu8kVHsI5OrnmHz/CvnIV1k+X7n8yss
xKRxMz5TiLg+JzS0naaoqtlxvAAu2GOQ3MYqJsa3jwZ4oRCoUgb0uFclp+YdNGJBlJzUXwAnwNkn
1b1ogFTpxD04IHHlJWJoEjtgjxdqT+Xfv/jGHOLV9ILf8zU5nrquTejx/IsLXZ5h1Y9c1otd4EPs
jfkqBBeLvQeTCk0+NHbKr23AzMMedX45GEz49R+Jm0GPI09xgHz4dT49W0ae81oPAvVX/m5SldNt
UNEA8Az4HuX4DWL2CQzEBWesGe/ff3fjc/Hy41G5XdFgXHnlBIboLAVV1MwlD36aCTyamjow6jCv
wmUc3hcX5jQZt+XocPcyw/uWfR552SbIGj2j9er7XMrnvHJX1VGZtSyID+a9AqZ2Mi3rHd3OxPyF
nquktuGXTvnaAuAAn90a/DemdULGSY/wOJegWAqToSa1Hd707s9t4jKfYI4hve6TnkFkNCqq9w0Z
zGdju325ny0RWgVWc6jaV7VRsj9q3kDtVywmPT/sDdYuo8eOQzp/h4N6MAC5LooZU+7pF1zBovuL
O9AT8AVU1xi/T0HSGL7rQlEGNfy0I/QgkgJKUidA5aY37Th+mo3IMi0sAHmxKzOYur1XYmXYX95u
hYsQdTV2j+TzPf2p+muzcgcYqr44mQasdsoLkoAN9g7e7bwBJHcinMhYI6XWfdNITyNy3YSETpZ1
z6AQ6rPwLEbCMiRd8cg0pXjg/AMb4CMQWI47zNhox9pJnqoEUpsYmC9SIDSJwj3hmevQFD5kAzWI
l/Rzq10Zjiwcv+5DhCZaHiKydG82K+HbPs9p6DAFT9nmvPl3M23ytkIOqI0ugLFGy74Uar5JovKX
hZGctP5GfhF68qfBo4lwMwNIp2UNKpHBXN/6ZazLxqRcEz+nzKJschLCVrc02BTJO6K5doaeJOz0
D0pvEhiCAmbvfIV8gFSxQs84imQBXMmwCpEXdJP/DffjIVVhzHJw5DRc2o3NDjIxpLONwMIspGDY
CAY6bte748iYtZ9xGPFcSasfXjEDNRfFj7MW23iAH1BqjTQhul2+Pi36vtHBkutZmri4+Y7CUynC
5XM6IzAtQ7xuCCrdE9PikyGh5Pa4pw01vfLWFMKG2miu3yqxe9o0V2OEkAKWHbDZ5nq9bnUGOjRa
WbQ7bzEcrn4IMGx5TxpPPyj6Nv+PGiDXcwV5JGiPBZuynPGQO56HcNKtfaVc/ZgRQWpyFzcsuBJf
zFXYO64Anm08YzcNTmlIj0fi8otP9Fd/irr7Y04pV9hutnjDG0bj++71hOLJExlOIpnu98mKX/KC
CRMOI6csvrwuQUoTVBxiYDI955cmOqdt6X5MlF5OituJiLQTkQiymM+kYEiJ7jGqAF+lt4w0ZLre
34RIBDfaxVCDusoPiKFpCGaytTOAElrBl4RmiNxulG9tRkUFmOHXiNIrUlbK0FStwEmL1J6xJBtp
gruk6NYV6GC9i/FFzgK2oGcW3w3n3Nkq57KaeEm5x1ZtB+7GLdVcFbZl2VT0mQXLek6fP9KiYSoZ
GI+9EwCsfArahwX8mUWRGRzZZ+/f5uBh9bP/33nzhbX/6O49tqKTYHXQiYqHNap5d903fEjxSvXd
LgriYeiiCzvC21Pmx8Uq6aKRAj3omSIb2y5kevcLhw6G5RSJHEBGVJJbH0+AgYeN+YPgY5+mERph
FWi4dyYB1TghdNk1I5191MMIUOO9CHXlYORux2JG8BY3Z6XevqZzY0GuNtD0NMqqj5Dm5ydKVNT0
V6c9idsuC6eB3/QK94o4bKEM7O/a+yNpgc7hoLPRZC2y2P7oO/RGO4DBwuDljdcplTl6FwgYkLDU
s3AdttVRQ/dNei+iFR/GUPsj//M5YdDLZYdPyb6QaPpIC4hQ6NXK8E+WVlBlRqsxZ54gT/lY1wiU
mHqvdrg2YyV3Hcr1sXf3zfty9b2+nBfudAokZ0PD0C30tAlYDLZtKxvHSd1D/E1i0GVvhggfyM/u
ysNJe+/JQ7OhTnz6VvaUAeHyIGpGTx25SkfkDJLli1iZ3kSrFKIH3nXHsbOyafAydvkPkMO6Mfpu
XbYWuBMMzqyuvbwMEUlxp7mszy2OJqHLkpE4lZFSx4Ay1dAv3G9pzHxUdgFJBDGlJyp5JeegkBRQ
0+xjYHe2NaX3n401eqT7YuX6ex5X/JOhNt2oVQ5EG117VeKFDxjjgWoGvuZfNWkFxr6umvLu3utz
MAzmK30bbv1nJD9X8pfLj8YJL3PfpVlFt8sRf2FFcLLQomRrO3zl8wuEQgeqI07uVa4OMDqlZgix
yRqHOwVdZ7CsCD1Rl4Okc5cVS5Z+CeFGtUo/oXG5MAxnoEVh5g+Z2eHJJ/mZQnoJJ5/4SYNSZWN9
ux8+ZIPadUQFanwJlq/M1So6VLD7FI3k3Idjl2r8mOWWKlDRqr8B4iHOimrJyPmatjgUucjd2ARl
tam9Y62YlcttSgomhppsGj/9jZAM7ik0X2otMnWoU0QIgrEDpbTr8mMv9hg9NxX0k1NejrJUqSa9
b8txdia+MykDXdTj+XlEYnS9ATswr9j6wWl2qcWu/4WXsu7oHgjqRLbtxBrzYQgbJDPhQnuUANoS
yZy2IsdyxPKZfm7bNPRlIdjj8GTbj4vLyLOMgYEHmNNzY2vhzasNMYdojps/qPguChhw7u0EDEzc
RsYpQnDM6wsoopBZntDt/TKMLxB/73ZbMKJ9OVK15E3dlsHxrCQxaO0uQNHC1bVWDdRSJGsgcSqx
+QMZWOf+F6OIJoAek3muJI+q8QEZTE7/lstnKXky3TacM2ezgfYoYJ4j5VcONOOcavmbRdJPDA5C
KzfhBw6JO4HlfQZwotcEbcT7vq1XBZxdIBVo8DeI2RsfdLjQBkYDAMsMU39sipZwu4h+v0891z0i
8WUOb3lBiVjpesr7L/dWuZuQkluLadw+ScA/6QeGym1vv3dDnj7u51ovkZ5Lt5g9TLg1TW1HQkZx
DXdpJG4FKUYyS8o1PgenkAZ5ZlipEaaqeAlsVQEhu23PLGKdl30IvsuNQciRZjn2YwdO4q0e+2vg
koIamALahGhPsIaBU18W54ucdPJZrWyP5GsidQZF6NSCvsGhMQwMpw1n8oHaTcWi9h0vq3v46wy1
xuNNu1EwVETz8r/HzffdKt2EVbpTELGu0T4qjgtcMtc4wTrnXHJ14I4W/WFySS/Th9O1ARHL9gn3
YTXmr0HzZ+qmHlzGEjEqi9k6+WEhPXr21D4IXub3Qlg/xOJfvZVUG/QlO25YhRTfQjYXNqEgKzaQ
vFZPJcavZaxKD6k61FBmxQGtkL820M1yEPUh7cdM4oYEsWLarvIS/+baZO63Pc4iQjM8wqm/7Y08
/c83EhI5JmO+7smw9yIePJTDUNLopD2t3YdDF3mTo/fvbXsz64dx1qnBsqCOPSaK5tOiAX1yK4dK
MHbi1a96x1gXcqdG+lU6q1iDtwGrmUoA5lQJmoliHX+uWS+jClr10lhYP3Sx9xwFqm5vc3xe3Uc7
YRf2g4MgutAhdCWTyxSICdWwg7QUmHjqszvZGhgamztPdzgH+B634sCwNziUWeTmdP5C4Trj75J/
B9ghz9A1NXfgMjbHumS2soMhr0IkuLiyLf8p7pE2Cc6+XK19cnmb8C/4J4XZg1nyTVvEwVQ1xsAY
ee75xhbPs+nhSO134c4zoY/yo7vrVGDUFU0IyPHTBr/Yl5TOZhH9SG4KhTDIe7VDM4bopm+yuqgS
1u17+8V4eLwABt9UQRkN9f/zljI7oMT+9mxJjXTEjOVXpf+nSG5LSimNhBOcbFOSUVsy/mDXuyv+
1hy9yBc5Xuw7kQJDAfw8x6c0BF5fr17tMCHGBMsPkY63xzKSBAn1BQA2c77pBKQfD0FHbF63YhlJ
PD+ditRbN4e5o5Ey2Lhyh9WkdOLYkXd9JkVUbxCXwDuxoRVO506smWU4a9LUUCjq2FfTzFyAq85q
bb4SFWqjDLNpFIB9Iu9E+JjanXpGO0J9UBf2Twt8lQ0qjW2mIMOy1sjivqIrKFSV9ExsuhYGrQrp
YNh5dh9zQEI+v+kpYdRH6XWuYDTJaVsh/1Nc1j66regUDRqWr29H0jf3sYs7hGFI3PpZgStSDLWh
jj3v9yzWlk5bh5YFN9oeE6Jy5KGlhONs6QpigTnKrkWjAFPJSlTRvsc6VX19gEOvhG7M39tMtS+q
7gQ1qEWgSks8d/0Bd/8JSGNJy2MRfMRwPYAwJwcB8TqnYWou/HrhinUO/BuYoBjohQgLCaFLgINc
dKcvj318TI835R3qW/OI1ZTAid8dUIGDUWpIIFE6Gi+6V8tgIOABQMq56kwgNON9sWxtAx1gH3tN
NtLTUOiOV/ZDvNwrf1zLT1X3O56VAT6g6QuauBF4cKK3/pyY6uqxl/Udq2NdYU9YeC/uwp9cj8W0
FNfJRV9tJ3zY15BaXB96HJ4PbwHVBDJvoTJZRI/xRH7iQ2b+3GOYn8EEeT5SqAOOZyBuQMMCj3Rb
AtNkU2WqxjS1EpXYkSFwqT+HTO5SoJEAT9WK9o/SbNS4HiEIlVL68wfbj4nSE/VbouYoBdnzdDpR
PjpDRh2+gC7dph+K0/JfywnS9JDO1X6BF78oV8yLvME48BAT100aaBoTWyL339s+cJJWEocIoyLG
eXTvTK4vtkq6tOhnbTVTf3w8L3WMpv1avgxSuNIJ10oYZsJA56+DvsQn0pCx4f6WU8HGvMdVDNaS
PTL+VtUVAC9EbxhgkAZvKAG0JoTrzlbpMtn4hlMGTmFSVanwUHegZ5+LEnWW2Q20qiva8DeaqULx
e+7fl/BAkQjtlEbfY6lzVO84oxg2TTPtX774XymLCI60uZjn7e33Nnsfj7B4FSNfTK9NVHyKIDr5
LZ/uD7lHtk6By5OkQ98VHDNlAHKEXhVDKj6Rr2w0l5P75++FwZOwtmAd/11XjE3DePtuib3gD82L
HPAmdpHyFqxp2SEv28d/D/kU2+eWTzmEyzLnQM/8jQVEkf5BhGXQpo1MiSB9XZnRfAT7WnvkKRXE
zGr3Js4q7PJmbQwEI1G4CD6Vc8W+husYcw6jHYDF7htJR7KZC1Si2DsPBIF6tsZGjN/6MjYYhBxw
Ty85kPVGW9+wfQCvUq1yMHnISjrBhSefJgyeE3oayiQa2jqfKfqJECL4Q70AW8a+lsajmZ+hQwL7
1fm/PhpWRZvQFVFLhvHKIK1Qjcmftcr4F3dtUTf2Z5X1+3+KhuZYkkHIgeHn5FvQ+NAwCTysa4Hu
KusjYUSItRi6RnyPo8txO+ejcQdyGMvsJWn1qd4qcGy+AJLYsklT2vz7qHo4WHQ9+fshD4q2UgZS
H5D3P56soFiCMQga+D29mJi7jxK47eIcPaVllClvAsBonvhU/8bujRhovV0SgSmzHrE+cyf8Oc17
B4G5wxmAom94sKakPNPobHcF9hIC0MjwSF3ioZO0BIAjCgS5DtxmSzlaQPU6NsmtM8bmSQlAapyX
oMREws6uLPV3tZNGQ3kbbbk45uh0e3clbtLJOD9zMmyrTezcvXpmAcpKQ7lf5NUtKxJB/iyY4PCt
eYAIzS3PMsL5Wrr3zwqozAXaNIh1cz3IpejerMFfiuA44mrlg5/D82Y5CKY8yTH5LP68zPgIvtvc
T5X4kjwetLw42YmeX0fA9DlNHFkC3BRQe8YYmnSGW8iiV3f8VmCgJsf5jkftlzn/XyWkDgfdX5QX
UJXwGWfkqfb9oL6QCW7ObxaSS09hn9fEOkyXYO0N/nXoN31SAGkRIPszvpqYtst32bR1U0af0BXr
LUZ4ZcBUdK+W0hvlY/QcHh//yn9B3OSMismaHa26edOZcvr76ttk4kFChcUxo3wgt1Zl08DRJPkP
oXlbO9JpBPYbHZYhI8eWW3BmYCI6Y27FYqhfVyrEUThPqGhJmaa8kEIgSzyqiGkZOxIK+eDFxl9R
oe+XkFvSDoTZH8RO60glwt53Cn1P3XUv4UaGRt8NpcGA94J3lVmyvoau4qpPOW9donxhb3PBH52g
UAAlh8AW0/wyRbhYrR61Jkcw8UEDR/wsoTm85FG/0wZsNke03fYktkFrDyeTaND70zb6QKeXne1F
FcJxto+RfcFTiSHR6VF5LkV8rQRNO/WAE1mMN4aC4WdKJupewongqvLqEMkbBRr+9oMEmf6eZeel
1sWfBUPurBI/yMw6OtwWf3slMmncCcp2KuMtzdJ9BQUx2rD9y4EEBP1Mc1WByDp11Wy/JUFK73hY
MxitUynFPmOtG97VP9vpQfLWl50Q5VxQ8tzx8b1LbmawolSLUFRdT+lAdNMxZadb2YCsV6Z+DkjR
a8WJkLsI+g8iXtUi+fVe7kPZmBSTFxKxVO4i8xaKu7XBdyM1suSiCxZoMEq1zdXSh1S4ulNL56cc
tphEy7IvILmorJOjZ6c9DvGQH2SEiGdIL4yxN8rUZYLBM4GSxLf6ECXQdfZVJAe34pReqDwsZkdK
xZrBPZwuUJmIio8gv6LEqq1kYaAViS9u3G/ogRkyJJgedJGivvN0gSwr+TOGOcw7lU2ohYpo74Yb
4fmAY/WPiI0GN3EPGyG9Jxs5Q+pKGQyr0PDqqcc1f64dprVqMo4I6IJkf9adSbNjclMtq0fN8BQ1
9W/EmFrMNTqbwegHCOYrXSDv8ClglX9c+dIN6pyYYWZgSXZ1XsJs+D1SWsgVCoNjY69ij3C7lErI
hRbLREI0dcC01zMQQ46XO+2fAsg9mHry1PdMwqpgu6Wb/AJcGoz88DbViAk1oDb/IGU5oGaoEdhF
r3GyTw1HW5hVqvpuzBorgI3Hqa9PSeZ9jqVN7Vu2Av8PIsf9ez4WJde9PLHsuzMLREumSNspwMAP
RHgsbcP6CeNCd09ZlVuYyOBXPJBoz8OF1ugu4eb4Aa3mxt9jtVKog1MT0Y1CjBMvKToiA+BUknVq
i9FcP/pgh7B8b0aNmcyUraIXWmiQWiA7Ezf04LCAqas9hIyB/2R5DVjzaGUKWN2PYEHROK3oLaWG
96eP5ZeopSZ5OfNOaNUhul36VfGm5oDLr3TSCbXb9lRdNgxul3RnmWpysxlBof5kVrGW5pzPmWXZ
gOEjlrVguTLj6eFp93cM9f8SGOkgr7V5lZZVMgPHVzPjnQ6MECnp3DweByy43sFup5vbmzPIrv6/
b98bGFyEtCq3jDu88yvlSyLvxf6QTzyz00ULg7CWmMWBVlTCI/0+NXdnkCI8w9I6bUA9ZiXsiqq5
7kC6mS7xVWrRpbLe2zLlvXUMyVi1wwVvaXj77yfXikFHCwd6EakjCcx+EGYvNk2SqhpYZ56BTvRn
d3dyFm4H/+CzKmBCOaDGjJ7HDqbVJWUNVFSbieYfNIjFzPTAQaOury3md9r19CPrFxQtM3Jz1+PU
Ui3/7jawOnTv5z4g+OobAleVFrekkyNsmuiZNLC+gHaYTqahb8gCV7U5qTtBs5tAR+u/tPxsbHci
vJGZGEOfabM7Lu5PFKkW0ybJEFgs/Mdn20kAvbzn5lmRwKrQ5TkCDjlmyX3sS3LVbknPZTolm4b+
4QJt2NBDe4efUZq6msMXtM6kFjp/kOBWv0fwccFO0dRTRPFtXAi0Q810sKTwWZpPM+kdItwHaQXc
B36bB3iWIWZOTOkCxoAWlt1KGVh47mUc9tf9qS9IayDoJOC9myHnDEHUYWiXJ4DfRqtkM67mxcid
pEAG063BrrNmXmH26nO1GXKbr3l2yxIWHPQoExQBDN0qwjgbduK7ZEQY/+UCGCHsyxz331okttDD
4boQkTwa1YmsCQGgZsvtRJiGUSlXIDNqJgxwfSLl5hjHJM0WeSdAI5e1VohnpPI7EwGQPMcrJfSQ
EuhdgoqQHttu7h5oXyPiHBsDkdDIqu+9TBPxThuRLs4JoIh5NOAO5nnrqVGv4BGq1rYedw9meVUV
hnr3k9DDmWMEr4H1l4UlC49NYd1WN6StOJDTGD6pl3hnMoldKKxygi7YH3teDaz4R3N/XmfmcEHW
k2MUkQJ1dxA7pMVOHxzD1TsW3ReNFIEXukiU69eCZ7LP7pjkduJHCZPbrzttzsq9q8ohQo7EP1TR
bemGj0rucxDcl4JD5z6GHjB0ABvYPCsEw1eKpaEx639jvATbVajwu+J/iUKseLCmz0TnI7VZz+Q7
VP4vFn+FTbrdCjnCsfVa+rM2R5/zoBu2rLl6gFuTidoD2r+oEQFPwTZnv13zv+0EN3E6/82YQs6V
7LX7ypqdYW8w+hMQl5tz8HykjODtmIlyPqF3903lalgdmKTmHV7Tm4YAwkLeEeoy9+D+7UIbIkMT
eRkhQKOGcCUfbEHQUzFGN+BPztNdLGIDyEsQ0Ty427jkI2d2ceQyOmtsATVnLPFt/SjuaPs961BL
3F6ZuBEj/JZJUWEfTGFTVJ0LbIBuVTAazfCdpn6T9Mf0v4HFKCE5FWSjtH5nptSjyUqPxBC2xYtk
Mq3ZFNAYecZA4aG/likpMqkJ305aWBDl9thuEciM0Wjf9f2kmWbzTv7lq5g3MIvlGXDdQJKIlRTf
IbrWIOL+o5h+bgXlyNabvkNy4QKtJDzLni5f260Ll0/Ky+QAiwyJ5UyFf4xMHvn8is0ZMd4El2of
jdaZk9c/au1e850+SfgXSBBJGPk1UlwlafFDWHZRLLy/9Q0C2v4cQh7V+d3kYLtUTGR988+VqanA
KaxFXIiJImfuh7vXukGjhJCiM2V3fNJFtzbFuBz8a3okHN0GFGL7QspoYy0uhHq/N0Jx/q33NsSr
D2JoDy2Tm/D1mlnGE4veii5sjhb4oT3GxTsRFh4gjT0uBfFMzRgUuEUwyzzcKqLHM9Ud6s/1ptEo
b9X/aiFSCgHJQnrheRc5xRIpN1hmvHBkU2DT74T7Id9auGOEIUsUR8aT3b4hQ0kGJEOKoZbtwCY0
JXqhZFgXTidScxZ6M/i+nBhWYfu20n5/m7uglbGsfsN1u5yJQJR4CMag+dmIdzbcxLRbBZ3xc+oj
860A8hSsvxE49NBqraKmNjPo/Lsh53vPUVCO+zbnxifQFqIZMxyEHLOjyW4mW8nO++qffd+pY1Va
6SO7rsytpdpqfQ/ny8edNO9D47w16h94NDg7FZ1Ah0zCmEvgYlyS5SiMmFCOQffQywyj96yuQVJm
Dkp1Kdq6+lmw0jHy8c+F4K2WRtwFcwSc2G9kG9izW3mu32XDJf6N5oLW1Uyn6ot/odcTRs2EI83k
clNUJunnv5bS9d9zhf5rtl5OWmvoQZ1bW33DitFRmMbjhGTYyapZi+D7o0wDeGckWcLRKXI121Mt
+BftRP2RQbPoksHOwk9QT0ZqWAFoJQbD3dGPY9Vl5yFQaNEKaAaaI4LXSjh3RKF7ww0zq9nLtikX
iJFe6Z5A3H/IqMSYx1iYHsMhTzxhn+g4qX+DejUMo0qOlNqknQXKmF/m624FVWeJ+2ZKsrfAr0Gg
uh3TSEOQeidO2aSQoEGvrM9RXgacX9jyBHI6w5G+ju2FSYifdmBL9vomCTYMD+LIhH7erfHfQKC0
KMpTvlUYbdDAKORhlwSv+ziNQstKC2cWypYJQe6ErJU++Q5wD7K+mZqbDuuX6OsYMr6pkR3ZgGJN
t9XlXjP5TiXuDyAdFqvskPUMTUZA15zvGQ8MeNPRaMuwMLgMWFJz88HDkYbDQn9OQL2nKXHvKvH3
M98WAJR+WH370iQrWZrJ40Fspcevc1TLFAA/yRBXm7YkLoy9vOhZkWKrHLOvFGbI3WbrDZfwzOJf
P7ZoVnfbp6dn+D6bM6oof5hjxKGsVsk9jmmo2za3u34b3FZlik9SIgP7BbauQ0/vFciWE2HPskum
CUUNs5MsW7+Bn24dzTAppLn9maJIcdPzkJx1KAbLUKQdCfaPIodaTf3nJEdOqJ0X6qMBixf3y+L/
CJs0XRnfETkt5JavFuyWln+tAs7VBylp9vjxZNgVsCyzWI2YveOohvLb1m9dzhymc5IiZoenHHyk
VK3nfTBQiC4OqXhmbG6kv375KYjAq58bva+mInczFcrsYWVYA/TQbPrr3pe111KJon0uej8CNPCm
Do/Dyh/WpEyGV29zndg9WYAwiaUX7N50vQPtGsWbfSp2z6IkJFZ832ZcHBi6r8GuWyfIjl9EaU2x
57WDWYhArizOAqubM/rVVxUQNKiTVI66iMDoHrPDbBTA6dnGnIgK25IQNrCw9wQ2Vy2mrU3y31rg
d27L2mdBJZw0G8J69qUIvlwsttmumFeinCNdxK4hgx8Ul07EcodwSd4ZW1Wqao67TMbd6jpRwit7
zZKLhFMZI/AxBMrpuSgWtTNzfnPMuvXKiLrE+qYjJ2ZTWJBBX18DnoCNXNOia70SWUW1l0KVO3fz
5CrtiVrI6Mjh1IMP4VgGTLrUeMES0vfJMMITwQkeFNuPUYquPOs7JXf9jryZsYmIwKyH0pEdbDoY
S19xLCjPDwk1Zcr/zSIZ/M8qpePE4kRdvymzJvCHAcAt/4Wd/Ne7b1ig3Y/WrvjF2aFQsJGWA/2t
bS+AoxufxP4N/6bApMG/8PWnw1sYOR6POaXROT03wD6MgeC0o0AjoZ5a+DiyybORJwmtabDge7Z+
/8Cqz+40V+2TZm9Dle8jbdDz/MObBcc9A+8EEA46p2ySTE5Ep7SWTjV6xJFJvs2r4EsVd+IxY11J
7L6tzZVpVd8FaYjBtSCOgZBO4PhljLAzfL3wwjmUS0ic/uhdasLEU7o5297QQTyDtyXIB534lCvq
mOjmlPSe2iOg8aEAjO2y/DfmAhSdNGl4gbOcthaPM1x+GERzTXuGvQsIgmWGhEt9/M6o4x4/YfOE
zZibZmI2vXbtwUU+s43OUyybLEXt8cwXXlx1mxQFib7BpT+Yuw4Gf870CBr3SQX2+Ljr6BW8rwNN
5XxoPVN4lydJ0Oo0Qc5n5BeDxW4+9wEQA18Xg4HUpoU6oz9c1WAlXHpj38ZceX/wlpe9CePQn/Tv
dijk0nZyt8HTvl/KHephiLFC68qPK6X5Jbyo+EpNEk+unABaNAXixAOCNTdG9IHptpOJy9jhrSAk
YnkYVNfWiBNBrSwp8qEI0Jwx2tNw98nMzfE/QBgrBBx8bHG6SH7XausYw88BL+2SCbtwfOM6vBrG
Qkectdf6JxyGToo5/mWXZNptf3mznKjhVkUzDNJHvBrtOPktdNJopLqt9DYmyjjHJ9vceBYf4a+D
wmf966GBfy5fwEJs2He7OOk+HaKgqRXKth567nw9NsSgl4GpAu4EoUJdThzca+F0/nh/NFNcRCwX
eQMQZYt15yirr5N1PQlkhpgofP6N302PA0Uph+U1TX8Yzp7RTznO/MC0VmGO9yM/yPF8ijSqv1GM
4JC1r/1csjzeaqDdmtssn6Sk9szH7z6km8RwjgBHzpLMmjCG+0bKjkfTZllTmClnuQtBunwE9YGa
1XvB5uBPYP8ZtVS3RFZBGt7VhFHUdp+87pNvG4Ra5xU4baczYKl2qMIMbo3UvI5ssVVlFAcXwjL7
pwD0bwgwJHJvKU0QwZ9JQ7BV7e2A8yZDpQ2WB59LYXAIFX9XTnCV4Qa+rGjHm/51brreQR8z3AAW
c04CiiKvkXmvoneejMw91y93vKjr1CyhQgGlUJ+cet/9uZ3061WnI5bS3AKvVkIyLqcxohBfER+L
1Iy8T4CMZMfNfLtJXk7/BsZcwtjpPwYQTAnLFSDzSjRrS8qB+KJZiwpg7Al74DTdQiBLuEzFOjS/
HCg2i1ArGUqP63BCMTDhkU785uEK7MwpiqjPdvVYt7pHUKYRoLk11JFD+EplfL1e57CnGN01C2UT
9K9664oLz9rUleITccSgc+7Y1j4lJS6Du+BTLNE1+Nw7jL4Imf1aTy+IaW8bsJKVeGaOeeuJdZ3K
tLl7N9eR1fqkU8ADLqy2bQb2YTQHwI6ne/wzFTO8PQCK473HWHMhST/7K00uLjwPrfXVcnpPv5nE
LBjNMt2DGRPNT9lAtYl2ZuHXxUk1GRiBe8Pj1uFdyNa7HsIqoaRqpH+I6WPmUgdF1exJeSj1bMbA
y9eebjXFwhOv1rYadSWMVhiOvVnzR8XCyxUrhuUB7UKM8aUyyMfypnlCYFwNJ1OxR/7AuJOtZP17
errZchj1hi86723aX5JzO1egrVjXTiR5GvLLqzpvLotqanLSvdeKe1mNoT/mC++MiCHuapG4rEfP
kK3HIBswxcX4Rm5Sn6GLndu1yPWSKoF+dhmUnuJEGik/XYL1xtmHnMtV/beV3aalmEqW9H+ATb+M
RY6ZWG9WTaizh6KGKAhdsl6BLmhbBEDIFFZEmtNox6r8mNPMknwGQSJHJj313uoYTn+A74Czh94g
NpAh2uN+PVFQZTzltZAgDL2cxw3W6m6V/o5AAZ6+N1bwFacTj79xf9mJUKGM6VdSnEGmHGEwcq8i
a8Qoghx6cx/5hm9bW19n6A531mA5DWOHQ86wN41+NRGMyoaDpwq7TL07SZfGdaDLrRHXFJdOQEos
fykovW+3+TusGB9cxaakxF4Ce4wmFOhXgEAh6JofLcZQRWZBT3TbxN09EPsB8m5gVSWazfkboA3G
FA68p/N8YONEKIKD1634jxXCu/PmLEZTXWQ9nF65kkE7Nf4FENUFbpUOV72DFpFr/VfnGIqwePeJ
RP0hzNZRHjXGb6Ld0AFoFwWzr7R+Bli9YZJjLKORAuZiDeQD9kHPQdFFm5lgr77ow5M2Do4leJuG
+bSn80fNMFIKoF3AFplLnvqeSMvF8hY7g6tMpbPFMjiffH/augz58XZO+aeYDTw/YJgurN7ZNmFz
+H0XuUCwvt1ZSWRZVDsbMjTq2Z4JPGsPUlybU9z6Rh4+t7JYv4w2t63jfvBt37Qrd10WiYBTe3rG
+luclixx/vQx5QkUmwrG9Sr8ahXHphlc2EqxMO5yCgkYpuaZFvRaVFASxI6sqUA9J2t+e324NoNv
yz7SR5p2VQRVVHo0oBiFpfDLij08JyL96d6p2L6ZWj3cEY6R771FxwKq6V6+8OCRlo1yAb4OuWwg
2xOTALu1xoht3aP10+lD/9F7PEqkwCa6zSdcC/5/wD0V/MGFVlOCtDgIiGafIYENar3sW3iUMjjN
14BE69OspGBY/tHXZiWPKi8xMDg6IJmnLZIn2kPp0/NNv1Pg/yvwyalOQjAIjyZpObuKWYK4h69C
nUTAR0OoS4DgoOo0pqbVOPqoe8xE27dXFV74ycpjX1ZRjl3gqmRz2uiZx2s1KnFDkwhV5G8KaOCx
s2D+69RBDTxCgTG8y9sFhBdcFg1xBU89qtmj84qvhuIZgE+nQQZQqyrZREmcXtXTCmhNSrQ226Wo
6EU0xXllhO1+UZtW5/xf3dHt7fyncs5oVk6Ndj8+NbC7vArWkC/hObBAuf6RlAPmqRNlD7NBMD2D
uGdFbnnpPNieXiZWgebBYuq56vv3epowW/zUrtj8/jUtOxvyVzBxnTbjMdVx2AQhZyPOksCvXZQ8
jdZRnjylegFQOKbVe7uPX8RMZk3SZgqINdkK+TWdeaKASI2yxLA+CSC96vJVs0MNZY4wxqNUL5Dn
YYIp9yJiKyvcuq0BDUoFHz7MSa1fiw0uVdAVX28aSYLJsjDKZ/aP+CzuvL5YBYbh7D1rvRHlcA7A
FdCYgFz27hM/lAtKv2ThdEZEzkDmU/HTZ3B5t8PgVuvRhhyDDEZY6E/THckqNyF0xXhZZFXu+GJk
a/S7t1nsjZgT6Cqa+YI6EHoJ5jlJe6P3PGcFu4A2xiR27fCdc7m4X7vLZ296pfHxEEgpKNPvW3+M
ueXL+ybwlmrTI2vidFGpa/FlOqSEMySsf3m6ze3SwCV1H2dz6zGZ4fx4WTNvQXsdhcB0Q/AdDrzR
JZOZxVpM7Ro/9Dv1++OFVItVHhuhtmFzg227f6Gh7fWS8dy1Tn7vAezxNCpgOJQYHmcyN/s9mTZh
cWDbLpEtiVMbBuyTjvuNvng0ro1QRXy5IvwkvIHhd+B6C9Ie5oqX7NN/H7nA1VxnZtF8ZTtMmqIc
xjt4PGHR0VUcBY6KOYq8hp+rzLTmsJnoSC3Geugh2/px4OnmqYSUZ0LyXT+qHrD172RAFhZpxUt1
NwsfQKoVbs0B5FVX2maWiNGS+m6mRE0iTNR4/UC6JKdoPH2WRxm5qgMcuDJmJmYXh0ebhmcLbEEb
4R90LstndGQXPNhIooRGIvQYeRtwf6hgTHQ8ybgZInRGZo+QMRGG8mqc60h3DZxwg0G1wTAj1cjk
+fdFaGRjM8uYAEWPvJ9+wYW7gxLspr15QE9xYGgpg5qfivJQfA3JriI4EKyVZ1WIdp0YU889O41j
Q0CY2j9YfxwcSNe5Iift69mjAnYbRykAYAWj+rPTT+iqOPUYwMWyNm/yCQ/OChYo9D6wU6V616XJ
FOcKbEbj/Nb4GNkEIg7kbrp+EEt8dQX+Cn1IZgiT5w/istOEzW1nwUp6rHPzv9/xcPY6fiFTPmBG
voipkJaeGSuRqZ5vcsfPIkYOv6XYYypRlcJDUXIrjx3/+jD9NHAT2avRD7fuj3cLTDI/JedzsM8x
XKug3x2cs3tVUhEQJmBEJWrf3jrI9fCZlCKgUvnJfERoI6tjdjJwqq21gcuH+pVddCqoLTVp+jc6
A8OuJuCzKVDdeAnLtpqZLy+j0pBvz63i4olqJGEFz9RDJ4eUDpLTJeQVrBNw+E/r5qwrtY9NiYq2
NrUsTiUc8BDzjJnmDZNvwm2zuTfUTQzSS8xs3u4JMx7nPeKgpado0fuwrDGxrYR8YyF5SlKUIvbc
9wEhsPsF3ZcOL+DvSw+KXIto3Ns4nNElj+0ADM60NRMpi09YRQlyMQrDxNiiXs+Ga0oipOE8tOPP
Zf5K7yfX0qv4jGK0VSSawc/sDvNeX7EGsoXGtTHztVUjNg8nWtQ6LWw0qVuKkr0NcCZl5GSCe/RD
6uCIIkJxHqcqeWOQN7II9zxRxyXFp1WP4z0ANAZGUbAzV38wNBWA6zpzOGCj+qCfon81LTPdlJfy
pBy9Qs/XyjIihvQwfISSBEyts29XtJZalN+VTtuwN4PpdAgi0sQ9JIz1US+VrZnFkCZ8BMTIfSpA
I3f1Hpwz51y5G+uO+OtDQ9/LQsQKeww87PkQpjN8gzBSR+U4idzm8dbDNkCDKooVTZlKa4ZwGwei
8LWNwzorn18JnFhG9NP5dTnrB8CjLgmucMsNljIQouhK6fNpCFTankWLcvnlQOk2Or1pV8V5se9r
JsWoqqOVzbfWVxn4ct3fULbdqoL7SKAgNWCm0rRAv8AFrkRdvtKH3xKH85FwUI+SHn79wyiB2kYV
zW05OYQx/V4BiI2/f2sadRmBJVKoB/i6Zujx5C9l3vOytC3hfGmTBz1xci1nrRv1/Nr5bi6IYqfu
T+FCsiHG5xSEhUip4rnVCJ/oyrOGUqSz+5t6Bm6eQKVQ40ilqokHRFmdg278SjdHxjN2Un0cKRkh
K4HVjLPXzPwDtz4gVmTyg17bvx1vjhvUacLwn2m82zYipEKvpTJIJRhEqwig7GDSD0cIh+tOK3Wh
RVQfwjqglqpdQWOAcBqCDGjjCTkSaEUar1kl7fT9gAXKA4bfXomZP4INtfF81/Vc6Rew8d3ZKgBs
g+eiL9OR+xvxfhnHL2/9IOuiVyhLm7zxCsRCpXcEtC6lhl+x+n+xvZcVp38/MZX3SN5vDBpxAEGP
8iXYcGtzJbolDPlUtTogBHG+GzIrcXbdWrt9P/Gk1saurzdQ5gGWWVa6PE/lsXoQIZWT4CCAg2E0
y1VXZZa1miKsjW1DynDW7N3Iw02d8Dt99mgeWpnHFDklPXvSpmO7ArlGbMa+qjkXrVz+Z/cGFEaH
aLiRgF1FhjskLJ3xn5I0YSfwo58ff98uOKlu6uxXkVyXQRZRGiAmBxjmlPflkmZ7csr6dGCpq82Z
Fm2W3TT1DbAPAfnQvvryidSfd/sbXJHxpZDto9VMvb4sbOa9V3N1942BrRNW3ge9ZAJQqAJhhpa9
mI9ZgV6lCT2uqEsHa1/3cnE3cUY12ux5hEpNJt/tyy7OekHqZ31tV4xLggb292Hea9WgQPAT2Xs3
83cJWVb3iDnpLDylSSSjr+hrJPUrzVQ5lYwjVu/RqV9g2g1mtwxUrhGNXs5HyG3FD40lpX3KlTmD
bL3U2moORifmCePz/MfiIytYNNTrLsTOmzzMhZ3GDNMgssyGMlM9imx83wnH000y5UCNjTlMmE56
h1YZStje69Q+D2QNaMocMfdY6vabKI9vk9Fd9+9pZJUjOmszuZt52k23+2HoDU6yAT/F94IFqflu
3kdTX2cYBX9gQs5/sh2m7A16gwAT/POPdvhqJZuDPoGM5fePcl96rSyg7A2WVkFLkIh3YbCNyYlc
K3WCAG2I30XIJ9k2xbe4xpjnx5FbnKIR0Jh8LKMsUtMS81Z55Y47ii/PEzFyvSg5n2njGkol97EC
QObO96J4EW05Y6oivbovVCp7VV5Rpg69hymTZVZvK4oVjt5lAfvVT6gdooI+zpQzzrVuGk7lk8t2
1yoHIvcbSohvDUqunqgqYR7UeO13wZWxjEIvyUX/WzqaprsdceqjleadiJg1QAm3fvEzvrxe3tdI
7aRZN/cgMXG050zM1GwtW3J5ijAf0xBb0ZepOZO02gB7DrQz1Uh01t0mGFOQt2lNbaex60csxHg3
7BvqPOWwVEvjeBWesY5W6mroz9+Be++2h2vnBE/Ocp/3A9cH4DNLrEMiNqmy3oXtEkdKYSvlE4Lz
njBX6wkrz6HUagKqgjNxBUM1UWWxmk4ctSoIdCZpCmRtI7feE9ARKbYIB3k7GzE2Owd8e6+EF72J
iRlIJJoO1MphuA+50nh8e9LxyAoZBmc9Et046VkZyZWuBF9GdsvT5nsWBRWKhdYfvfAm0nA+ZLim
p4UU2L5vOq5iWpZeidBwKhMw+YcmogYTVLs62Mu5jtEA23O51r/kP3XWto4X5ranuPgFBBU12Ttw
5wPWlRgyPoU98mdq+zWUJbfS0TnMuHAsnFhfi50UzhEDsCfO17TBYRLs/+T1o5lcNDG46549GQFh
ucG8iQv2BwBqYtEoQW8sXs1wIZEPccPyAAkQ8i/2v/lnVe0sK2UGh6/ZwxterwpPEV1haYJ2pqp3
rikwGypy6Yfag/HXCrO6ewq7OtdhoOQD48BO+5qRVlZKMBMcnnDOaUHV3TW1EK967i4qdEGxWUpO
d67NXtwQkHqg0aj5M1ifXGGZmxN6cV2WOnYVc+17innvgIrw/iMTv06C4Rfl7HLW1UP+KBGpb97p
EYz3MYItFjz5hWKlZjnKsOg3EiQcraYNGZX2XV0YUDcSN8u1zoq4kdC8JVfv6mDSrkbn9ONElR/g
KVoDLRiP1r7p37WN0eO8FhUuAx4r/zNpx1GVmR+71fvXsQ8i/XvI1sqSErct20OpY9YRjTPXdby9
O2YQrxn7ujZpF5KioFBMD/OGqJZBErUM66dcCayF9R2erBdQHqPOEPj6wKHQe0/7jYmiN/WopG18
PdmBKQKVqSJKvNXlWwlkQLHbBhjkLmWhP4nwUaSFZ43rTvyk2cIXNH+hHO/TXAaFchC8BJRHyKtk
0jk07YyIDieKGds4YJx7sQGEkakOs/KTjoJvpdJYm1aPy6io2dHHkSV2akUzq6ythTapQnpgqj79
G2BL2Fn0olxqJD5f3Xoe0tMy7/TcjCOhpuOCHFV+ovhnXuCO0XuMmQ5WN+X+2veq7lL+S3ckJjw0
zXEyLhT80lUE4ACBJqPrIHoYoP6p+9C+lQ7l0xIAWXR/SBrDokQk2835I4NeqyIJIsWAqOtlgduG
crduy6y4btPnqHAcdUMN1YIcN1bfc04Vx1ceesIDU/6iSKD6MinaXtlQN+vZKqdXfFUDqoELgNUm
XBACkZOXDcttY3Th7gtZwKfjfAXPgORoWBNfNEs+HNpXJYhWygvWH4q/Fy49c+hfQVla/qUgu8Hv
I0+WRF6ClbAtnr43LqSHGKWtR6GyDyQ8fk6iBpdSax+Gbxal+lpMwtlUQuUrQe1mLxsaVBXQTZoU
0A+A6SS6QVGrbaTKtiMWoDfMtA9SFiwt1rlsJe4cNLXhFb27pvfcVVIR0q6cV/bfCe8Yb7uuWrCU
sZPvzy8/oavQSwQkuyE8aZ9UBLLC+1QqzPyeK75JWieirPjrrnUhAs36OLXjttQ0DRlD8Y+m3hvx
M9W8qHkmSeURzACymI//jWPQT3CDLNyBYnzxhN1FttR04Gs+KO2+Pdc27AE+L8r15Xmu3R8sVRbE
ip3iTzWY57ZpCxuDNG9G4hZoUqnLJT1T4EWpqQFLQxmjACr1PinGfNAZWVgb9y7K82AjgNTeVgrM
XsoeZDgXC6yPs6/+PnpPbVWHPmzrysrxFPVw4anzhy1RSVwjGJ7un6WTAWeN1Lat9bCm568t6NTL
LnTONrsqfpE21zlf+T8WSCJIaYBNOZLuL4gcd/CfkAAFu6f0zz2GXXf9n4bR2Dq0AHMJwlFp4L3N
mQ3DwZylB58EAmJ/4UI/DXsliWKBx2uMAGB6TsIzfguhqgRip1Ja1Z6iD32ObMYMzMW3WR8Y4BPB
48luJ54RzHmTVkYoFZnFzbAat6bN63B8wIodrSzKLD2MKU9nXvuOCSY4reoCxb/FxrVdvsyxztGx
V0pfSs7IfGDMkkDFo7xdVVdJ3xVWFGAOuZgwy1ozhiFsin/DNCK4rh8H1gKurJ4OkJtiyR0V18PY
ZF795k24irOFJYx+oxzjGV1lrsndYKslnV3RUYdZJk4eWUNZ5m3Hneaf3RJze5D0Q24BFEo9qp33
RwuvGYIwDOHITtt2nK6hrR4Sl9K0wCa3bQzZrSN03bWO3rvFtZDUh4MMR/Mtg/NcaE535XvvZdGw
mdwnpCdkt00EAqtaGJU+ctGLcwIVMwBZa4ctyeCQJj+VlkuQg8t0rFasCXsYt8cu0rRmhpa5h/1X
baIRYay2DBFvKukX3PEdVf5Ejpm4kyFFUbTbXGWieRY9O9EVmhaRPd3M9RODTh/WUtp79L9wVpEB
/VgYbejvO1D5QQdrszQbdz+oZ+ipyRg4i4fB5NLMIOfbBQhYxsUI0/Jx5xeLQ4RT8PIGUreVmBCD
zivoqjkIsCfzFPfphIH1avldLPK8vwxu256+OJcG+62XcAKG55+0T9Gibr8Vr17Mt03KDcQKDkqh
7/2sbe6AUJx6I8tMLJPh5LEWVtK5ZdvYz21Tge+OoXNNTl/qxKUEMILPbuHm9EP+zTLeD2qXe6hI
Xw0uA2/Cu+Z+YRh/ITzWPgkJICqjTpTpuEDBlmITxzndjt2cb+2bOKLs14Mlmpsv9dxgwPYD9duP
JtEBUCCio9swr4+EU7xPxeGbifCj5kuKzo0Aj9MfxB91j37zc+kDU5IYeg2QlsKdOlU+A0SsnPc3
XUabHouAIxcLrQRObS0hUt853v5egi1Zqpy1ad0UaVNRMO1GXG9wwM9OwwkEAGDjZk7oZixpvnXf
UCBQvKLToFx639BC6lgPupe4v+2ItYqc+vEraD61Oya34umQdVpTC+WkyNiWo0ripNmXkk9nGrxx
8XDW5161DMERStvHJ7MX+d2TAzcu6FCG/WO18Yry37veAZl6TROCpCU1/uJS8BnTaCA05hUb4B4g
XJQ5Oj3jgWuZQj8FFceTW5agoK1LM4w2/Oh6aFLr/B96/vHWh+vheu4JXeXCUVy36vHU3XKrxE4F
jHT10i8UuyH9JtK+LKgLtuvREL3BmFxeOQ4TYKj6apFuaTRxxnbZDFRXbKZiTPjQmKgeDFCijSxa
W8jzJD5PHMtG5L/RvgGu2GNEgNyrcoCV1egoUtO1GxAsFkpUQO9FjiO59zIaBLIs2X6W3gBqyGtI
fXfLFJyrRWfMWQk45GYvC+kA+/U9SamWZV4qNOLtcC26kM8urrcULFDec5jqFNqVW8EIQVI2t40h
zmEWE9bBWVID57DluLQcH8a8LA50KKprgoobRYpXAlx0NDL0UubS1EnveiYdInRMCaZQAd3cTyrB
BMeKAU7yqSwkztdaShmZ8dRghhBtltRfUUsTCDtxCHjJzU/7eDH0cJSFtRJ2rRKGVhb1JfKjhBqI
ReB2S5QPDuvE9beg4DDt9pyXP3MpFwDrSaYu2BKWD57ihoUE3zyWTuZdXRjYxBt59tT8FK/IJg+s
WtM0VQYkvaZMq0JTdjKhNn5B2P/nZgJgETP549r5a0LWofzwEpaAbtfYfv6aKEzZ33jk1bxOcZZZ
Iq3fgqho75r//HvErCr89HCW3E/zmGGdZOt+Hkf5d0leA4NwenM6zuITSsDPHhf/P9poz25ZYPOz
5dO9aTAJ3W2io+3WMC/AyJSdJbdvUD5BLDSnaqPUjeyVHSeUmsN9EuvhJOxvlSEJBwPaGcqJ5brU
BcqGneyPFHrIyp/z26bB/9WxBtNT0YKaAzjW9GFYKsquxWdMII8T+bBffJz/u2CWMZS20n6R9Ogq
rKnhjezfhAdhNPX4tRLIEwaLQRyljpuArxTGwl6h860rMuxGs7MoGKKS5e7UpDgF80BqauDpS8Ti
u8H7sT5bE69tjbKjkpQ5GOlM4nrZ9YNekpzfsMHp/qe71ZRhgMQaI/szGFbSIxLQTAUV7eVvgVln
j8G/PYT1+JrL79hnoPThY3mQeWQmS+FbSRiAt7AVKNbytKxFbekyMn0pQY+Q9SOb9fTxEKyNRT89
rMPrggUxNY4Nvxdbzo+XVxkAYURtOHAaTUBcSbSD7F2MnPJutxos4qSC0WPzQNj5FtHkwMmbCVL2
YyVaxX19ON0JVAnkXsFdxyfdbl/o60BXvN6H7bhEZ0Kvj9golbz4Vb3zpxoFjaiC4IpDNbc7zwFO
0x9UolHUEQeAQlfj+K2ZbkKicoybr8qbSojzLhj8pGjUsQAHf1s1f55QBL13AejyRcvgsROrP3iE
OtKcvx5tbHplrk0MxdPZB+9SS0QD4r2O3i3C65/25eVS6gY3DZzbyzCiTYjVInfQYSHky8tJXiox
KH1uaSCH1fhr6C5LPoizgci+Nu+8GihfOE4H/q6EmgcoJI8Czh3zLQAWDwqd/TDZcYdoXeqXA3Yl
QRX1DsGHuKb9csfSt12bi5/HxJPVxAG00k/H6j7+thsT/GU1WS0d/xvaRhvroxaeI1Bt2DnoTUAD
TU/s1U+q+wu+SPqk5jAh2hucBCb+UooZLFm0LOvxpzDIquJQ3oh0R2kWDooDhNveCLLE2jlqInFK
rWk5uSES19KCBYaW8CIAgXl1xrPGHGJ/jx7G7j+iQgLYgAuPGesNFYu9ZSQQlR+t/F1oKAjQteQi
tnYOfJCtr4C/t4pq0ro9rxvZtiJJwA9/f0O7ud6wauGnPefSPDlpcTa4ZbqGDEz2S8SlH/uR5lah
TnP3o5zbA19EYDMuLC992KLA99oI1PQ6dit31NOQ9blKOzQnyjDjQp3UK97WQCVoV32bvBHH/+Yd
Bwtop/KR3OvHRA3mXu0M/IF2CC3ZHuNazAM62zzd1w2rIAuBhk/iUx4TK0SHHr8kRjYaz5d5oYxW
s0ucLI7bZoubdWIuy9qpTWf/FcaM2GfUy28ldFqRD8Ue8VG6tXJgWqz0IRDWDDTWe0iYiXBVjwpt
MoeDyEk6nSrX0BgAqSYWCMjAZ1ahJel19mf4MFyog2vlqxRVFf6mcYPYQT9S5tzLMNOr1cFDOsnp
B4zqpjYEPocNpCE17Q6bYnfjLhBdn9owKN+GguvMXQcDunpFQOOUz7Pq2noKuUkpvbEcgGd9cFgx
AmiqSMTZLOWl5GjEHeh8A/56sFgLDZLvaZx4Df+z7NVEEMKgSMINzElmGlMQ6cQ4r8k4JtGSqcrs
eJm3bj/9jCFmKKa3IYqIu63hFDFv/1tyFu1N+xvM81OeRIe7/soea2c1jORzr5vgmZGp1EKQUW3S
H5aL/lhFz/LDXWt8DfzrL+iLw7vmFGlV+7qe19xJYoBzC8Ril5kN5x4eEZm9XvPSYeqfH7uYcvhu
t2piWYLJL/vH+/vjWiP05PzzrN9/aiCZNUMZomuap6+a3OKU3ZpH46Xn1UWkHAXxoR122q+ihQRu
vcUawhzaQQvbcWJG3+H5zV+4InIS617/o6APGYdPvffMaPGAf71sjLTcQiu2KnsnfSwtvoDewOm5
w2qnxHqeq0FFkkZB5sA0r+SbTFEqpY62XDzh2CNGSGH2XLDgVLBrMHKukdCebqvj8J2wPDQnI1aQ
g2KC7PlI4zIRuPpXZRIkjtAPWW3lGtuIzUEDFdZcq/CohzV8t74MJTUjXSV/HC6BTy3qVlvD2WpQ
GTkDeAJmzZUo0WH7f5ROVBobYvGKQsviJ0VCi1igFRIZ4yJYOtE4U95k8Eemibf9Fvtfg2jbMDG8
MGQ04YGvrXOyqJswzOvCZitPnBghUgJeQPpAbBxHrOYwBnLNYr+b/X2IUlALxrQp6TpOBjTLa5Cf
cpENrhtxx4cZe/qANC+nDa5EUNTesIH31c4idDVFm6MxF1uCpuoaYTfg2prU83BEU9l+GQsmjbf9
6nvUHaIuZL4CN+BTqJ3tfup/OAkEU5x63ooiIS8TpNagZoNhCnXfoPQ6Uy10X+B0TRZgcU6ttCFy
fkZ4TjaX2wMlkH3GxmlZstzEzzGRIOWNm7T+UJdDu7/dAzoGDgTPokNPKFzpdBG+W58PQJ07AoBW
yOwjfvkUbee+/1jq2EOoFNcDIMXDpEzgIDGdvezIUGAckykqAt3rPCBQdNcxY7Qo6Gwi5zTFsp+7
e9DX3fap6xqYBT6TsO6mk75rG/EHlCMkeHs6jScxvVyDgpfV6I0QmRTGVkhNNTCIp0anU4kKtA+Q
E894800IWjwC6bu9z1C7UP21G33OdlcyQ7UxWNyOh1rk5Qj2/gE9yxrhqiGMZEZ54ujC+i5sdEQF
tOfXX0OWKGyRB7+ASBAz7UJjcJBdUHS+4kmTzxN9mZt2aqoBucQYEbpvwcyJdjwmAA7F3bK7uAsv
/8vl7OQKlLWAYztF5MLKvqbjoIQhg8qDTXzd/krv07atGz5LxW55Coy7GbJWBm0E6k7FxK46NxFr
ifoJHrkaoybh07NmYdl6P+imxRhlHsZNKXI9puoGGR5NBXhTIXdt7WrREPAuRJGu5b2WEIPUgr76
vJSxIXN/A/cmHsiYJOPn4Z+mIfbIvhdPLpuV+CQ1n/IlIwXRbfDyA93fw6/xTv5uE0MESnNHV5yM
CVfLSToyNG+xKoRboFC7hr16p4Blfs1CtoQLMSP85WQQJ4ebzDBCCWM28mZO1Znff8JXgz7YDlFB
0X05fVbXVDNk2y3Tt6I3tbFpYzy/OETvIZm3v+MJkJWNgJwaZWQRudmmme33bkKAfoguGPUr/vbL
Z5yFXNsBvXPyg7lPRsP1HYQ02OHExetUpcANfPE2oEi/9KkGpRivZlW7qxcoQLcISrOxlNbzFq+p
Br0bSj5sIlxSzu68UMKKnszii2Ru9u1iDOsUvZFrg+/vG7ShwcS4A76KckHTP0OQN+5E8AzzwP28
snykkH7rAqFnfqf8tCZm6/mt3VB1irOtHFKgstuGpYLZqLD+Tich/QeqTHWitJsOJ94CHw5uFBN8
EoPdYoPPj3I3KXqSUcvfdruXR46JoR0BvH0fyZVzvBfezAZRIkKz9tACX3F9lEBPhPKFqJC5tBNl
fssl6oj/mbWMn+VoG7BU4icpIYozzO4w/8ETm45soDEUNDK7OADpjCwYdGvYfSe+Y9GLR8z2+OmE
GkgWaH7N4Ef7r83WXwoBzwizReOH5hCqmqs6/2XYuOe9IWYNtnU6qAXL8mfdLMTULOqUwnQExBX5
f4aEXW1bDkMLKftWUOdxJbF0+7ZEFN/6MjPJ3zLHf/pvvNBpGczpT6Rsz/NteCMLoGatoqMpkpOw
W4WfXnQeM3ORhCXa5xj1CxuTv4poccWSDdoOKLRFU2oeMUUNfrTRXcq7MK5keHg237tv600b3oVO
B3hGIWApetZUi+8ISSSkocI9YsG71zLUX8uIKSgAuknQPA+djl2GFM+cECMuaV1w6bmqULpmNdiU
WDgnfeksT9tRSEIq7iPdD1ZpJlWGqw35jigHGdWYHDdjbPcdFdvfA+Gul/SDCy9wLAVjwGVPE7BR
gOoSeRyyQIaw4Hvx2mequyfC3UIeKBa1l4deiyRoaJkYW6Tc/Xi3OB1oYVizxWlaGrNm4zh5+1bV
0zYkPfKJaOOraMSJc85BGf+LzG6NaZziJ/q3Lz3o4B/DpqzfgP8eDU0j10Csy6LsCM8O3eYfF7jS
mNVyTNwr/iLZYSJmKc2a8jzacLrO5UK9HU7L55BYU1c4dAdvpdI5Bkl6w7X0sMMtsSafmIEzo3w9
19DtOu8o6AprydYT5KWzEd9d8+bxqYgyFraBrHZSEri0lFBwDQJMBlKq8DRYIwtUkLZRTg+XUaqX
Q2W34MQwVJUL9xWbvjHAkMD/9x41kceA0NqcZAGtcKX6RB6k1jngKe1YLo+YukYeXxjwRqXOefzZ
AE/qRwCTansPToiITJ1H8WaaSRmgYFtZ6wusBuVzLi08n8wM610IBmyT5XTxZLfFzGNAj5R4pXs4
xbIb53B7gP21qhSlMFfgZ0of8/RLlhoIebMGl+BISsni4WvWpTLJ8m3fpaRg7RepjRza1itwP0eV
MK2TdouZmS33KbOtlPyT3Ks8doyJtM2TDYQuPdbTuMLBpdx1gwXAccPR0LK6XU/wFc4CirzBmXXw
Ap8VWywh6tNfVjRBME3B0iLZxPhRnGmQd4l/2w2gCB0jAv9IOGUHXsw9AUCvjOsaOFxQyLVFvijl
iX/9YQELzqCqnszaMfQi2RkkCkZVeDWsCea7fy22N+3r4rq+ET+OqrT27mQklec6hpLIY5F4hxH9
+iH4nJ+8qeaPVfzKUZGhpwyYlAj1L7z5KL3jS8ofvsiMmsFg5UjNJfEFc5Kl0rpn6P9gdq901ULl
5DMLD9Z327eysnBDPgPq8/qnyF1ntdBbjvRZRF7ZeUC734rTMGDafpUQCAnDJ99iKZLq2C2rqQiP
/w+ckXBWupknIE7Io4dfHLw5ba1ZfJW5JcQJW1fC+rxBFDVSfkf7RbxesXEL09PDNSKshog+31FV
gGYM4olLy9pDr3Xfi1HGtvitlZgvm3b5lyc2iP72p6HMIUqhHBxq2H3SYJGaTscNjJ3vwEyqJhM0
AVtaS9iFMJG4sgk9VECnk2ncXsUZ4lAw5RjPQvZwGu6/m2aE6Nl536JqJeU8i2Gxj9z2mCApq9w3
iYYMWzBHgrYLSFBxgHa5f5MWtWHREM/6rnN0tos7oPDAsTBOqmjCZzKXoKZ+rNPos9QpsVFB0ukg
dugopXV0ydBgfI9zWphbMUibhziwHIAiK7DWLUwQbXNzRb7vaMfILoz8BAidBW4kNY0dRlWy89iy
sjfNH/GfKZ3/xWffrQKFuJ5kBa5ibiwUQNUMs37xAaOtlf1con0mF5rPFcGOxESVwKtzF9ZXyWPH
UcPsFZQPGlJDvPTVpn0ftYpcE+CDxXXCqIoYtpEt+cy3VIoFIb0a7JvwCPp5nQxHxhzYR0oTBTHU
WwbRpChzhVEG6h4lpN9eCksTZh3LQPUdJrOh3CkpXzos1UDooINRkpCFuzt0mMO4CDTZtG3tGD+8
ElCVD//qgvIV7LaoIcl+YnQfM1p7kkFwsY8tDSDtMtrd1e8Y7ze5tcxr/dt1h0/y223uH+aSe/+Z
Bt+1X/cvt2chfzwPFS394elCOuexQGQrVmrq+o7RNL/azFbNty/t2Pz2T8YnW8W57FY+AcNp/l4b
lnYUi/b5ragpe5rDAMC+3KXUQzlU3scjjubTcwXaSDKWMXTKz/1oNCJC4u4CU0OxIlN5hwXtWLLk
qBnJ+t3yo3LfY/uMcbZG/dmtXzhe42nlsmqyrxu5lsdflNbLSEouy8pdUxaU6mupoDyWCJZHFZBE
g5ywzrhPCCj4TTRAhWq+0UNmZ8IdfHMeUfNaIX1to1YHwuF5CkP0r/bZD1QI8qZ31humQb1snGU6
Jd+Zfr1jnP4sUCXHeSh1BYLNaplXmAf6bXSqoq9ZvUXAziCCqNByLRdlrsuNSO7p/w1Agt284321
y1ymML3xKtMAoXdxtUPj4M0oZzDwZ84yAfNbsu8pxYwXApCRUnH9GAUE1wQHzWP4sbDuo7OkM393
NaKl8v4/H755c2vCu5my9IwkVpwUo8a06UeheZRO5maV6hjaG3LxXl49aNNhhFNiXTgj7gmMMPGz
z4FzLQNAOkcwSCBWXk6rR4a5ncKFuckk6kv3fYTBx7Zu5C7zqZmHfLq9826iyMIeBQ71MmQSWY/Q
tu93vlTBZYm1pVJLGGQI+zquGWrGHvNRiPyjVm0XticWrFe5LjjQbXbILpHH43sWpuvS5asyw1iq
yGW9oHLkgiqNfz3EjNo1xjc8IbDWvkGdQio0pHq/n+qlkTcHr25aE6EvcIGUpY3ZlTNS8mK/Zond
DoqxNwKZSz+vy8jCNLZA66LErbVtq0nVs76AwTGZqoTQJ+8KrPVpbFMJkIiX/iAWg6Uv93nLks4T
vCWIvSSiiKGQaM5MmeQKYIktJlS112nAn0GsB92ERw1doD61YAsLje3c1VBpINebuvDpSjmXZJHy
agqtaS9k4Q83cKEwB+eh5tKHG6zAbciQlVhec03e43YpCnIaWUaOLDTGbMXmUZzIKkwai5+svqIq
5iddLRzoF8ZH6VAijXiG7S9jbrkG+1gloFEzrUjPihDfJvCXCJpocWdnmbRRA3kXj3sJpy8avpYw
ET6Wwk+vtbEK8w+2oOKoBaZnlK6ePHm9k5Z24UgfwSRF10vjj2/wqsRaM70BH7uYjOWp7JnsW9hm
JomwZq/2BOijyiZCOHlLuzR+I+5jFkVi8bfFhbm5Upv/9a0OYu5aLPu3eaMV18pByeJtfn4xKEMC
E4v0Z5s8Bny2VTXgGvK4C9CEDwn0bhmH8d4vSLGOozTq6Kri7MuVJ4hzZW9hBO1jc9/ees7C5Tnp
CTyVHDZKyl50eu09QYvpfiYFb2Y1uDGZxndPTwZzNc+lQ/MDCrGfuC4JICq77h0lu/k7hsrmBxLS
bg8fOiYWFva6lyZQW8SAqR0CR9pramJk29Db354oRtoBS6aWF+bTsG0pMVkg6LUcsyuMXMx8jFK6
B7JnWCE0Xc52J0kEcugbcw+iHDmIvUEOucXUvEOQqU8gaqabd3g+JuOQmUeOhY/q/MO/wKPVKpOO
+FHX2w2vy4qBAPmjzB3wEe927Yu+738KRnPZVIehOs1RVPKZ5CHxeHAx1nOsNkpGqih1iL1Ept0e
7/KcAVP+oEFdMcr2mylQ11Lani5bjHQThe/oNhqtw78aLUKDw7W6nos/Go6SAOnrywPfRpIq7gU3
/4kGrcAt1a/XxAh0fzXtAQqx2XJj/K5AcYsSnXg24Z1XyLZJD8LainrNODC/49q8KPfLgvPn0C9g
EADnTF/6qC1bsBbHUi97ro3z4eVzw364o5f1AmYrwaMQ6OIn5SjGsM3fccYI1RE1apOELzZkFXnT
Q2lZuyxfbZYtTsnyVkDeMvTjuCAxAmMMsrt6GJjFbJKzxS7ybfH39DbMEpAjpYjutVGgFwEeQki9
sT+cXIWEq68h2oPwZAvEicGki+YG9WKaqnK1j3N/Ro4HZMELBZIU04H4bIOnZxZQS4e0FfeczHVk
yvgZKNZuOeMqhX7VA+2LcQUrpDsL3g2Tl4Y0VuJgeavmdM7Iob5R4LFWJPGQLLwnvQ4epF9XAAgr
X+sgHZkE0wa8VH71ITFuGUYCaX1zTyrML4IYse3S0hjU6K2w5ryAjKG9es4W+Vplh4UpE2vpg9xu
3Ac1f99pC2BYEEzsPBVNddUrbDEagJx5U5ny8EM9lZaAGiehlyln36NLvGwl1AiEYX5G3FyzhFnw
5lRnoXlGtlJ6FzpyXfkii+fpoWhuJF/6w5nfeup28PKRh4ksFNv9oL+kVFVUEfWjvYdbCJbf6UJY
qajwcMZ7aHY3bWvlyFZ0EC/IE/DmJUe4rZxiMAjdvz9o/wBA0khb/pSR9KLudWkUBEM3/Qh/kTsv
YmFdwP5UaRisSkXrAdpEVA2Bll7LtqUd864L9e/UJ57xJkNkAU/0biBVtLaebc6G3XJju4mUIxIG
noIKZN7i6Vo+MXOgsIFXAkmIYxEwjap3kKR31c2XHkz8we6zk+iRT7yQ4h9wfdGXi8yvpJArSBnU
iDzFmEWCoBnv+iQ6mj5YV57my7NWyjNX++WPrEL9PetVDHhxFNfjutSRXNRXbnpMfRtoksKPrmqU
g9oBe9EdrcORucwsxbCpcKJA7lcF53MPlnRUWUCqa0/uXE4C7JDz6BL59cscBfJtKfoTA8T9UEbC
TCOiBmR5Gql39WOH3HqF5VuwQ5V0qEFNBl5Nm35t4/osbTcHeB+KRFYZmklCBFCbOyFptPLlllmD
OS7QHU8v4rzddbUhbHc4ojP/ydTSqn9Jxjdhd3ysWN1UV/DTqtGUOBl7dUOgd6LqwD8XJh0hTKi+
PNMd8sPqxFk59i8cTx6nDcyj342IK+JmDjOrOtkgfRd5yLJCPuro2jkv6F+F3uNiVS2AmaK23A3Y
7/+uzVXLcacLxlgJtBS5S/EPkiuaawYuecTI4wMHk2ytp/ziKdRdjMf1mS0OCtb7k0kI/61DLG5Y
iUCB/lBKFGlTzHlSaMK6AwA2M3MNPFfTmCTiXZ2IMPDKhyoGsKEYXuLLWpOiQRzR5+i7G9nn2WNK
bv638SoBIXZqi8srx4QeotwjrV9T0WOvh5ARGzbVSuyk824Flky/T0O7oWDpLqmkZPTieWqbZ2uE
4R5g68lkBa037bH3jqNufmkEAbtcsNzTp2dFHm5Rx8mLi7N5X59eJfSw7Gixgkz+gDZvQ10J20/y
dncctoopCbjigtHVXrL+KcZ1erJQ/qAOkv8BfBESQMupiD+oSDTQCnKBBp12kZ2XBhHChnXZD2Dn
RMMVtpwJKNfVDWyCMwAA3e61Qyss34KOt2rcCinfLLTpsDjEoC1xJ889sLzAY5UYTx/u9fWnX0ag
kH6OoUFfG27nOM+nU3j4/Xe5qebQOp+e4MxXP6G8aeKtEfG4PM3bgsxPtVSHVS0Af9lzQDktaHaF
YshmnwuHtHLdwR1gv0Sv1FSj+g9inN0UEbsuUxJjrQTt81szNWMRAewDvbj/CTH5RRQvvq047Kby
wioxjuAD5Y4b3EoAtlCF5XBGEBT5TANXDbu7NO5ZG7lKpGOwCLOrBSl1dUqcvtRz2k2zFy/LL50h
jfgh1Oli+WTuQqj9uh2oREvvm8rq2/WGT91UrXzFsBegDAlHpEJDGrjMFXCRL8/7cQeXK7bVXKhN
lbzNCK/egprNsJYrsiQeK7BE2VuRcscO9NkKWC80VXE+5o134yRMJg2CoZdEAKmICUE3PFDd4HZh
4YLZ5CNTeC7rSvjTjQnCsKelsz2yFJhbv+lib5wxuW2UCtx6PK7Z4McejM9wT2seGJEsHCq0XZW+
ynHsbkOj986iyCJhapTTVeUzsVlwb7vqJo32Q1w7bjUFq3EptXo4E5eQarxE5mZnjNIxaybagisD
QSR+lsQVgWzOLF6EJ4BmaVXiNcT9ZdlzqNQssHq1+Xu4iOYGSWILUHYjXRikXjgxi8CNjAi2vgYB
gSuwQ1Xrn+yVWWaE7oHX6+dUmTHrm0ezWW1EOfBgYJSxLGeTsUHgSPFgIb6sGbYta7LyXPxeceaM
CF/MQjwqbUghxpTKQAfMocgOCy6RNgVAWGYzlXzM39fJ792mCUg/q7PubYW6zbkoPuCcoCUm18eh
vm5cnbH1nOLRV8Y2hClcJEV2eg3j7T696ABMcBnuv59ayRACubQ+OynX31DCTjvbawfnX9mWAzhq
b9O/Kkgl2DdY7FKh4HvzukW+YyPbtBvbbbtD2FPFIX4z0HA/NkBvqrXwP53jANA7FjfZRznyUHrI
ERV56C/AYeiFbDLr0vPg33W7VNwZRDnrk9Vv8Xv9O0ayQBD+zi2RIgAQNuHOg+FKFnQAJdchw5KW
TYLzCDK/0m2qZThDoysr2QQNq4R5pVncQMPnjA1XqPRZqASb7uOZk766z/fSNLNvZ+xYZsVQMJnH
Gc2+tfCRK1bar4FTWq20kwGAUF2I1+ZSqqvRqvtFZ7Vt63PWxU3NE9yXSa7vgPp0ugRYkrNlF1iw
FqG/WPQfSq59ml1mn0VaHp0gWdcOLkQt66mbMw8F7BAROnO4VqdvqslE8hYjVLrs20V8wTzA8oGO
BbvAFK2M3usOVnVtCRwVWufHXclyPwU5ylIwlJO0NBhGtaK4UWnDTIcVM/67rdd5C7F3tPVzCZx/
lVhyVUMFCRg8wV5+9O0uwqNco1AZcJO53IwBRy0n5QuS3zY+3OGo12FaFOcz/L1axGgqrl4Ega1m
JOMACbAz5iCEET1aclhq5qmHjyc8NRgAHrpqW/qJFrMGj/eTYnrlfWp4KDTcfUygC03HWN+L30lH
cbhjQfbnU5TDQ0Iq2R9NIrF0eIGEmQ/6qOfWo5c2hT5CNFdanAXhZ3gei9qVpeRg1VYcY+HDtL8/
p/eBotbSVQY+9IOBO/9ED/DjLHbYnRK73u94884d3l4QOTkbuuc3zpfyWyxRmmsJhF5nqIhwAoZh
kd+JBuympJfssNX3VdV9TyrMigocMGRBEnlK3ZAWfmK94f8ekb7Sv+Cyqq41bh/F/30Kam4tg900
893wkrnIoYkbXRjZH4Jgs6Wv8O/VV1tws52lfm2fe39ShOg3OozRtRTPHySVZCm93i+uG81R3HLK
V+FzkCZ1Cgr9/Btp00DRUuuesTSoQyM9eEdxtAx6Lo622gx4293kfV93IQHQshOP4Khga+QoO8fu
+mQFubRYjckRi87EDBStofDUqUZNP/5pUg217gjjAieJS7JXInNRpOzbuB3tf9OHJFcTRcP/BcLf
sw4TtGtwqe0BO8t1Acb+e0ixTjTeGVWonX9NCoGiip8nBV3ia1M5oWuFMOeFcG2p5YclZKdsnwT4
5KMdtOxF0IuW3qlp5fwv8mGB3zgQ2ZwPBYkvXuzD2coM56YjICR0yk2X3oxTPZ+8wO1TqysJuixI
4XlMXPza/1jIHGXF4QGKnuRueiBJTNWcDGDHjj/vX+NXAW5jM0as3eOW3YLoxL24tC5LaqiaJkc6
CUnTkpB0zavnYkkEqYrvE9gRyZqW1eb3GpoM2vqhFnDBIaABKTZjHhXNyo75cN7tykS+QPn6THDo
n/7Jf5wCY5NrCHNn7r4jDUxl4qZwmnIwbcqN1vdbaokQOxdl5HYwkSzidMsHr6K8LB0xOBWJhDhy
GGB2w+MhgjQyQsKW6OpQaYrB9XmomTHxq0jQ+f4HYj/pMzpTKpIvIFuTPILINGuMhC7cn29mr270
BxVgqhjVrPPHV5GNjeXMXUuYyIUlwIzacSEBzslX0uBxXVXX1d5TAWq24NLrS+wxEbjl3Zx3BfLo
GqY8MCkJxJvQicgizs20yz7wBwSurnQzyeLiJnvw8YzhR4i2ip3CsaQajZ1hEKMVz9RtVLqKzOMf
o/fQG6Eon9LeQBD1AQ/IIZPXst/QF06qEV3FHeDTYcfFTeT7PKc4COwpSQBTmX8uhXdWod4B9cvY
8Oe6uG+DFMqf4+f8U4XVS7xHhof2g3H4DxHueecoK/yNIZFMcvkSst4dL6B1FIHu4Re52QLjpINI
qAGTcP8iIa5hfGKTdrDKfZ1JJcYrhxJ5nLvbGEflXBpbThZOGuQLrKidF0Vlq2M2YIKyMxZ6b92R
6RH45vU+ZgCLkunSx4tEzTBiG5bXjomtbuohD7dFVL/m/AV/JsSWJmtro6NTXul2KhU4r3I/KeQe
DMb8Tg59NGUthanB19B2iefM5zx6N+oofXXdhVI1LVDJ8bLYt/0w4AtdNBpPcML1QoPsIROv8jBH
AoBMA2h5ZUviPQExVt749csaUW0llwZtgZC6Hny/GmuN80dyxLlFlDhtniI/858N/xqAmhy8iwz4
TY/YZTpUpG0F0oSNM2cUqToO157kfX7Ras3CnFc2HnkWo5CCQKjwjuKoo6Wo46euXtQauw4FBhbT
X/bFtKZ99fC2T0HxhmPVrd7QrklkktzwgkdQSqdi6B2o9PCFWXMDf3G3JQUOI7Rgj6QtqLS0EFWS
AVlWlBuheIu/VTepDs9feqF0eZ15flrqyjGO8tHD3HpYNhUpsuUmZ85P9x7EXhvLMNSx5h2N6foO
4kBOHL63u9ve+sveHK3cdUCX1uMNDsMvkwqmdI6NlvnBa/jh+5bzxlERx3D6fMf1ZWSLXqE8KmU9
qQtqclD1ZhDT38fkP6kz8vPzv7LoFuAZ2xNRtqFO055IiP5lCHP6b61gYNYpv4X+DHW+t+uhRbe0
SzcD3+uqQwxAP+ipEnvo66wBiO7SUqZuBz5uihh3U70f92JzOxwe5S4aIj8td48pVNpMVuGSLsUE
eb4p46bilHYO3JjPy+vOEr9wRp+a1MKWQUetAqbLqtaaV0H/cs550FEC8jXXgU5NxXHRB05DIu3r
rWAwq0cC9r3gCSEfdPMUutXJ0Fd4OehJbpCYr54HaMu46ZpiV1cJQXq771aQX2bBxGPeoBGSeOfe
ymAUbRc7FEW538uOagd2s5BX7y6aB150v+xrMul5u5+FndoxFEL3Da0WGb3fO9k4ANfJpkP7m6cG
6cJZjnMUElt/Wp03kfJogAmdSmPZZRCJADMRsIenF9+43F6lzfQYijQgoIf+tUyM+eSCEuusZJ/J
BIWvihqj/h+kJ2cNApAFfzPfqve425GxNsbj+w9prdOrbH1HC1ZT+6aqGx4kons1+Ld6Mkf+qFx6
b2qeC2/LKUs503vQwjhd3e9+OUDDbXfiJTUg3aw8mjV6et2TkJTnfMAjaEZpmKUXpWwMBLJfh5JD
y4XqV7h6PLoAUrJ+zoiRoj0m5L2JaHUB+rKYQXolSxpcfGjtL+/wUo/ppYomqSQtVdlsBi7MQMK0
1PbRnaoXcIkYD8ZIZENvrpcFohz+eosGJfOfTQRaqUh8YYoP4xf0Dg/L0CfLbG8sighADNVpiNiD
V/cCozNOvn2WYgNH/7Z2CVJ8aEqT6BJ2wdoNduRe8IJ4X11aKENBmbAxx/U5JBa62efZTQIjtd/X
JKISJajqswHFEH+ijz+1tsud76SoaRbmTjt6xOF5Y86AIzzVHK985fMTw8R3hDlwXTQeWdVcDu8f
GAeQrpQFE809zUVvyxvMeiN5NMv9Q0wk8RD6FdeqwncWkU3LXlojPdiMz0016zwKe65Tka/0iILS
ETX4kNO6V226HYpoye5dl2sXXmOD4aPArHwfDohPDUEY8RuOrmAegd1LLT4fegHiqipGavzt+a4L
P+tWLWGZd4gKW8wVkBm64yCGJYEU7gQ2fNh7h+5leGHUHPFoM/WixFlDn6lkkQfrZg3GWUZnGIFK
SkVlZ1zcxoQ7i0+8aUdi4K9AOR+ozQF54x1AS+EkTR4PC9YYM58mzdFD72q9kLr4s6J1EGOnU2MO
sje32mnT9kHd1ol5ZceVACVBGORULJIjupRJgRnZRTQPVRsMwlzWcdjKT6nOE5/wS6PfWs18Rz9q
n/YoLGknzbmy3PO9nDVEHjEf2bnV5R/NRpgRzZ5Y7PWm6sv9HuGDHqiEoDHpOjwdf7kzHenCgpy7
ZD947ZhOo6eBNAw6k1TGoD+05GiH9WWqtTAN1HKdUUrgnCh7XPpBwlQvh6IaPQJUSszSHrjlADtu
ngclhQizaj6a8mGjh05seuorgZVUlGdv+omhM2Hvu4kWyo0kkGs9dSaWLYPXrHPMaOnyOIMuGvNN
777+aDLDKiL2vl2sPQzywFsr5e4FtjsMVjzMGvog0GCnM/ICSSnLit41qrqfT+IOCcsSFX6uIT1X
lPLykgcIAMBO9RVrxD/s62+Sz6DtwQF7w2m4tc8PER90DcsYC7qABaXU5MTDkaIoOXxXH3kJqYTz
5MG6ZuC+izU5W8xRtT5c02uKRRC2vLFnJTyNO4gCUo4CHFbHrHpSaWndx9uRhZzd1eISbR/8S39H
r2LxT9YFD24k29lQkErULnQ70EvDRI4i/6YpZLbvD93LTXuRdRTUSzpPRrjXETGyRPRcggkWWp0v
N6NXCfaFeDUl2DLHI4y0IGV6ztFhxFRjgbGvb5OLqHKk8rqBrQrbZP/Wn37+Vh370iReoosdUezV
CdSCkavGjQqHDmS89WNGHf+SnYDUOPkD3We7Yew7P/MnWNVs6R3VqvVMpD+tCkWcQGCA8MjdOrdY
8SJfT2Ji960r1TSbsQZG7QVJw2acuA1ms5oi7etlUqZ1lx6vK2J/lA4v5hFig76flsUiGTI8JgIo
pxOihHK3EY/h9LkqV4omHDOqiK8LVyP8LzOikYrxo5m3sdi1uV2wLYYEof2RHP9X72GNXxBix6u/
sRl/DjOVV2kLckOP9w3u/Yoplfe0NN9hKUYDNwPDW+KpjYEX4avyrlDxyr0nHJZjWHAchIQBZi9P
JxTugfsRf6Df3r/fFBZfHlH83g+Hr7KJlGH0VpkA4utmBKCv+8pJ08CWYcXOWTppljb68iYYrLFL
QmYlWYh8+jyR0Jwk4FATugfOWn4KK21eq3WTQGVXwZUetsD83tEjo2lF3MUfSz2xFJvo99eFgUw7
kPuW4xcj8VdVNZb7C6Xh3hCmRYElZcwgOtobYawqoedjINonFpxpNM+cvnmzih1gdkG9dsH8KTir
8pgC/D0Ps5GSFc/VzjwxVUTsyRWn/NjKKUu+kCIitY3cBlDPNqN5fI8r87imu/TekYSCRm9dlZTx
zkRXah0EwkLmwE+2XvInWgjsftdK/HfUmGmNpxcR1XgvHHzsewUpUqh+0sc8+dWDuYgm6pzrfrjt
PsQJ3eS4RbLIkC1QhATt9qb+vrJ44w8GcYrE2HNA46gPYLhUDUxwss3LbisknA1HFB+1nwPrXcA2
Ys/egiJykOhD5GySU1Msw+FX+QVzKFik7kpNMkhMraIlWzwsWdWUKW2N3kSn/GUPv/fKhABq+d8j
tr8wcWaAaLwheghkoLnNwS54oGhSMfukA0ksu3lXSCDnMUFEi//usNU/kawquM5F4i/YRxjWpbym
R5CORf3n2/L+ZAxsT0nqnvr8aMLV5WiaWRlLdcI6HXbW7OvPs8mH/9VcDEp1Hi6APmM2VXIDmVv/
hP8Zm9vFH0h5bHGEQkOHb1jyZ74mcRxt535A1CxAY0jm/bHEE4NR6dog+tERjuJKjv5wLUILoOSr
iU/VyadYGO6cj18hCoXXjlpXjcAGhKA/unW1t2vN89m63595vLlAuxADpcY7OAli+uV81l9SlhyJ
vSTv0d0Vq1fYRqGnreMS7SoewbldygPy2cGNFb39RlhHktXzKa9qL0XpVEnIJ1REZAh58ldQB3Nu
/brgHoEjrnL2GNmiKrphleBNoODbQSMW3Yg8mQogfW/3n4oX9CL+E991kx5Phx3OIP/+jgT83KF5
/DrQRtcBqCU+deqYSjpBoT0DZ6AF2RIRoSIgS/SnpUtUA+M3hsgoaaxilEbe2MDtDfrPYKtxQc/F
K8zpS+pcs8uCV5AFIfahOoYLs9Q2TB4Ja5e8DZzKNixvYenwXiIH6+4a+4iq2IpdbuVPrQK8nDe/
Xwmaq9ynquDLbGMPJCrTdq7PXWRvCRZ7d0fsSXasZNHxvCg/jGcpdPZ9Tp5wd1RGxjIDiBbElrP5
c0N2GUVXt6pzLiDnSUmYr+d5LxjWs7fEf63HktxUK3daCzAwTVO8QuR83zwdKuH6YiaECXJN/8If
G2VKQvuP4Gb4wWfEstsUefPMI9cRZTmv480ECRw3KjLzroA5O50gEjzvQ4RqJMujYbyqxtm+cZPe
f0EfafMazYjH+XxM7byrrqpmzolUzXWqImAjfM/jD+C9oDEcKh9CTCciI0R/8OPpaVq3II0fKleW
phVT5joaJkh1y+J2+Y7KWY8Qc7KmetcMYxzI6UeNq9fk4RbQHOTf9WX3ExY28Ck4YK7Fe/+FgDW7
JaFQvz/ReGYGjqHoCeF84JHzy347qOGHI/EJ1WtTAKUP34RG7a8CX324CCuoDQg1aHwBdjuX6cJd
vKbcvcW8JRB8EMHsHJflgXzZ8EFmzNyIN5iRfw/1gRERiTXLrXZfyUO/W01EVEamqz6nuAg2XAX2
tUTHTctBgQLYi2uCQW2Ad8vw+YoMgHQnQM1WgQvAqK7Gr4DSnJ5IaQkBsvGDiQMBAItYKMpORN2/
tcq42Y95qJ2eRmuhR84JRgG4/zyevOctX/KCO2vp4BjCfVxxlnNPa/ndRjLCszesIeNw0ZqbxYmK
H1xpakfYXJb3ZEtj+Av2mMqVxO25bAN+75gqttWJynZZGbUtZuwIVIC61rJL5w1YrjLQzgVThMwO
ZjQQEcq2cfoLNZcFRSWQSm5M+W3whz5Ay8OkyMFBAvxOkycIZG3J+Mi55rcpAx2ODBMXb7aTMQtn
ADkjKA7uYQ4151jiBvA5kw2eYZ8qTcohR/oevd0mZSj3u8hwdS2MmD4GbCTvdWMIhvSlFTM0+hzv
oxmGv/TU/t9vEwwr6D5VSwgDx8sBJf1IcgZV7sp31yhG/O+x7REKuWPSGgHN+VriIG8aS1z/Se1B
FIDVwNX6cA9DbIqZ3uJPfLFHHbQ9tWDTV4ph1wOViMau2ho2ej2EfVUsUycbo/cc6eSs+/uLDl+J
jn/fz2mw2CwFarAK49UNOAh9yCjMaeS1O7jc77HagB6iQq55pgPlD169gHx5uYNm+A25F7sYIlA4
UQz3+go6I3E8Qd5YV5ES0/RFy1iFqW6NKKKZrC/GG76o/ttDjHZ4WUFw3S3ZTwW9cPTBxkNdTnTn
txnJV6cCYR5FmPjuoKAyVrKI964fUP46HSGSv/BxB90xDHZH75nkTrGIflbl6Ku6gti+mdMqzE2i
c3dwSFC9da05ifjpe7xa2qQ9VHasvitJZoCaaoZwfaVf2e2XSdwmfrf+ug0aQCKs2tawlcKugbwt
5dUtCpU4fCJsbpbJYfr30s3qUTiW5BplJnFGJ7tBn+bcS70h+PQ0u5DHtm4eiPr3ZEVI8gBpwbgE
rkY/zTJwvAy/y83w5dZPrQqZ0+Q6Fgi55Wwht7MUmkcv0/UVtcengIl8L7iquHJjehKdniZDkCyS
ZBpkPxGKucHBCHWr5LM3zFYNaAC1CvpJMMcBFm861lt6TWuHCn/BjALik6zQK6uu6DXpJLqSssfn
9vCiLHJyy7RYbrl3Of2Q/QkT0bkRWxKOrzcoRVlEIHr3nA11LfzueXDD7AACjDt/lKHGsqvTBqLj
+AuA0bBPyYYFU6yhAgtXjZ6SgxwK6HQvIf48AYIM8Ken8MZ1YENLpS42nEvOO42SdOrD++N6/RnL
skHTGHC8+pmKNMB7LmQk8EPij8oSIxSXMmQ9e0uPQnSr+w5KtExQn47Ufu/3s2/OBs899xhyENf8
RGZbj73m3i3/bJ4j41AwcYy+hAxwsNqga+/209vBKd6oOmfkjk6sLDaum5Zhh8nvPNuF0hqWQiyH
T7qHyLITbUy/v7+Eo1O3BtmWktjEbZmxsjX/9LgU6AyZM0AEtuHijUK+WL+CpwE1QDkSLmRiCkDz
PWu8udZvsa8rwIYunIl5reSJzta6UDvemxYC2hxHPIw+Sg3aUEAWsxiIAB8V5CSv2VtJi41718mt
edHNdnHU1PbZh243SfMBLSK6THfb381M5xLQvahv83b1sxEOZRxoPAfsqeppr4K8sNWfhiz05hDr
IYOVMOp9wBi8RsNgWu4jNf8830Ai7r/9TjknCX9r90PsxJriy0agEprCONkDueNCe/GBAfl4HcN4
AfA2ky7QI0wtgJyZFCkSuWDzWlp9Ms1+r7hy4r7Pirhr2a+HOqU2GGmGJ49IGbWEkQsL3oFIAC2R
UM+h6R/I3AnKr/o07eXfd9h68HIn8TM8pkVU8S3SThsYAHSTNsNgS2ETOxGWHKsawXZ8A/C+n9W/
ysVouJBnoUqDxkVFKPkoDgyK8oWddEU7XVAwEKllK7MqfHWXl0fEGE6oS1QHAqQm+IFThgGcCZVX
O3AZVCh2HnfJ7PZKKwNfuUKPaKQxLiEBkp8JXbQzMKdbfdcZffYgmGjSFRuWZBFr1XbdpABakrN7
L3j4Kj2+0hK/DRqXVOcjiSry24VtrMKMoZngiWJY82hH9i7QHPCelSqIVN4YXXaadpK9wEmW475l
/XuZtxY+ILvDY8FSyM9BgUmmGoZBHvAWd+2XfTN9RD0AfNoz/2q5IiMyCUcrDutEygsMIVTBhTZZ
CgWnilEM2mVP/1wSXhpUycA1KXHCAUCTjyDNQCvqUqLpwC1O2OSxdHmGPj//vHioWph44T+E9KDy
uXyCCaifhDL8FOcKJBN+MXMMnFIKcF3q7xDFbSPyikT2xQxMk+TvxJ+Nw7aJ82rZZzgDmlVZnukC
IxOg3/cMflAKnNT4zWfHfSZ0PXEfB1w/2A98dpS43Ph6SFZDa6cUtnimtXc6cMDSle+Bq1P3sFpx
1psTzd+skycF63tv7ESbs/rhwV4BMklFsA0+rjY7D+kn8XF2VpQFL6xsAOd64QEzC7FZbzJOFg17
BXJKwjn1QvDyQ5hfzc51Wgx0QkvqG0Fo0QYQqNtyNvR15NJmGzLycwucnKyM+2hgVpswl+Ifkcx9
vHK+dCQitP44sonTWjb6eRjT2hyprDTZ9ov70SetNcncmeLrLuE0iD0mb0nZE49PR6+qMIMhz0Bx
D/VwULdRyZ00cmjMv9BVM8hWdi3vz3gefirsjXC/9sysV8siyo0gBaqS34MLU9lfwSP/g9TFj6j2
NzmL+veAwfjmZccjOSJyjOz9TrLWxyOvN3Bq01Bn2VGWCO229j9CubzlXazYLzBG8yF+EHUWeoZ9
8/73VqSw3L0bg+tFmBLNoef8P6vmCbW2SZPJ0OdTkMU/xXxJ8BEQp5PSlHyPmiYjxdr9GhryrXQM
X4A8TPajshHM3Wn5gStZjQF1DrMoBYJNrGT3fJx1zV+PnPb2naa7eRw542yjF4HwrFefBWf3IGZv
K5kojFLAnEhKlEqqk2xJ+LtGOeU6YBw8TGzy5krURASfnM5v9URPoPOfnhI2moXsUhUY2AF6IxYA
VeSbPAYMG5j35eWEnd8V5xKrJ6n+sbXEPpHDkMHtYwp8KaeK6U+fNummnG4Sl3AnYSuK/wu4CYQJ
zYKpIwWfOu8cKThESVvWSUOdbJnh1XR5hPYfBMvRnMOordVV6w2da6EhATM7I60w0xC9J44nCbwH
PYNHMeGL5T6mCjy2mT53S33ZjLaLPMmMXQuJyU2Snlk+5lDSmUsIfOlNNhtIiSLswjFqBvJMhOuK
pECsJ8V7EDzELNey+nX6p4VCbfb2cT5NpSbyAQoHnNcVSTlKTV2YYDNnVWmt0CYxIiAQni3AweMf
RCo+Pz5WN5JyUMWLrfEzQ6awwN92BkzKWZv+olmKNip6fAGaHXlLBCXTh/qS0DRdfpW96YzwjNoG
u56FR9qEpaAQyZdhuMXOI+9urRf7YzHOPBc+X5s2jz08xXbHR9j3jCL58C5/5SivDPUybmuYrF6P
g4wqTEYEaXn8Kls26naCQ3qswomtig9lh9m4UumzMO5HS9eibHrSit6TQbwl1wOKQIojaG28Wh61
1zr9BfMqqt88blGuf0xzEVDox4WhWkBkWyJXf1FGAY0bfbF6etXzzRwzoBloNHHumqUO3r0UFwM+
pZ99cIqW33g0PxTA7yOWtf0ra+QZP0FPo9rq9/MTEyCArhY+FscNWRO+D66aeq5HeI6p2iQmrm0J
zshn4DqNvCIitOpk+6yjaxfA8GgV4PxQmoUr7qMhjkO5Gb6UUsiOV/ftkqd3E09qp25hCgxN9hOr
9EOba0yocSfpF1DBMwPasoUXXznS+sOR4XIHQD+8XT5N8+tcWTnT45NbFI3puI9NqoQxRLtZDoSH
A9jEyfEnNwHS50D0z0Bpa/yQU+Y14VS7YEZrLfeulXpAdkUvAmIwk3QZIKqkUfQ8YY49+VfJPLaF
v731tAg4kL1FiFfNBTM5xgDUeD0goc4YkZNHrXjdycPngMF4/qFVZB8QQDqmq87w5X2Gwbb9N+KS
5U7LwmxQmcd7LxyZHFxal43fxqWwh8vnmnZ5Y5RyN4TOilv2a1nYJtBMbrO0SCd3+3sb1VXVRGUl
YexA58hKrNEpIGx1IgQRgivfamOkF8tnUAHFq/BwQRR4m2u5UwZEhAh+ULdJxOEAbigoyMfVPR6H
T2v6byEhFlue2K8gqdZarDW5dSUg+p1OqOSprPzyx41KsTISUXkBWsjcglUF6x33xQEf1q8oQOO6
G5GEOKUUUhswZJGYVQGGHdL1ZzSRmGtddoWVGQyYlZi8zbISKMEMNNdYZtalsEE29okJgapVtq+E
SopjMjUQezVarisMJ4eKq+bgzE05J/5+faTm5cUSkzs4hi90LtguyY0TP02UnJ/F66adCBPKKZJG
D1MXZSxqfVwdeE5/Zi8KAZNj1vbmME3IDQpXlFlMZw9NardMwxTg2y7pQRR90x9j4U/aXSxwghPM
oMIUeUxlweESx8V55Zeofec5oFCYSteM7SEjHiyjmKftDX2SnfruElSq1945PK3NRCI5FF4s+TCF
YxOcFsJEM8yvQGkcJ91cG5l7xynyXd2a6VzWgmIroD5ZaQzgTXQzHuZLgJVcT4mrtqielHTx7TdX
YCIOujn4KMifhqtLtCFLz8UodrCEok7Vohf4l7W1C7dnFg1aKUfmzOhi4puZc06KTTerxFrsJ58g
Y4n6vUeWLNZKgfj0zuFX8MuSPtGKfRaQDXZFy9qFhsBNSwpJu5bRVM9p/8LULLNOffkIy3dHfxEV
GprFblx7fL8xW8bL26VPwnPe9B0zIxl94Ow51SpMi4NsVCI+5jSnkdIIhbo9CoKQR7O4kLh82pni
9078gr5AaBQjnS1o69QEF8I1H5frOOQtANGYqgRN6o3dmGUvJNPhWrQyAP7iNeXQz4Y4J25auodG
DhhDAIaiQWY2jAegZ/4R9Uf5e5L5UVOizZenhe5MWHMt7kPt9ZX32fwNzVi31kx2GfKMEmezVunP
2m+mYjg2rfQiP0ma4RE5Sydgpe5dlOF+T6aKLF+2zAhCBP6kSvBgnVUn9UDcXVUZC/jYgD0AtcFY
5c9EDmYB4BZF+P8HsTJkz9MlyykH5kXmuG0kJsy9yIx74rhlnsiz6I6yhRtdSO6+eG9lgwePwNpa
UKP5gQ38F2ymB4IQXFjZVDWmTrUssrdcVr78+Drx7Efb4VSJbZdTd6RrFESTOpNjZgu6Nx+jrvBe
RASLwGVdyNkvKQgyO7K4cKWXu8IYhTGDogz6l5Jt4ZmDwfK5hHNBtNYAmkipKQFoxmD/5btFLX6y
9Zn+WKmfJ7gR1HI9nhwcrT5gTtOaiEeD9iLwApOwJ1A4kr56L5iYUOafVl0xx+xi8tWt9GmEB/Bu
OSDMTIkZ8bUKlCX2xya8y4nyxGYmjMfVMVErPtZkx5iyCyDTFrKp+zvh1/ETyMvZKs28F5RLUhaj
O9NOSDtXzeaCjpsDIJTMlck0my6D2BfiSsb4aad8E4sPQOgsDLVHfI70f86z7ygClPuuvpWjy+LN
36vbQ2stZ3k5Q9QcfTFy7U5pQT2NQbk0Xw9NnV+beck18QRv5DbiyNOq78T8T1HCOpSSS6B07JtM
ZSHkTxzcwm0N5bhJ8K8VOKZjz08KuWaICSSFNpgfEjWrScCvxaOCG5Ijz+fszbAXvEb1yKyny93E
lcbhBbRrjcOE+JGKCtq0a6RRSvn1VxVxWh8A2FEiBimi7SL/mw5SiYl0KjDoNhBddaC4axR7XnZ9
dTZ0N7ZDJjNbrfXvYkm8Ud8HQIaLF67A1XaaZM/KYm6+3K/dUKvPHRK/fLujD5AUHZKfYpVZ2au6
frtjGfKFfQduHtRs2iK0ooA1mjF4N5TrRZXGtLbNSdStA0cMB4eR4p6i79pE0tBvXIOx+U2xEq1f
o+EgZccoF62PN67RP5O/IXvEBIXXCQKRu1eeNA91wuKpwcjTqKxuqkho81MAjtJVuKSVnpqU9czh
pME/qqlUPJmR41XTWBy1xVuioL5N5t2w0LjAD6glI7PBoL8ayjh69JIDrmazZOjpVa512TS2ddpA
oBVdYowDaNrpCrWf/ME8Ji7bhekQk6jNSCUfKOLuYipwTymVyVsktfrM79/d0fbSHmr6eQDv8Prm
1xwC1zWF/aReqsSZ/ECcu4tJWUQueaN+XxSD+WYCNBT9OiPb5ln9EarG880LZ5TEznsb+YRFzgX7
OPwNIv0CX0KPeyD6vNAxq2rwm9HjveabTxU+h1wvrvZ6tokMFaVfXJTH2bQJSQrDGaHSVIPreQf/
eE1hNCtzUwHKQTjvBmzeuAZpJl15EgHCiUA4gtqqqJ5C2dHu6kfEt5SpizooyrXExuXuRPzH49VR
uphbsCKELSKaImOVUPuNc9FmZ/evTEMsDfaCnCfEQ3aGIpg81YsEeI7O0duAjDdWF0A6+dDrz4n1
T6+hQEWDqtVPWT1KI4y7J4TlAt+UPT7XuRtAaeieywSE2M2M2RFesYWoRPt4clnjM5ofyb76Igi9
TQzGYPEK4gV0A3wA2umJuKm6N0iCwemH3GPQGaZ+mqQCz09N8YqtBgbF2Y4nAc2oMGyO3X+QhdEV
eEmdmzxcRR8Voy1mGau2Tm3wVkz7LQvajkV9ivV+25DgyKKaO0+lR2n4f0pbociQ2HdqRwPfNtIo
/7n65dc8ifECxcVnXmnkPCQxSuHnRPxELDaoxwM5WvDz+LyC3f12bPtyk3OGQBd7Mza1XUxM5vqv
nYTnfku3tf2gQV9BmYSPgp6I6I8TL2csQsPW7BWdUIywDu80nsISDzeAOUeeRENntCBbh6b3njOb
xc7o1NnTCCG0+pUNgFxOfMeVc/3/+FrPR3q+fRmIpGDNUH3XlR6AWzLBglnnRLBBKJiibGdzcKFJ
vHZhy3Mpp3vFIq8xUNyhBJOxkKSzVkvU3ZMnEGZrz0xNTn3hEo6v4MnR+a83gZN2faU6bdblkeSH
MjQl0bRz9DKa7vPpUSb8AER0hoVa3hs3SbjTQDEEV/0pZGFt8uDe67WMMUl2oS/PanBhks9knt0v
VP/78eUy923x+SNwA87VdsIgCIZ6+kYcnrtuEEWdiWiogKiAmbkLxMGPZPnpFHN3x7ag3exspGgK
C3FlmXLoHZqAuj5Ik+udz1lsjJ2l1UcRy38lsXEyQOl+/irTpgX7lEZHlcb5vioi2tQnr9p+YMpK
qcS9JjM6/ESMtex89h9vsgDLteG20JJEUE8nGl+9aMk/Ih9+Ev4lvVcWWBcFPSQrbR7Y2jFIujNP
wjBhM8Pj+paKzKEWbzar28uNZYYtNJkC17/B2XjFfLeWiATB2b1vZdMVrzqD/RFyjIu6jgDx4MsR
1+aQxLzyMYnXL/2N5e1b0lnqs/nL06P7ewKxzp6lKkhVfzHXK1hB7qc3SAqvxwdIQwKL39F2xoDa
m4bSqGhzyBB01hdGajucvJ/fm+cwTknNOIPiBzr8OXFvPCiewWGGv5ChBunLHBBiEuxzdHJdazsH
o0ar6sPVs2e9j6IcHk6ljF3bTWs2X35E/uU0mTu/kttmFj97SxhJzStKlDk/awaesFvmZEl5RACj
DOE/aqug7zhhSjGYmN64vRBLslivKDhT9/vFKuJvBbGmzMBAMBydv3c0uQ0uC4o+TXoZtrDAuMsh
ZFFq6epx9uVgYMkhAps4tJKqZlHWVLwNUbsfrCkiuk126im1jWGNwbnPuTSk7cBQmAoIAGLlitlp
L9gMjshBhdopm7vODppXtYfIPCV6bk4Bib5UGR/JoGNayv+Wf0d1rx2JNwD8w+WL+ymwshfswJPd
Or2wSKJMWKLtc3tcC2cWhZ6602XFKBG8EjK80uB3AhGXMPpH97pX0d0ZlcbcdV5XWJsecRARj2Se
S9tmDKUJY7mt/ZBDhDmqefcwaJ8BllPqbQ2sa8m0L68f6TzdbVDzp0pPQsN9ZQ5NNfGXGJTgThcC
cMd5iWPuyOj/8IF0+5rlUJ185cpbgNxq9rwptZRHxl5swT6IrrjSUQ5CCEoy+XiZEbhN3u9559M+
IqE82KcueuIan39vY6EIzjSvtIjTxnHfsLx+67P9uxqoMTWOpMaZfMNWBwbmIlYu1Lq0lR1/P0SU
N9EQ0m806TvGQQCy+hMYQI0+oUnkr2SAFiUVTKr/ru22wjU/mc5KLA6lvRZXE5J14zCK9+nArbZg
hfcTZRsefbl6mwc87brAY/D1HVFyjmzAreJVXljk3IEn4N6W20V1EhB0CYXwrIL88RSj8SXJdFkj
bY/JG4c9zpFXM174Z/U8qP9meT7GQLkiMYkkEOyN/LZPCweSD0RyfqXAE+mBJ/yI8ZI7k+5G3TcH
WeYw4eKSOGGr0vYJYqI/33lCEsjKJprt/LBeJCyECXR834AcNd+u4IBGv4H8R2fBnVrkSmgvTwgR
HrZxLe2rKF0VwR22SsD8QziFtE+tIfI4S6Ph80vhFDSgBwNy0jtaib0FWjOs52omBdqBQuFA+Acu
uw3yLZKfF2hnMYahTdE+AyYYIXNOdAjaIKLUOnO2AHUlKxNAPn1EjQJ4UUhA3GQ7p3vWUAPY6yUG
3hzQdrCUKLR6QxgBGbNht7fDuMBXalWNVGMn9G7MfI1ehLs9NecUAWf5VUUE3Rc83XIoCL7VLdYr
+QLByV0/pPR4HTUggM2BZaLogv7pQRcsKuPxV51v4cZEdOUhRpm+erQh9QGhVT3pxSe57O3aC99z
lUn8QJGhlZbcsCYk/XUn1pR4VeMPSi9TcMJt26FwDekLsfCErWHSQ+C7j4qxoR+2ybfo2TDOMCM4
h5aBWFoj/jwIqsSRhllCWuBVBv3Zt5p0iIEk1neMBgD+ZxM5xNzgbKsti/aUMAD8I/0v1xvNM4CY
37i4Lj0p2Ja9ZOD7gdBDJI7kgF3itmnlcC3VI9Ms7o8nMQlFeLUMO6XeQ6S7ni6XU4VkbHCp+tQ3
SuTOky1omNZoeOvUwxiQ4JO6rzHAqablxuDof7T8EystzYRnUvFzkxF00B1zVUBlZ6ObDvYaJIf6
EftBL5xmIWh/SGymvJTT0+2n4byiq657MKMR1PJEPchi5ICrvCN9ywtAMx2S1ikS+6/0/a2iJ20g
Ydavmv3tHdr/pFlpqon84Sq5YSe8mRXVZb6zSisKCeLW+By+d/rDMG679n3+qX/HcfdiWXoUAGEe
GqS8j40P172hUNeSoAH1+36v0dEtxM5NV5d4zOXE/AlYtGbrDI+e9kncRVIooAZHJf8vSNUJSezw
ESf8m7bqKOOCb/BovHoCvDe7kpbMMqX4sjwqnY6+VkylImBCvLdVQIExDVLqbOK4f0m0oBEZdSB1
4nYGNZPaW8V4yKCkmHIIbHLIHZg5FCPGy1ok+swOY6/CnNkgNaApzOGkosTx9NNZNtq7MbxiFaXY
38/JACDMsJJMvMwb2K7IJjZHWVyVWHZ/cbMKEQtd49p72jdaNHlZDQR4lcI9u/CLmyqWQWohvLLL
L9eb7kaTuU75goSAyrvI1CqXdaeRZ5jNC08cnnWT7/oRTk0QYYGjLgGa2gG5e3dpkSZ3mmq3xkqS
5Aqt4lUIStB5Dsshy8OY1Rynx2FWunpJKCjUcoStUL4Smn8DU4XvQY7Vc4oUdlTUNn3j2MWJP5eu
ZanGADeU0DodJdOd2baNCS6WY9p69L8nKxLYlsEwmPnsIZygdkrE3Q4DXPHgEYqAoHjSGUNEkuVw
/Tbkb5vWZoaJgpLryQhT3+EwBitLMdMsJA7lsemBs6Lir0vsJIMMNchjWyeBmATqHnwRFOs1pSub
Df/Lm786cyqsasAei01L1ecrkdqQ04HdFOLLxX0K9USDW69COnO1PhfujqYW69VO7zCb3wwj4Fnv
7JQO9IiD517DWU4B1OQ6nzHThuYrNvCCcwGQt76lEPHp5nvD3Z3AYGph1oJeoKGWNqgvXMudKXwM
i78I3TLAQ7HtUo/UoV8Wa3PhoJJvvnX6Etxl9vzHc+bFPdPxsGUnkExl3D9YAvKHPjf08Fp0+2Ru
afS52RTINSZQgV5kvkbOnj6eBeiWDE/S005bZR770h9QHArF3+SmX6AMtYDsVutkSnpiUwu+xtCu
BWVaxwMSJaXo0cIkJAKAZ7xGBF5Q6lhraIvcacgj2WVFA7C3bYVl0fvYK9c6dTKvUb8f00ZlNTZt
GdSsBz386F58oIk+FV0+p4crGjnk4NDETeXtl+o/at4/CfL5aN4cJOf3xqHA0FXnK9vXetONyvet
w8PfGjqvCn+UPZXXfOX122TIHNBxSzfiX+jcVmS9P1vKl76xlAeytp6WHMla+RflTUbXn6+b2yPo
47dley0FSMbapqewFq2akjjwQXFd4CfVjQLoOML8UdEIZ8/U3IcQo5qFqs4qlmWkNFGbplb2HaY6
YrXsF4LPqp0wdoVhFMAuZkiun6eZ99dJPHIqXsLDh9GdVelxpIQGLPK//SKLcIIJhHCvrHsp9HjZ
PYrzTj1ISgaj4+8Wq6BQsFmaRoS8aF7qRs5Z9O7BbV8Ye+ZNfKHWmIDhqMfJUmrSy37WdN7Uc/cQ
eGiUvQSrQrTGmMYp7pbOkVGZy2CjnY6BkFCzI18icJWElZkdUVho+NHnVnmBpBgfqNnghS4kyaGx
P7XTwt3uXDjWP2WV7osAi6llChhrwxeNk9Bz1lsy5Ii8UQKgJhk/fr6MV/S6RHtRw0mqLP2fmSAh
mpRCsFOPUDUIgZ+ZaVn+GRoTVdWDHqzBxYRTxKdK49cfNWxXOneGyC0vweVaMBQjE1puqgt91fE0
qUOUy2b4eKURFNEM2XMr9NlyvjU0CsbjEzp+MmUISMYmw0tp64LXKGBgLuDQ2H9ydJnEA4XzOkrp
xDjymlBl5HRWo4wg3/lIEVmALHO0PGYdgL2D6vtyOPKaK8xaSwBsI2OjOMbvmIDIJwt29RQixiGb
3GvnIZc4GChV/at0Kf2RPICPuKCxiQ4GV+ZtqDXSvI/nHoby3ASLEwJyVYPyTCkJtz6uEPp15CpW
6AyE6q//ffRSRiKvz0XfnRxLwHBxr2LNF76p525xm7i3AnkgA4ANQf0ooVwSufWRmlP3CLY9hZYS
vgL29xBkVTX5ZRvEGf2q6GNUXL8Cvt3nQU56+KDWFVp1FJhhW6pJEySg0cqS4/iN04GaXULnxOTt
y11kk3XxN0eW6SrDa7FA3Z5RU6Bw+VARCvmCFBcCOEAosEKRxkw6/xMge4WdT8zhBBcNVUavClEc
if/GFEaS5NwE5jTJ6xqgtO9R3TvYyIoPx5ofxCxnEttnAOKLNgJiLyKP75zwi50o21A+zc5tbVm6
zzH+jrf1rwdBruD4dCo1eBsUcuFzV1R60Sry/gVUKOeiIc9kP3ZyijzMb75fDExqV/MQDXoFhSfM
38ylmHcEGS15GYx6ajSem+dzIrvbeMGExXoQMQijTBxs99M8z5OFImL+5pv/qD1RvBeNmhgHiz7n
E7bH2cmf9OBdrCpMl5hqquVhFplGVCAr6J8Rs8d9Ki5rSrwwN23Ew/eHufn1T+W2umwiBAIFA21C
pOpkYDBxrYHr7fYKwnDuYqZWZMDyYXxGKHtBKt4byidCn8qWjECznhK+bqN5A6Pb9+AWf8Rr3bKj
8Tmr31VdxsCdijEmVhyGr+uEeP3dhNfBcbB4IHiJKB/LpAR4TNce+6XONNQHW5bSC0ggzFvM7Dd7
/OzP52TYrUVZbCQgPrrs4lPcOqgqP7oh9EuVKjPZu2p9F7dF4cbEZXbjHagXpyQWRsJAH/3usi3W
SeMsKAvXqqkED9LRF57Tigxt0ycK4TXpFihkNoABwz+PZHWC1TnOdo6XnJ+k2+cdDSf5GQ0zn5c4
iVoBKH1ulfVD0gJw0uFfwMxdyzTtwny1ERXtbnLHiA5zfmdXByzuoom7ERPrDcUNsKIoRx+k81Tk
MTRxeyePHDMqLbUV+kWmuAr+9XCkQ7cpcv8BK03hEjeD+MaThJ5lgxLQPCCOaCQbJylJNtoQHxuT
bDqLb+acuyKZ7atKtH1tNP8mHKp2nYYCBpBcpOVkcs0lYXWkmwby2NT1P12HmNOcbS+KLmfQS7Mn
AZ0RSEAAKWYNIc7OzlAiaG0dXPu0joTAsUrJbDQPVtXeLDON5jOqoPPbfUL6ExDmKYyctGpofw78
PnbaGi9t9MdzrxPKaXax1DhOJzLsqJs19+aE5bTmVvmlF8iKpWhX+yQcJQc6mCyi1MXGfUlG9i9m
dolUjLus6+BPNFfEBdtz/FwqxwzfsdO93Kgwn1vkzdjZCGsJ0kvIHV/YgmXHBDq42TIol87blM8J
Bs1Grjxs9zwnRMRj2pneHqssBdRXJDYnyh2FGw14GOeU67ONZKlAcQi+4d5FbuFPEQNLp+7Pnvac
zskM6NPDV0a34Z65GPk62RAYoo3k2TIwZDdiC5nPY97lMx7FSTCAVHZ57i/ZhFBiLAKOABYaYX60
M567eVhEUvmg0pak69siwbi2PgtACbJVTdXh2zlid5mLxGe3OIcoW+QJaOCP0OU+b1qcIihYluqU
6aQ8b0yWHERDjPiuIw933GFSLiL1fax71Hb8kNuad/ZYwg6jAAzgNfb2wX7ygEmUONmZGXZF6iTf
6MXnVr/BroWzLr1MYBIyISTMIfsFp0ouwooMXWYq3XenUPc3M8URxXC0v7+/D/iT+mwSWue3P4I6
x5uJmQh6bZNryw/xwNuH6s1Tq0AV95zv7Wk+TfZrlNCEt0UGIYicPeaAYpnsXGScATpmsf8keMUS
lQHZKTsm44zP0G87biGMORZhiDzEw6aHt0utgTFXPfpVHO9jb3DdB1JeKHAgSBwod9T1hLPrF6RN
Q5cV7AEMk1PYTgkc4uErkv1RjwG5hC5n/zgxdFOQc+mhltKRezZi4IZaxsNUpTC7hKKusQnQ6z4c
nwL+kR8enNfvs783BA42dOgcl2jwgsjI25ReG/wYc3NMT4L2Kd1C1WerOp2nPPjIuK1jAs2pPGgQ
eGmqHa53Y6s5Zs2y0maiArBBTDeUyKgVazO57vQ8obq0Al2WCwGygR5XOVj6ZfAEdQr/qGkiMLTG
qjYmuBfhWCHtKUH46EZnJ11NEd7afkDi5QZsoWPlQEof+tVjtz2BtkJcf1mUOQHa0TP0P5iLOU5e
mKz6tbbv8qVir7nJyLwNWvy+a1dMPwfegQwesR/+wbR400ydXwBz0fGJ4oqFDyhE08hSAjNU6NwS
mIj9Jqnyjgpt7Ng+8Fx3ZXKoScZiXEMDVMAq9+3hXqT2HIvX5zZDsGjGOZ92c/IABBHjwqlxIaoR
GlKLWtnscX08dUiwTFGBp+hbpGB/r0TgNB4rJMUvoU0Np/t7MjSOtVKs5JD+H3RstmFAW4V4cljW
rQ/6NlOOMkyQW3U7rmjPGSmdSV+YPsiaPOerCPezhcuskJdlg4OrnEuIaav2ljlS87necE9Q4e25
/cNDDWqQt29x1sq86nExtO5Z9ICbLLF6Te+eIXHFdDSUHKWNQJAGIWOcw42fhcTdk2bexELXLn3F
Kq/CpGLPPtKbYCTLF5pF/p/B2kDJoa8r4+9WHvMfHe9LgtUvC8bZozcJlN+jIgf9AXYu0Vd3RlVY
ZEmXeE/zI6PcAKirOmV6uJHk9mnn0wTqkIaOT4eRcIWXF6nyc6wnrGlnuOde3Cjve/nslSWDIpNB
A7FLPOVSsTdyfRJNmomlA8f/YYBTNMbO3oloyQ2DpR2L9yYMTGfC6Doa3ZAAvKGmCFHwFqSUu/br
wSrRyMfM92/5mF38FcIv4ZzQ1FD2RD7mTZ7wErz0VBDTR7vVRxtesMNO8EPkMUV3+EmYsEXxKD4I
ta6ngZY1SFC++RIX0CC/7STb//CSgHF2+FNmd1fg/4IQRHDT0yHOhccFPa2IZWW+H3uoRu+U9u4j
U2yojxeozXSALjNAd70CiumXEoJszSfreSlRll44Dhgod89mPI+M0x3f95dhZTEjrIpMRP+CVu8J
nqPedPFXMpPdnq+JyMvZBWfwCjQbb9X9BDvDy+6T44bRgUlAaS+lNpt+h8d5s4Brg364NKk8jNfH
kOp626IvgH+YMbsDWSEdRRYX/EAv8Q+T+JskdKuf3UU0CaakHgsAOSpTA3HQRz4NMxQTx3BEDwSS
9kJjOhJcN3lKJgHTJXPAPpYlfclVj0uqC/NFEmpCP0Fm7geC9EvyUYSSYI/a2p4JLWCqjWsKv3zm
c/Yll2tEnDpN60SJr+SKifh5qfeV1ToE1elLfo34vPrll/hLsS07p4ZaCTYpKVZW/nBUlfXj9en+
HJywteYWzz7ASHN2nq+b56qvWnURHvaEUqMOHiO6YHfef8GAybakm1CY7jcFy0ojhUWy6F6Ij+Au
lY/tyff0gRCwJX+XIekOknY4JYQS2VV5p13RI3dXR/kEiVqDTWdskAYT4eTzNaRiI4jdj2rXjmxy
v7p12NxPbdNPOFnGsTqCoXhNy8pvPCwKkSGtE+dkN/rrm4U2TYCmq2O1TjIDAYPWx8oec7HtvWwy
8P4g1xS4FP1WgXjsXNtztFe2fpaPo3PmleMBT+jVs0fE7L7FC+oyzweaVW4P+PZc9luy0mylttt3
zwOD31vEGzbE8TM0AwZ83WaNgWrIrGYkBx6DosaV6vX/1BL8mJkCOZzWg/ad2vsKNh8z5MqO/RgR
LpSFzsPinB1wgNV/KIv2eEPGCIzgQWqJetPNZ1X7F0lifvfKypG49tyjBSoWbIbTfQwbFjA/BtA1
sZcp/qJB0aGN50EFim5XoCAS10ChnIrx5zXsWTvLl6nHp1JCz49cOXWI1qBp5XKI0L/HUWyC7/vD
zIekPtbxHoKzEqaA7jACAUyInJrxXWWL10CSeros1q5OJ8x6vZ9O/QTvR8aFa5FtvvjE+05mDt3T
7x3uImCrcIHOoY/MgERMdz1KIXbvmFm3USwhg+BYzqeA6/uu3OzFX/TnZb0xBLOZYoh6wWi/kU4f
glFt85p7EW8jpIN536wGn1DPjHsUPFE5N3Gx7INj0MV2fSqLS7xYh9XGS6+3LYkEEevzvwcHZtbC
6y/yUZftUBRC2Bu1G/uTTZcuFmCClQ2S/y/wvPIHvZ70grT2teafCxy2mcTT5Z8VPxop0ogTYWyP
w/7EQ6ntkx6vOqjnfiZ3CsA8N2hJ0BqsXTbjO0hjmx8ATq+wKDJVQ27k096eBn3/GqoOy27bogtG
9smJeyETqzbNDozBZUyTIY8YcyDhyqUSA1cqOli/ML9qkh1y5xxiik+3VdBzo2rXqD3PwBuXwcUY
Fv11NEj8WP0ZdgYpAeL462xHiikqkx0VeQI96yqgdaJI8pvJR58Frl99AE0zmUUHFG62x0fOT94y
ZvxNwHTFRnqVjSus+3Pa44+CiMYrVdx8l3KatGdMHhlrqXAeEzid2YiV2wVIgkTqkvVFAQSpRd5q
UxJzbOSW5WxI8J1XqBkwv3ku5MLEbIo7RErvHZXYRsmuq58Tcb/F1/77+7umvR8vXOr7JUpDwOs7
nIch7Mhyl+yYZ8eE0kqZgQ7T7yUeTVVD1OyX+VfaWFtqT1oHjXBJPxsfgii3hVNJ4UEfetrfPeLG
BqiCSTSxt311142PSPmSbQyGv9i9lhg5Tb2qiEGVdcgMjKyTHyk5vj3zmDuT7UqC0xjfiDMs0C+U
Porh9PLEURolLxRU+0uzHoXJX7xe8cvqDsOZ9iAq1gNOquxHwzYrPD9KanRNR1pdXd5tFfYJcwHJ
1YAFfM+WhbK5NybhYJLaWN+PqUEWfNAUo0z8IPza3uYDmTAMyPG3B6Wv15Uwy06ZWbarQ3XsPECb
jASiUOQc33/jUVLL2ZWf+Sbur42k7StQ1NcXlVmU3rB0cb9yJoKhlErEF4Z5vQlYk4umR4WfW+LV
0cqBhImUIZmwUA9fj62M6p5Io7vnWd4XD0ccyYXafg8m3/cilCMqIJuA9VUKwzCOWHZ3Uz+fz+7E
P960YpC9TKaf2uBkjUuHS8SEjCfIWVQsZeJKySVLEe71Js6bnC7eZGZVtv2VTRs1vA9WW+b4MVw2
EGpkJEZXzduPnis+J3CQFgLHOu/mLB5sQiJJ54oJp7IzcbFKfMdzvTlhG5e/qduZLjvSfP5y4Cxa
eVmyE9sDW9nGIxebTvqM2SypV0AyBUr4/4NgQAMfgO0wmqMrTRa7S52lAr894MhEmQLvJ/aboj9Q
yd6TAzuNRLAjtrm+zbg4y/SQf4IUyl7eubJJ0U4BIK4yPyjosmZDsBjb+Wh1Gn1LoHh3BQeAftn6
Jfi4KKqx2t8XNgOdqkQXOw32YJ6AqphcJ10W1bttqzO7gK3Mn+polLd+R206/rifaXgyfJ/J9j8f
dwr6S6/7yJ+OTMw4WirAJTEiRylAh8x60PFewePLelTdXt7VMxMPHBtlUlfikSMkPHGGu0WPMUpj
bQd8tGrv0x/xsmvzOsp8CSR9hkyEcy2kxTvYOqvHpY6d51VeIXsijEJyT6oqBX1Jos8o7KaUfcJ4
91nI9XKh/Y3y+arJmuKs5+pBXPXPOkY2fv4/DdnEJlVQsnAPdD8JZdz3fzBZS3OlDEfyfUuxWaYm
BFXadYDPeuWqcIhXkgzr0IZ1XYBOVoj0eIIXQK9KrUnKSSl845/b/R3ORN1blNwWBuZXhFMcFJiw
8GVNfz+4ZBAP7WbRsrEATwIsMZxkD1GbA9XIr6NyCDnNfnRVYyAzu8FW1Y4bqDhuJfTlStFCLdMI
NFZqLLbmSa/rQX8ztMqngQyes/G3tSr5Df2oCNcUhVoyGh2/H69UvCJ1K3BvZknBwv/Wf1clmaya
htd21fcFIwmG9Z2LJJhJ0JUAwds8NVK7QxJnTe5Nojj6tezbWuhyFoWlFQe8LHN+ADIFAabcp42i
GRpRIKocOUa03Q+jS0eF1DWEBdnjOn8z5nj8dNdve4oE9vcIY6GHHY0FDQoeRCBEuqLRtRRcp5UD
SpWEdpbh5DQCjKsjvLdgpKrVTA+4evuUgJHRf8BHZgTPf+VzX8xXw39/kIIISNhdqi2ZS+JpBxRa
bKNTzmLgRngCEwKD+F8OOGgNsW0kD3xR2RA6WtOPWLJ/PoayLmCufmPNy8uAgC//XGTGLk7DCJnq
ClSWxlsIljDr7OgmVgwLipMhgovL6B4A3b9mEoL0e0FBJkq+RaH1l5Tch7gxs6/ohHr1SnRiEWtq
R2UYQSYUuINeOfv/PxSHZdTadydqwf+HBjp1EtLmEo6JRCBGw2rMKPwnN7abIK/0F5vjdHfaLAio
9NubxcPBh4CJQc88HM3YjcAgJdG8J3XOg1f0q294tL4ynR8MhPqJ/sfzXTCvYRb2xFUfwNb5P0im
foOJ+EpjBeHWeBmAXlnO52By9Bdy32Q+rCXLf0tDXLV+CiAHdbmjVTw6fEoJEtzJ+62gU8YlTFQP
KX921SWuGGB4Sy1VXwJcPJipWm7WlG7NZGwFTelQyPDzSdEtQJ6MbqDWW7IcLYhWyUcZxCJ72OWN
4Cf3Ypjyq4eEjpzATrxNctG0kwM27j6xqRGHi+Tubm9FUiQ1Sgc4iSmIrWuE+UF+/wQq7/fu1p7o
Q0QjVogj2toohwthuESOkts9vfU/K0ewixfOQBfJyRILxNqGYhxFQQgmIVTKqwjcfgB9/f003Ck3
4+JynT10KcE4GsWUkweS/Qq7R1rn1O33rrqb97qjvuTtw1m11gxnZEy6HWfSBT0BGxTvYaovhGd8
LPauR8tM77zfwwli17hgMVvtVTuYg9+15XrOEf/Cb7g4qcaRFuG0YRZze1Ma2iUJPniFfBsowcVO
C/5q/C8eTzhnqiXYdPF4+R1TBmn4o22bOTsGbbISeS/Vto6o3z63i7nJ15xaXwgv1FEw3mFMeBEn
sWBWurg4a/cO1qSPLc6jNast/z0xe1eo9SvkI7NzvlehtehKfOq02NlfHlqWMmRWDremYBsqzfeW
9T+CZKyhAT9MK6R3/XjCHDknh5sqfXVWmN6d8DavE0qEnEBbdFabyWEa3unVZCPSxe45WF1jMiDf
nrAK3qBXKdSjseXOXolR5evGBC4uerJSwqYTpkhLG2JT0dUASvphg87ILtm7NJoORNmobfYDL+sj
dI+BXfah5SRuf9ZXh87BCtQnpTvL4zMxBKnw7tbcybLL7TlKuHdct55qdVhOJIhsacEK5mtYdOKK
PkUqZhtuofFw8vFz2vPoFSl24M/24vaTdkLKMMhIzZXEQuJVGmQ1ov3/RwcpQZ32MS8y9Q74cekG
PuakZe7/lArlraOh9UUvbp4kKFTNQDzNU5FmaLxk9u9PqyPxQgM+4w7IHXC+1tg5H33zbPl05F8Q
4qNKkCTKYPkYnsS7dm1wKZSx6wj8nfaCSFoEX6EIBnT1yr6D957UKmpsoY0bkwaI3oh/IYuH19Ay
htXzf6qCy/zYPjl0dTAnxiRQxvgjMsSRX/IT/lgF3aN6LVdiHEm3PvdUwQRLOdoBBHhhH9aJT50p
KqLT5e2/RI8bJWgDVaWY8qprgGaOJFlGwEtCZW4urIRiFOrN5aZYD//oYr9/WvsA2ZhK5Dok0tME
WJvU6jgg8fNUTOGGb+dFOZJe25yi32mXcZBppTAnNynjReRuDFquxb53+hIToZmmtEqJrRXJomUn
gtCfU+4j7OBmwj3OshtLawoYpqC8PRY/+LnaNBaVJl3pvUCCREsSgvVUJZQApfAXrMOgZAeHPE/4
shhPciMSKvmbRqYkCurnKuRY/ojTo7ybchO4GkaguNEGQyx3HwwXL9aKLBZTav/FcUYf91/JzP61
SKBXEw3zf44kANMavAQnWFSAqU8Iby5uP7lJuMvuNRoSwbT4OfvA1/uHUjzxfPbwsMujsEf0rnos
O6D62uGGYf+KBnkuhK9y0xJljSYPkWmsdJPypYSCEn4AmSdoNctkdo/YqDFEhNEHhWi1PDoET+0l
NjHwHM877tgH8gJyFzTAzKrpAqfd1EtLvMhURLq4+MP3jHSkQPohHmfZ7g58Gtwvil7q0M30rDdD
A1T4KPk8yppORsiMBfGGKCVctXnCYk5o8XvWivNCmA9HpYwJeSQrVClbHC7eBoDj/RJE4LrHeUyU
2MSp/G+9MZjH1TEcftPWlltxwC5knQK7NvuPMF9bKCuvDhUexKJSI1hwRYPAWfjBaCoTEZNPYyeM
k4HkTLghaLcQvOuuLPGVNhhWK+kzW0KdIBjqKoIy4Ks3SynY4muEQ82KVKvcqx9zVj5idO+btWKa
H1VoQZb1UUKBw3avn1phi4Kmwmw/CcxpXK5UevavHYOaooFs3RonRzMS3HIfP7WfGU1WsDOVx/ag
N4qXEOcx+zm9SZ27U5ZdD1IUfN+xKE7qDmZVDLdF6XQJSD9sNDWTCcHBwMHIx3ByoY53TWnyXKxj
owoth0zHz57H3vI3iAWPSuwLj2g94lpmE8n3awwI7jbxGWmC4QtpN0RtTXwqoPNm3rKhyIec8gqF
FC5Vd6MZ1lX67nL13xfkwQJk4zulKlst2y4WTU2unSUyyszb/OHVhcAiblY9xb2JSSAGzfAtkE8v
0A6eEbHsHa6wMz2Rqh/+2mLBdwD37oAvhmHvB6ntzUiLs99W6tx5QJsBLcmA7stBDqvOkq21upiU
x54eemiUTuryK5zSW/FK+4AlkYX3w6ESBeIYNhohQfwLUhfDhBkS6qSE73gt0nho7qDKfFAdPsJk
n2zJpgG2ooYpQeIx031QERgTUUMlRZ1xFrigOwgajYUrSqGuIrIsbzVuopCfQpnNg2SvQWncHGaU
rpIJAeXem4Uv8+jUz6cER7EvyajwTLxJFavQx2aNebb6IHUa59LxgPIdYskHtGB66vJJYiUSR6Ua
ajfWYSpkKBvEQkr2TXbpLuuig7bPK9fXFnqahuoPk6gLrugQqIwanim2K1h7qnHWfX/C69m1R5yy
gBK1SnGtSYX7DRYIBwBtmv3+zomaDp1fRAvDTh94vegJrRK51Nfts6uyjLrcDaT8Z29FqUcHAKd4
1RK86K6pfqKF3+sQeMaZFDzdKcYB6n2sUxTX3GKMGWn8iOXSn7JHk3KArCbG6KYMZhfHMAkQM2Hq
bcXClsDxt0nMHflbaNOW0mslL/r7+hioYqHOCoOUTX4Ub5s1jkd/Qhlu1n+Y0fhAM8aQOdmZb5CI
Ore9TxnHHyZ/pMaHtA+neUpl6OU8Z3Ui1j8VEMor/a3LtqwrtWzLj2XuUgwItQuXcC8OBMYkiUPA
UCnqQtbpzNlatgNtn/4sQ3ZInAuWXJ8d2tX9ZElbhLPePjmMxtyEIOhxBFs9O1EeqL8vEr25h+zs
xUqeLxsoFWyPDd9aQt9CA/pfa+TE5FqXucGHJtGFWGze/dxh6/11GIgelHA1zuDIUcjTvoaVRMbu
WOoyu2lmC0PqdIZGioXvNS7HdO+j+5bFxe+u58Dwr25HKMVuEj6ijE/hzn5Rm33D61DzcKgo/bXJ
pbDQFvuKthAXmqXW5TbgmdWxCCkhLl9PMpSB/9lf18PECG4tiMW0cRjJ95o6UIeg1oubGcK6EFfx
RW2wtHzqBLJgu9zA4CT63t8vrlfR7NR5vksmJQtIvPFICDhrKeaA0Y5mf7onR5vtvK8d4XASsumJ
8NPFbWdNR6pIvwLAZ3GqBLxA7tdl5rom19GyhoHI+4RuH8w/VNRan1luoPjEnX4bt9KR+/bhbWBx
iF+FyWf8lbtrvPy3aF3XAt6XUP7bRz0aLwTTveXrjnNBtYi5o2jFFcp8twtlJiwOMz3sooQZgCBg
5a5eABj76B/sU7DJlHnBhKH/Uxko4znkx3kcnBGpigkCFm0v39lP8Cdp3PFnPtxifmBpXet9X0xV
8+GhmH3kGclclbRLm7l6qB67nazirTYmjDkwQztZX6EhsFyXHv6jWVuJPMUkplV6iBZjeJYrdDw5
PBhudKPaHYHWql21EwqQ3kaY5mvuXp4P79OFOLnzspnh/t6jnsD+a3dAaSgefP9yeiqh3panp/mw
Hn+RBV3VBn0DOsDJy5zvyBwQa0Xj48YoS7PP0mRRb8bfh//QA5oG9NNAjQj7sAwQZMr2jyOmu7PS
k90hz+4GdZR9vHMefs7HoEOVdrV0Zk6I0xJlUH8G2txFPE21xTXy/POId5Dh5g033Eegb+JH+Bbd
ROQDBxHmidZxIX6gT+Vtx7FfxBJEjzfLxYEiYkH22aWt1/gdd/8UfUxaD7Pn/jsIBlVljaGRb6ug
MWtUON2Mif0c/QLj1c5iddFBMt5vzgvr2/fNYGCHemO6VrsXtY5LRjEyRo2/u2MRpXHSHxitf6t/
abyBigQgzb+OGgEzjLL/lrOFLHRmXXaKMbiA8p7Z2DYrOuOFJJqWrqVKadzQdgsLOdVACot3uRmw
yUegWSqCbVaoy3TkStDqUOySW9yRusbUTrqEL8UE/EhnXeEzWqtcUZrDg6AjpzNuQs15Qt69E6Ks
f2W54iYa6RibKlEAtJuhuwuY0yDv5o1dJ/6W69NoVSraH2qEmiruZeA7mKLuXQEbUhv2vof9EUi6
rVMshyCW7iCT0dwP6329hpFW3gPXcYF58B5xgAwxHPpKQwrqks+4EAoHPp5ZkIKbM6zcx7Q+W8rm
tJwKHcHIE1uELWwVpqny/onkFmZcV2YjLTroRowohvGcktM/XoMKEwemFtyBeSC7Mkzzgzgz/3GT
n6CDA/IcVn4n7zBxZEcEdnKWdxAc8+RNr2FHGvxByLB+szDKscRVfSNE0m7Cl1fuRLn9mhus5he9
5/CXtp+AB9+sbqurkYA6BFlRLtXsWkozWThTwxegJQvPPuausqBRc9u+vEQPpu7WUOgEG0k4qIyd
HdhJHV5Mf4KWBiPWyAUFDg8lv5hK0wbprhz9DRSYwdNJcNrrxwpkuI3WM7yuarChVWfAxd2HvGa3
z9KVO2ZM8YhTp1H0gb47tIyQZAVxSR+GIhUpn4jO2eCuGLRwZSL3/z68rbo6j4OFhSCAWY5OHVDc
XPD7tg0eLYuheA5KOnClzaqH2rYjaJsn0PWRsRKhLFmfcVU11e9qoKeIHQlwrQebh8XNCsvyFcEh
8zJDv/zVXfLlvCUpUmPkEqpy/xdXsCsaa9WIbiyanfm3vk+6QAZsNLrn2FhYU/4AZ+Y0NdcQRuXy
xtDrkTj+yfMqzalzKLOMRy03yU8blOCpQWTO+ni0C+W30r09E1QLC4k7r8CJ//r33evgO/CkmTJ8
Vn/VU9aXvVJ/f3XvwTlFJ7rs9+SHAkziAwrfc5yL6nBwJ0IlTf3JmMAQxYaJr0lCTl3TNLTJvqLv
U0tphVA4iYQbPgUPFpzaasJv4B7fmDZnEoyZ9ilUeIS89wMr6dPRJg8aqKQlalBmDfZF2TSVmV1z
kFRts2lT3plWJ5ADvFsujHeIoZ2n1d+5mZJn55ighB0vW91Snyvg2BX8JWs+kLocPwtf2WolbJiA
G2deyTy0fgWbFcCs5urURkJHphls3mU5Z2Af84DY5f6kAztKgs79/F7hyHQ8dpK5BhbX7C20Geli
iPlaw74wzAZg2HbYv/oTap4FDhFEJ0ONxh6rqwghN8mAlNlqmRjoZwQ3LZNfeC5O2BLcSQnLFcAr
uJ34IZaWQgO436rciYo9EpSzoucRWQEdaLXu9SGg64MrY+xltTiKF5hg+4l1GygXXOkpbyOcOjei
Ef9wwkjhPcUzBsor8hKf+5unKmZ1uhUHO7/I+0e1veKnXHUDqmEXYx+443epblE/lZDcCVSWaiyl
r4E7EbbZWncV812Qpu7tTM3bEpG0caEdpfIFB2I6rvST0Rctme3VTxreld083CAbf7hLMv32iwfJ
Q4tSXwmYnOfbf8QakO3LJ1wVy3Bw9Sgp08WIp8Hl6YWRDqsGVtg/nvoJrGkah8ceT2XhGZXvNasE
IafURstfblHOnPhs2UYaUk+kwYNaWZUyybHP8EayjjRl02aArVXPfAqs3/ZlDY/NPdizVGNyBLSv
qipsRZD3pE3tq8SLjWNFPGra6d1y17tu3zTXUzrcGvHKF9YJoS/9Octhbbpb3L/hakfwYA0WwUJ0
upylXGyLMAIVQIvN9p7npG61/S3mL68yjFXdltPclcsKXbw+WkzAsBs8DtQbBEcWYYc/OWf0JF//
SiNycdEQCO5vmQGz0vA3NDP8nSeS8Y+XJDGZXuvNEjRNNZkxEJaXCaXuowvhuy6knVtJnYL+mGny
BIjqz/eZzGYpv1ZBBzIYnbfdXRO7pMz9Ef5yfxmfDgLW6Q3+H/hyu21OPUQwGSqNK++iPED8XH+y
suCoTTXDbmv/+LkntsyYFncFzoulS4p9+mi0HkcSJXmKkfe53N23uy4fO3F/C5wLT+d9+QeYRnpp
RsFTd7yxYjO2TKFCT8WlKwmG5uAGdfTSqhkT8njSZLL9MSvoG0SHiaY5kehd7o9a8U2lGe7V9dEy
G2lY3KuREnNwJAO7cwcPhoXlDUfBmakmpp7qvQ45u57hjQcahiWM7E2KAyaSeM+mBohPNmhICi0u
P/mrNSGKuIYbCTBSVvHgg3n16cJHAsOX6PPFs9ETlx8TrpIMM/4Dib8CKb915T5KzIOB2473ULGD
ywuOuLpi5qMG6kIKf3251ZblXOUZpU0cctsVDoiR4cNCHsHSonrYu81at/+DXsXcUXCfRNTIBXY9
UoFnXW9ztTKvIJCK26fRPxqEBYrBwyo9NZhos86azxSf0a5SHpQuqvbnr+zBuYCPu6+a19Gb8FKL
zMRduOcGjaDjEQ1IYiQPmAoH0CTw7HUrvQH6NO1oF/wntqH3dGF9uYtT7RcWeQZF8BfPlXvtLg9M
nYJEn13i5g3ErWTEvgqCug0ccpMxz11xfN7c0f6jl2jSGVmwMTtfLILwD07jdl5bsS8AuHTqd8YQ
T7nBfheEzaMSQLFm1Djc0JnrF5pqGbPekcr9bhMqeSPZBwuOFaIEedYro8sJ4TQzSfhMgssUttCJ
peAki7XiB/h0G0r2FwzF2nKDAxvgzC6J0z+muzQEqmv3CHU1F6hXvV+YAeVCkqrXXjYxhCBo0x5K
OnTrEeOHUtjNTmcfxo88J+TgIR4G8RQ8OKb29hDUWOkE72Wnmoljm41fsE6FE/HBSJ61a92zTY/w
Qk15ZulGkBl8hL4XBuJhjFepqHBwByXD2YjD/i0ay9WQD5HZ1ElvuJamxFxCyUsabgmY2WX9heWc
cOqip9hDniQEXxFZvkPwI3SxzjnFKMfkvTglYjJLzvQibD6QqfhEb6yW8eK2AE2cz9TYBF6jLcJv
rw9ZGoDYpPv5xqRO+Zb5ik5GP8igsLN7sEUPxSYgPbidkk7zMvKp6FhYpDYZUay6wyIKZ0fkV/dz
C1M7dohKuIh87ek0Trmo+u1mizInmwYyAWJlrTHRh2NxZ6q9+VSXslPPhQLO9H8ihX1VPpHcfmDX
q1Ms9vaDfBtAQ9pFsyDaKqjeaiAFmsqdBRvlWdi2ZHghY5hzi6M5syDwyt8jKeAQ3Upkll6RzFq/
Ybwv3Xfm7VbC9f4RicmdvsmL7x+fPaQwECXfW7Q+u8N+GdOIc11XszGMDDhFx1ZlHYPcDeiDEVn2
FGckvlIpztm/2W5tXhPUvMAHX+euz3T/Ufyh/ZRy0FWsREuD2d4RdXsdv/g1+oQiaP41YOmdUAL0
UUEApQmfoKaZqhK8453c/0SglXiaqGvUrjxK+QBtITjtePcigy8/6NPlQoU8jtJnqd0cSWMIAYsn
c67W2/++idc1oYNpjGptsH2MVM2g57FgGNNa+X0lQxcbrJ3cD9zkttfcDaXZyHuB3JyVBkjqsW57
MqQIH5daIP9l7/vaZ9EJBm/rMIuJx18YojuHZzrEnilIjn0LnrEtOZJ4fdO1Duk7px8KkXrAU/hi
IE6OcpIz3NyctUAY8tbWDvOxUJELKQaQJxK1ns/zzPeoeHjbw+vnx+PLzbl69C13H2TXAlnKF9b9
ODsiVQG6WKP00zde8ZfgPYStL+M6KErxgPaFs6MLo6ktS4uFrPCimzgPkOm48cNdO65RhSY+x2fr
QKY6KXSArkV9skhlwI5KgH/QEuqnUHKKvxh2jsZpNhsPQI1/m9pH/0g3bXbKpzmHCsJWaMzARhWq
XqwwYryGAiUXPjAcpXP9p5J0SsaPADCTMmZGSIXAHuF9OKB6gUpQxA4k/xHzTUG8OC3S08WTOnc/
gGmsFOE93L+Side2kV8Dtse0UPCTDpYbGH/MuSPt3e3QlT3wCdDDEFB90VoUHhnct6MZXYVItQA+
G2ckAigRR8GqzdD27oZCKsXVvX0OShQs+THY0zLG0fvDxPZ4n/3Mweo6BOmLAqesrnRYAm/Q6qh6
cynV5Zhd2oNOUv5wI4hdD/N4MaHHPxn5037EieA/4pPtR3kZUJHf+3xrtXmiOhMPVK/4KF9TJu0R
KVjukVm13LpWRLPsVDMwtteBlRjVbShCRpNItVDB50bqupo3xNz96zFoUdCFmYD+cOfHyFTgMu0t
IyfQZrU9XYyk+dpJXFlP6NxvnDVuBBnNlpF40WdWY2kOx6twehE1SVYvY1DSW6rUJRHHkIJXm2b7
dKAQ/0UZ0RgrNtMPrzlxV694QD9FICaTuFpIpZlaWLOHieQ3SdZ4yuSncO6KLvCE5GwyxVOlpMp4
mq95WgQIsniYisAY5oQcyEWXb3sqmCWWEW2BtuXyUeH65Zvtqf12Lv3PXfN+SDCpIOVr1bfrcgaA
ZqVAywFkmcP2F2rW4p6ZM7YkbbeDEXrB1BlbzjuAVNZ/zYwxzTgLHpV2uI2iRJz82PjqUyeLLg+6
6AEg8fGWJKQuN8OnyVfvuWHQsQ7N9v2pCCP8ZjKS+9vHqSYpl1Cpb48XgQ1MW4tXwhCzbIwuAGXt
L4a42zB0FUGBkUr6gi9LNDjmyAwyEDtmcJ4F3w7u5CRz67qQ8qWGUnSGBVnbQqJngeq01wVor24Q
MLo+A3+zIPNRyIt+r10Ns0uCfso9vDmJMlNvtIJjhCqD+3cDxiF+yPBsKNzaNv6+xxLrFuszUR1I
HFnm1JLvIwYLCbfljU3kzBtZEYeTNuSpnK6MJYE+3DijmnC98f3s1cfszpDt5+YMX5P/W6xml7IG
US2RemCe+U+oLpckNxa4EyGqq+yhV4qtRCJLS/fckBFvUsaIWJ1GxEg+j4x6qpK1nF/PVG6Lbc+c
4tTWfw/69a0HBEe8c0AEQMFVlBR/L6DzIepoD/uoBQWMCoN78D4cb51Xje0eLZHTLSZq34CN2BiD
sgMBrJf9ViaYqhetVfe5du4B/vD8Pp4pTd3+GTk8L5IB6rnlybx4IcGmI1rPRmdjJXe+z149cOVP
8hi8IKMKSwtjNZTrwsPciXweBqcvsf4KvzthlBpuZYQt6BGJnlXtzitlmiTrgUw1x3C9dEHZ8twO
aHo5MmFMvgD8x6BRmvcjpFmYleftAerawEBMufTR9DM5BsV1w12qVSAQyaLfSph5aXrV+v9C254w
H/kKJvAGvT48d0x/CfEMY9o4QH5f/TPOKSb7kHSih3dpsGDQmpmo/9UDzGYojsLhIVBFfu1ApvzX
gFPPmqfnHVwIuHRPVevijvwJyXWttgmJeOa5ml1J2efoGth50tslwLhsCJ54oRoOgS6VxwSK8jwD
dX4gbecACzq7YFy0yFrvTBbfyXX1+sONs80IllHjyNFWfhOzl7gDFCBx7MhbaMjURLyFvzznzW2w
AxHpNtm4bNmuwtL1Qh9zzI0VT+vFsoDHf1dsAFWHl6SYQ3aK7RyWJIfFXi6zRvheBYtXkTNapYUF
IYH9U/NKA46KGuYIZH6QR/7aKqZ/9UBmNwEC08Mqk147O3Odxl9TuvUNDKnD42DH/D10gxskoGg9
NTKGZ0Ka171He74I2TEp2+vJN8BD2DK1yM/bCn3t7+lYpQtn7+k2VkliL+FKGC8HMQhv168V8JAv
DhQKQZTMyp9FlcoPqcHpOu5KfhyInbx5fA1icgr6cdNF6EbBPxY62Z7qxOyPPb3k9NoHpr4CvxDM
ue0oz7KmCamCElaAUuqM0SqtNxMc7u8qUlPyVbk0p+HQ/jNZCHqjasQ47xTYMTuYrVCiCr/4hJNz
DirH+VpNI9PJmS+GYd6r1er3X0t3sWJIztvjnciEepJsgtebZfcCVYpEQ3ylJhNlCfzorryAvVsQ
c/0EbRhQoY0Rmy49TSZfV+N+7mszwChdNB780LW6GpLo7km1klL/OmFgoAdMXuqfhU9aSyPV1Acs
J3EZA15bJdEdooVhTUUur5rLTGQ7Img/KHGkL04JGAWZY73Kl6jXBL0HvXSF3wB3vj8LE+qfZhvR
WiRTGf/2f8qeIGvfJ4V5ea8+RycU89SYQd37ncpqTa6hxj1tkXESeH/7KX4yOfy7/z17nhvwBZLz
X0envA1DiqA2N1B2mywsloNQ91I5CQ3TptXR46z+mK2ZyxUHNg520KTDuGliR+H3DKdXLtwWwZKy
X1rET7HlVcjIxtFHsCG/je2vvahvowtTdWBmx9v308ASaZNJ877Tah1EGCuO1tSTPoucEwtsz21y
VWWOp+dSnqZyESnTR5wVtUho+OMZPg7IrxCRCktPlA7nV+vInY01y7b8ZU8Gnb3tKpboG01RE8MH
RGfbOl7e7QpGdEX1XzMH7GVwYp9nQDkesrt0BHaoRfSQftiNgXrsBNSH4wXZk86Lj8/Mai+O9x9k
tSQx/d+43HPTlU+IsiOKwHiR/ZaXUwFeopns6ZTU1c+xyzvunEyiNmtKrKm6URb9vLQaee2hLlDj
/0Rfdogznjt4Le7ya4kfDouQoXuh3lir+x4QPHxCUBxZTxV0HLR0h1gHKFz3v7CnlqaJyIpqJypX
IKKZ3PlPgz/YxONjlza7TeWwBzC2RrDVS5CkK8n/hUVuEHaZeYbDYL7KQblT4sMXTtPJhWJz8ypD
oem9Kcyue8zJRxvyGh0YG5i/dyFDM4ixKgIMudtrGlxaH7npPPH0uD7IZ7fenKawH3v1wa40q+6E
YX0i6asb5GQuSFczYMd6GUJV94yo44xcBJPXm1HQivv+YScKljiKCJJwwak1Khtz+cSEETDKTtCI
VqpGiLXHcWtviILlyQzMxHdbvcj+kd5vMWVfHkRQ0sac0k26ysZ7HW969IvkcQKaltF4B2w6Q9ON
mbl0Ivwf/h6kzJ7BsADTQDu3Nkw3D1oJrAHqAxgPAiQRwEmGcVipkHrxstKL/w5eGsYfmd/Q4eHd
rXYE2Nqgfzr8De10OVEYl3VUlaPfOVfYxIlDfagjWt3x2J3EMOpS5y9eKJIOQsVFyQTKpTvU4DW2
FvR/CetPvK/Xl5Ijdqeer/9P8NV12xt9oe0I5UxKm5AKKudysKthIEB1EuueBCCLkL50yYO2cqtk
+By2tVWNABSI7AJVFxWbVW/XrSfiPmLDXgcu6wFwfbf4SKq/gzwcfz/wgnxCpXP08djJaJ/jez1C
sZVsBkUdldiTjD6vPp5ES3qqLWO8AyrciC+hoxexXR9VVI2FVppJY2ZF/I99wNLm7mmqDw+Xk/bX
kBcEunSU10TdViQ+YK5d6XC0Zc180WpnS2CTDDgh7lbo3AhEWVa5smIN808/RmrTo+PgH7qwRghm
R3CH67RCjI/DYY8LatVV+/IpszndlRKSV/1tJrAUN80QHgCVkLDoM68YlEjE8FSHRaH7+b80fhms
XPmQyI5+ZMy3/iAKtTdC4ki4iGY27Argux4q4lLHo/Oy28AJDXjDGLoCcSKqoryf60pLpox8/zID
WhPJWsS3NQ5eUtymCzacfc3+ihG4D9NkTvPxMNo1nu0VXbkwtxbTOVXpybk6yNbRgPD1M04RKZ5V
bO0y4A0VNeOxaSCdVra0A0gPiLasGmcp5P316r/ZGzCe3WubveXeDa/F6N0srAk2gEIyjobscw+x
ymwsnOJwEF6mBHZ7NSJ2AFxp4fKmutjna7LFSM4iTWj/ranqYVTeHI4exZvAVXYktBJBMxwqNa6g
wuKgEZuRFb8laJPVo6/mvXFY+3L3/rn6QG1uDy8B/AWWe8rn8eMkBl+H8L4Ak9H5ZhBZp9KgfX8p
fK03LuFdi9gZxh+hjBQeC3qAeePTeoSaUqAH2qUy8nq8HjiU3RYZkDhzR7tIDR/mueNutroekkFS
tW0uHAxIe6G1NDb81N31DZYwgLQu8o5rjLKba99tBFh4IDFNHH/qZynWU46c7s+0AkAaNPTbrN6D
Xz+7wMcDMvXeWcob8vF6S5i8t98cMulLWccfoBYY7fGMtN345A8mrWOGDaYiFVnknpQBhIJqias2
laCBvKmSKenWUHbPQ3riqMAXdALvFadsEZdl5gJpDzkI4IRIeAPsUqmTZYc3IjzwG2crqvguXTA9
Cn/QcoM1Yhx54vCJ8Y+LVDjKQeKNHuCIXx9L58POZpE5JlDX1Q2Yu31gGeG6jnTw4V8mlgCOttgA
n9Dm9D8gpybRKw1Ir4gpqIXJzSeAW3oYDHaC0N24vwT3xAbprsOf80f8FZ0ioG3pcdu3M2q3brHA
PL5K12K1Z7T2qP2eBvWxgzmoi9d9FLWzetE0YqCQpqmL6d6iGk6TY8dYMwgysv93QnFAoKtLVnbS
j/ka+h2Ccm13G5dJFstl6SIelucF+elGyPWncLKvwrzQHn3BCdOVWuRI0g/kUzZNjP+9IDErnxKo
+2kDiYGuxmovzLl/CFNw9lJMneKUEUxeQgxMLcDEdajrF/A7WXoCcBTo//kz6s0G/DpbO29S37Et
PVxgaecBEEurbmyQw1TApakXtGCM+n6NVzJUElllzc57i+yijIjq+thw3bc/QagzxI7ivuvXqZX7
h25Tmyfmj/ROpC1TGD4z/1gcmT/fP9+BcQaOtVEVfjwpZAkdxnlCFTQKKfFULF1KmdhqMjiwl243
85hbR6Jk2nIIXWhi+61EJz9cCG1a7yloobyLoLmY72AtqrVqum1KDle6t5QaMH+1eqYd0vH50unL
SeO2nXLEA4jf/PNalbTmZbKCVY0084WrFPHiefbcm7oH4RaoEpk5vRIY+bedyal8NzUGZAyj/HUl
MEPUY7A+uGG8INoyAq23WwwsMpog+SGCDgKRou5jVcuvEw8wu6Il2q/EgKpECG1N+D9wV0oFZupK
O+gLAhA8p96pjNLaJbsk5hYPIUQ/fI7+BbjLIcFsFbGKoxeSUENvOUVqLteoxEhrc4ckeIw6Kjsz
x+fIlN3TH9U/GunxkSn5tsHuJI5+pyogMDpEaaDQikcaXX0LycwarnKoqqDePoc+a3A3I8YKeMjY
iBMMxFUNxcXP4qNQQeasa2tMvpKGN2+yWmOpWWUVrX89zz1KUMzaruIvpt0+0Aco1bsLqg0cvSPG
RCFn5GmKybG2e18RWrq4LVsLMCWktdcbV7N1PrdqYKJquU57vrpUSIP2+Umcj4uHZTjuuukN75MR
jB6d28/4tpBxXAgHZ1MsnrX1Bt2MJioFmHI50e0Radtf5aPg2KGzp0kxs3rnH0+aD3QMvpxabgkP
jAMZQM/+IOuLUTp5c2du71cS8EeoA/3ktD1cw3YD9iCWUIE0R7hsCpM+eaDpH9DXIzpKE6CVkXft
A4QNmAwEosg05bi3e6fQFN+KpT/Q/VOcu8SLWTRJ4iv1O8r3zcNQ/3HRe/WgveAjOplmRJE+r5Ai
BJ6cUeMzokY8fhu8lh2+pQx5QQqcCXbo7khOpkXQMrcakRlmOoCCfIPlm0v6uJRWogRAVRKHClrA
W0pQHo6NoyV9hO8DfqhLIMRiWQ8R2kXPyVwBiY4TvCaYLcshqWWhxgIf2+h4iLe9Tx5UTOxtrJNC
c7+KAEBqe6qIGCRZjjnPWSgrz0+0sMjpp/ljINhPHDaYdNPnnNo5VxiKgp94fL3n6+DJ39K8AiG3
hijcjNdRlPTHcyn2RcdnH8l72fVkUkyhZgzNf6GCTdJboKfxBGb6BjNInvvig5SC0iqvSA550+jP
gQh2feUrs8gSv5IePpJFf6IrGy1aFp2bDWu5kwmOCE5LZ4CeHFzTL0TMP1uCpy1XDL4/mBAVmeAE
542vyFp12pGPm06DSzdoHNJ+5NIGXYDDlHZ93rqCM1XTC+MuQhDWWhcKKBbgUw1zI44XkCXwGq/X
C3d/cOKa52tt6dp1rKcgB2J1eMMTlotXxEtlQjsjpS3ubhupA56bsOA2dDEH4tVjxLObedfvDq8S
tTYJmBEIfwOpQj96r/83JB/0oUVQODrs1rTvVaYpN7AVBTLXmev0QCSad9hbX8EdikpHE1s+TWma
63awONH1lZ7MZmzLreeMYmHagJpgvWVhIQVGyQgpVN9fnwKLuFbAAdaXnssm6fixvOsK1kjrx6zx
GK1DG0K+eRmtyvALENi5x61gPe1xi95qAfnK6fZyzEnqaIHM3mQvamsfJ1IPwrRzIeW0o283k4tk
6sTPFeJtLEoS4+Y2A9eREdaHDzyIFjqWLr1NZ/5XRAtn0i09LEWF4oXZsUarzadlJFHS+HtynH36
Ce1O5qWERzGU0eg8J5niMBOhBFfcWazl6SMiviLJL+8KZp0qvhHx2Kjg8eMwHcot34Rh4g+oqm7k
VvSgklstVMgJri4VC8vMjLogGIdyuTkpNAlRqgjr/axOGwGK2gxKj5mxMS+5ljOWcF5d8Tu7YEWL
hRmDyW/+X8SmrtMte0xpB0NlloGhC9VOXqJSZ5C38SMoyj9t4W0oDFUKncl3vOyeF7IqAjOj2Tkc
5pUucoU2hur6ldnVmAK9XAV4H5pGSMEsfn5fv1uaDeFb+ST/K7zt3KnUi1h+WFgXUEPYqWNTyaeg
gYEO2eiL9NESKu96bG2STihR8idTOsHh31/xR/2POS4k+GbckQAN95e2wZ1/WRtXpTHGsxgI0iBf
IziMkTlJMJsvGd3G1Dp2DmvWuKuW04nLUoDVaN4TSG4w+dlnjrgATqFl4GPugeBTw8cMhL+utXUG
pxLOB4PQaB8BM6vufhNqmuAyrUNHZAgMrWO4YQ1TvxidkvBz1dWxb56ZcbHPyRl/ZATH8fbyTKAz
cZ6pABXvXC7Y8LedLpNV9haKZLYnqR/6TIfskqWgts0YMDxkcn02bFKPZNDFwTTWP1CvR/eOru7c
Z3Gu17GEjN9MK09wH6RPOmDl8cWJuyVSQBs5t54XjUcmSQ2UX3JbAf1XCt2JV8LwR3diJB7O4xOP
AoAn5ICy/QRPAlDKQTUlTbG0MGQqI8RysN7Pp9aAoqokYT5RAQ/2Qy6tlWmwjbhlE/SkBaJ8bgzR
AK+LRlIaF4w+bsVky5vSfdjWV/duoF5duCpXZYWupTMqBYwkmEM77bAd2nlufU7b8cavxtjclaA6
DKSDpPgFYLjC+K6Gnmiuok0Hbi+AHc3Op9oJ8XwBF8LUYwq/l6XjCd4/sGVnGAufPhwLa7klC5pU
UWBkozVEU4ev8JgL2O/HXx/53G4tGOmYS6XD6+oCo4liWDCE9fWgot0B6FjBHunF1YEkHY1PR9TV
v6K3/C6xhn3n7IkaHoGmSoAtTXoMrRx5zX2blvjGk6J5HCvvYsY40H8Ruen8SMS8TRvcCoY6PtKa
AS8s7Rr+KpVajyfWK5lC9kuM4kgI90omWe+VDijjCfyWhHO9AGDzxVKj3Vz+jHm853R3pr6+u5e7
olhhikax021HQYORGoxIn2RlP4Ke2COJTlXPtyZ/G33GHgmWH8SpqiMszBpuuPElk9e66kN2kJhJ
X+K1vgIm4ZUhCRlA55iV5rk/plUxku0niQbJL+IHhvSYnQuMuhlQ/C4/ZYqftQuA4Qyt88B70gV+
/N/nIH9B7dqc57vEpNbSSmnNxStbcKOFzk2Dg1jRkQm6XF6cOMZm3OgBUbKgkEb05DOHHpgqsgAS
SKIO+0k4XgqmqbXez5BxbQoEHiFqRQucunYziL9xUReT5LFU5bap3xkNcU2Ge3yZ8oOaLi5pU2J6
qQ77609OqRkXmRqDPFoTJj2Wc8Pt5psZMxLga389BE1JXUrHe0bBOcyc+07rCghXHEIWYvEO4Di+
rfNjD0y9AqcOWwszFcgIDqJ2ZKnFLFMxJ5Gn1q/wZa+6q/ZpclSiMCEF13b7aNB5O6fWGvzf9KG0
N1GEB7ggcU6wcsEQRMwEtedmLw5LvVaRdD8u1iZZ2gFWEZuDU2Nwhb8bFlifjBHiovkY4o26e7wq
zxMzcyGzZdu0t+G0XEYfUywSSC1+rt7hHdFosTo6aOPpWkOaEHO5ue+NRej0ZxLKhhNAg+vDiY2z
cxm9/4MGxMPvz1wIENMszCQmkh9s+1cH5E0AWha8gbp+WZCJtCrfvu7mptm10xFn3lMhvdA7I2U+
8aj8D1aPfvkCdTqbK0rfS7r8RiX860FhoW8bTlYfiaaKFkn6BirUbAYVq95OdTGKK/Z7/N43SM/+
ZQ/0Krnn8FcdqHmYTSdBo0zrmmwCRfanWKZxB3bT+4DdxXRHlzk4/zWxjmxxmcKyFBgY7mr0T1mB
E4wc6EWDvwcc7JNScL5CnLr6WYYsSQSDtP1XtHVQd8HcQ5hQL3n5Pd3MwMls3hfHpu3S4XtVWcTM
jdceMAkMx2ty13GiulnGyCotq5OKooEXBE/pt8JV+m0q6GXmqQbqJwtEIrWamgs9IoI/QO+PFJKC
BkOz4I3/XOb0GtZhHSQIbIZtbOVuavdFk/Twrjz0U/kqEKemd4v4eBMZwwdvzjjdoKscLS3uZCpS
PYuyHghksUWNgkj2fDZqAPgXTq+FdShzwPa1JfJT6mvxjRJKT1M/unPuVkGjPbARx+E6YyjPUMdP
8EKGFbkCaa7QI9IZ9hRlgoyHN8Fr4/c2aFoF+7niauMWQntA7bG1uLzXL9AdttT/TCPB0HwOK1An
bfVjONmeFaWZ2sLhuL85Clfm187cYNVniAIB0Biq8yqr65x29Gr5viVaQSGPs/tTdUChlojTCKoA
DUrv6LaNURSelIuFaR3F07HQSSoj350v8KyicnPkDJF/0498Cdt8cvAjaDs4fKabPYvAg8dXRiMw
5ZEyANG8kvOToUTTRHClulSiSKb9F7iELG1Izgd0PgGraS3ez5nRrcIXF8a9eWd0FVgmzT4G0Qip
dVhDekx6Y4r8wJIcbNvGSOxuIRbQUDnwFyTL95F9mG6BsdVxOhl6OlooOeda4xMawi9ikgb5SMi0
HCf2Pln4cpGtnhyMg6og15YHGcf1Ug6Jt9FsBRtSPxlM9A1g9XRnH3mfmYC4h2XvM31cNBYfYMo9
XZo1UrW20YnaDE8ykdwW+0H67Xh9KzoREZWz1zWqEPPdezq1dGaasfj7ArXNoA1poEGUQp1qGGav
BRenpdsXrrQKqDSXvHQnb4AwIHvUM5aJQspT9it5UstptrHCZ9g5jRXyjF0eM5OgeAFjxL7H10Hj
AHV+wCR5JEh+Y++lsF7cfS8Mt/rUZIU34/DcCJE3zMRUhvND7uYVO8qcCohl4xtR5A4bx2PpHZoy
NUpvkFjZ4uma/ceMKADrYxYP+IwdsvC7VKXzKL7iPDlaAhtTVTL2falzRpbN1iJZzgMy3WLGGJeK
cBDYL/a0Gkgy5pvRpBUptR//BOQ/xRqOw7OkSA4lolcfBvfghxCrFCiP5FwA4pKOGYHHE8EpTJFY
xrPdnsAjYo/gwG8/YB51eEBEQ9Y7M8MqTAstaBtaBVQd7XXVDs3zuGQHhFPNdfLTFJ2ZUUUHixYJ
6PV6IPQAgAKrDfshf8/dJNndyUVpoMfozDz8BBSZai6z0E5/I0pJaPUViWl7Ami6v6KYJaamJPfP
OsqwGrjIBJ32/1078hOvFDXBpvdfnNugKzhMVGmeDYPa24ZkfI9SeCXofm9eNz7/wV1c799Burav
OoJGaRlG2Qe1E2YLcfdbqqJn3fxaeaBHppCxYfVXF9r5QhJ5vqR56MxWyaPU3zBhfOlnuAVbgcu2
Eq+ideIHfTtqQrOJsjnnFcluHYol46jthdA2gmQ0f7xfOZkaJSlUG5XzoAMt5MVqdkCR1yBbBjVJ
3MHUkyCJTAyHHkjSDRLoS+jSQ6PHDdeeimCwvIbPA046AjGDwupU6/pfDfZXegfcTNhB8KTkzXo9
WdxyCvdDjZbzUE8b3VqhQUo97sfe044BVmhknC15vBa1KSiqHyyZ0oIpoMs5GvPLOIlPEOc2sqdf
jwT6KQVHMdk25lrRAMEy/G5KWkLKzQe4Ppjid1GHn46lolR6BA3VEGpuBxVqIqpLP9roHGaC26Hh
/njFMnAW4gpdDZ6+1BlVYfaEamRIUyFNuGcxCAFtOkJfeod1kU4VWHVu7PjpAsBlPHhv63myFSFe
wvRs0jf8rIv7tHsi7ItyCkiKXGIVXBQS7I/l3xc9PIL13H5Z9XB43Z1IR65XgZUG8qoXdCo6jVsV
6y95veSYiFBl7EcLlIdWYVaRhmaY1yZMB2gITq3umJBjffsBEWHCIf0Z9/CteukhldN35EUDmtQH
yh4AD2Mw39+QkjRtaI52cAy1lV6GiNlGBCZIZN9QojRaCM7ITpvq07mPpYjr+iSWGjGd4uA6Vd6x
Qh9i5txp6aRIRLIZHi8z/QFX9Hu4Lu4kMRO/tyH6zrenpcwt298vpDQ/hnX/Wb4Ld110Btiyry9u
0T+W4ZVebkIjBAzLYIu23SM3l6/DQf3H4QrTpbgbplRrR8bP/IVy2ke+J3Cg8qd2b+HEULkKPKuH
XtlZubOadRg+/kbXKEGhIqrQrYJu/RyaTVqZdwqJ+ANrGme1r4La12fsSOHmpFH//KFkzuSAL6dv
+0lN3bK6rC+BbzFdpd28JqF0zhcmYiawMFJ8IPKxFcohlQ4wS541lIUCKOdYNZ57feogm0yklYBf
MBiNni4eN9Fr5d5b9t0kJiXnhOegvxAH4TmUl9a0RTEAvnjDsNPa8XMnXgqBmJrcOTi/agj+EaPK
ThHNvDrCuGH7q/b0Li45o5LwwHz7Geze+ZMJglnytCP91CfShcsa0kuEbSaE+ZY9j9sa3EZCdxna
M4YyCQUtVVXg/+xUJdcT6dgX/Nm26Kwxf9801B/WLV584pTi/Xr0NgD59kNZ082WFJg+KW5PxLz2
HR1HpDMiQ00K2T29BkgqRTH6m1BMFfB4l9umYu+gEYbtj8NP4LxIjE/vzhjP+kDSNCfr03iIosX3
H5FJCMmwdVsbT/pUMB7QVB0zvnZMnkHoe4o8vdpvznX/p2I9Q3XZlJJgUgrwaIGSow1YAOlpdVCu
g96BI3vU+iQ7S+i0uDv2baP+Ou/PbaP6BL7W+4FiIBUn16yY2ILZ+Q9o8JLHjah12MDlK+iWJvRE
SSdpOUhe+Awma7GADdvZLNLStKgsihbrV8DBZLtkt3V71l358HVaFAIYQ06Tje5AhnH6GdazuuSS
8zu3Ug4Bu7X4QnpW5QAOg0y+yu89G2JfPZNqwurB0cUvGLZRLP0uYKDDJJCJKOHHTBqQRgPXr4nb
vvOm95ml2zXoqiVA/2kG5hRssQa/o4IIf4K+f4ydaO6omPfxXCgw9xcj3ywbgfJ1y6BUfWSCLIWC
XXWOre13cM3WDdYKLOQ/F+BK4ZlKJhmLUWWFaV4S/HeZ0bwbejLmK2ogh7ij4U9PHYwbPwbJ7pMf
LmGZtZp4R0EJoaH4oIlK+vlBZcrfqS0+P8+Rt/yBjHysegrcfReqUumYvaingEp3HAspQzpYFUKC
zs8Ooj7i0QU+msDSLFv7+cs0mARaIkFQR4dZlXTLNjg4HuesA/E7I171fC/iKZ8sEaJIQyH8Xh2o
RnEe2ySCLbgwWjLAlmQICKDnzsdXK4bNzXwayIKVHq1B9ue87ev8jh1z1fNp3izqaLqkZbf/1zvM
Kvtvr4dvXgwX+kT8svL+947xWm9GbKb5BM61HY5oQLYu5oHP3U7EBXGeDL+GIIIOvg8ASaHIX0LN
fksI2MSpLfwpjgkTtgRf2QnEGMGcNH0sHs0QgxlM98BiqqaZ0pjNH0xY2KWSwJNLIc64osx3xPcF
xUMlDTcg+yMACg8DmrrIHVMDgOZnE0eNmJ2pXkx4b3qCf02ZYg3GZR9SaYUJAA6xAvaX1G4dC9NP
1ZJLTBtK+rQeBnHa918Kt6VnMAm0RSBybUb79HrsjqM7Zn1QG/5OvFzguOBhM39Ix8440enGiq0r
i0jqIZ9dH2Gp8QNAWo6OPIR1yx0/W5bRCYfuqzF5KY5UD11uUacVwTtIaSacayVWBZmW2HBTpUVy
PHuG6Dupslklg2KBcbd8BXLjuO4X+mkCZjtom8D9GgaPKZtuzI0M+R1eH9cCqez2odDessySE0zf
z8L4xgbUbmxRdMKMTqAKiPrymMGC7W3CayNyPa9dr/2HFFSzxfsxC3AhJUtiiShAUcs/9gVi4G71
d325VMFEjRYznY0yToyFXF/iknP2xhzaqPDcyfnErhYEkSR5UUzHw7MfxOCExHvU8Wpj4KiMLH0N
f4w0d4qtw9Mo6ftHgs7UCQT5UjDov7Rgo9h+MC/FqUmSwMjrFrIzRcg9RweefXyC/VLpKTJiInMD
e1+cTOmH0DK+vSbfwmYlXJj7mzH/RTTCduCPqqgTPpsUZMK/+oILmvc6RrcEElUmBqd2o8zwN7uU
L3b4bDmjQ68EFgNeKU9OkX83REsW3nNMsKxiWY7gPsTx75ONACT0Ct34KRVNcGACRoLniWXDOF5b
6q9BXmdM+0EThqmeC11UmwsSV1L4ZdgHCxVwEbbLbhRNry5JaS6soxIT1cjv5JbiBAXdkXKXsvu/
uTEH44r4PSuNX/GEdB/2FKAgrmOCdM3Sw9p2nu9cCIcS5d+mUgWM3cGSoMVbmjA1Dl9tWeG6AMMQ
33UZcM30PleBITVqWrp/X+NVVzfF2BYg2gzQZLdqBIpsm4YEF2hVTG9pOegBjqiaNazQTrux/b9+
sWo1A5zZ/Cu7wgGiOEg1uSrZsal69CWTINIxzDJ7yBXNJOoyZeX2vnyUY9im5w9c3kMnAyexlItE
/a6x6QEj9622rKc1xZdk+wQUVIBXn3YfrBso3NsovYT0rbQn24j+RXkJqwL7Q8MG1Tbdgpsf0rQ1
MBCkGosu74lVYelPyQkohTlFRfokxOQZsjdLgmyvcSAJkQUFa3DbYMQGB8cNLoGoNfQ+8csPLChw
9/Fr3bxDkHIGtXozNlT5o6T0g6T7NtPulavqorOL7vkKM8dPnB3emAS8vJG1hBSL9WORq5NXg6x4
eK6JlSDk9T8JKML8ZvHR5gdZKrBiF7c00sMY3twxHCT4N8Z89aytbQ0L68ogZr7M3dmDlwgyrfri
z3QYyE+4jtd1bidvGmmhKu3VgArWKHnikikK0SY6S9LSkDyF7WbE+MCpArHrfpzVhTNzGz7QtHk6
ftAMyA9y0K0GmmMDD2RBigWqG4saAtyy1katOMxhdklf8NlPFndiA8GSIiofWLDJ06FIAfQd4t33
xm2U4TQYolGCv29BIP0z1kUz2sw2l31b5jzUXiF53JAWNnYHFcshcDdkgV8999vesD48NY6FfTpT
w4R2DU2lu1k2JSdT6XJrPGjrJ1g/cBDmGu3q5dC6Z276fLdp1OIZMwe42lkHDGd7yPn1ZGPusRo+
DiRPbZaMVjdU+MupKxro5MPK3UybGAm5cOW0gsOAje7UFtqd7a/I0riSHbLEhdxb8ImfRA4OWh8c
oblG0RqvPYIQx0mcmg07pNCest2jEy/lZ7tCeWmISRQkjqP23N0dKjZ5d7+3knaxPgSg3G6jYtgK
WKolbnEHLftavTCxVZ/01lPczMr5bUIxOMtGJnbQl8Q/505aVZ4cq18/o0Pv4CqC3jsu0yb4pAu8
cUId70In0+ImrN7nGyI5aI6NXIldr3Qx518n+Z4qeRw9/Zw++fimZDZUKB05d4EEqOXvQCDh0Jcp
MjWqB44rBuwRBQBCEuIi02xfioXTQ89vWc/lHqpkZUfTeOTqpfVBwzNX3t1dVbBK0kqDgSLO6DqA
madiVejrcE+6jeqoFn63r4jWg3eQVxB+OpJo4fjB0YW1wOzB96IRV8afxocLo4Kamcrzq/REIHxl
8+DYqsV7YIWXo6v02h0bEUAhjjQlAOnPfsWGKWa91pebgJb5pvx+UJla+ruWWveQKbsaAbY3lyVj
IBuSDrL2PmUOySGqT66KI55+KTywWqMq9DDsNdkWHXwiMISkDnYUbtyGyaNRH881rt+cb0/JRPyA
0bjIcBJN34d8NRtPi1H1b7XqWX/qoj/L6AFoBR9OHRyQFpYn7lUoC6+Mq9c7RFBaWknHKcUClytX
my8jTYFIv8yqkD3j5jciA3wCXc7uFubSVJ48uPFJs5Za5ytg8Mx3ZbqxowbfbATiU9j/MEtfVd6W
eY3k5GP0NnqJtG6ZullxvTAtAmARAtVa45h69ZDJryGiCRodx0u36NO32chfjeoCZDWa55mZF/06
8yzotIelZwtSjOH0shVwhaCxoBOpL9b4BW6zERquNjhXxyyW3ZbxoecPVMHrjhBeiOtN9ir5Dgaw
gQ/m50STMLzY7KxUX6TJxox5Ysv0SUAX9FqTeREGsFPSu8F+e8VtFzySpfZZwx7tpeZHvs+Y49z+
0iwxaEbwnkDNHzmuKqf4PBnrXu8pBa2Ftrp9iztLijfdNRoknM9MV92kPQgtAveOeTGP3WdljJgT
191FNz1KBAHdxrwD3CSRGUs+2XvLsQhUxym5FIDI3bWo9tFLRGj5S8G5+sIOUQtdNsx0xWlzbTg+
XrL7ITMKTP+ai44QJxZNGxwVJVEPIY3EfECnJlz82Lfk7zqW6EjgKG8WhP6p1nWw4JZS/OcOBPoi
madGaWVnuGLYqvAtwV8FUrUysGxRCWpEDBFxfW0v1wr343uIRWnbP+a0iEp/7sDmKZtCFCYgGmfk
AZ6x/27dDdmPfolPi7A4X5G4GMAeH5MN2PHwpfrywO0o59rLEQ8J2aFSIoV1SLlu3TCVT+nu2gnl
WGXWCa51kSQ4iXP2fhtAFoX8PbaJcDHTw2LdN44YgSPaag5pIBvt9ompV9IBVhrkm58AaJQ9uDT0
K4eFfLR2V8ZN+A4NpsPKWiX8yPnfPURtwQmT1rdjhCHROCKvKHPWu89+VS0azEhFHWiHix2ILrwC
bnoDRjwWlReVOkx28QmaUZqmmz0e258BJpq7TBGB3XH06uFNdQT5wLRgRS7mS6jm2Q+cfMV7l1O3
Oscts+nCWbU24q7LFToNbVwA1gHAlwDwo7Hf/5xbKj9d1JLKIEfWFxN7PddNdMS1QoON13BbQSoh
u1prb2guuBWn8BKB3pOWp+qjCvqFwHiuh93mu0PhwRKyV5p3R8O2nA5lfejZk9PVbuVt1+fA4d7s
d02K1wZRODT3m5cMyPW57JO+z78H57d8vBULXS+sjgWurxPgYhCcJLxdzIA1/3qPkPrz7vYB6Ftv
1pnmApX0k8WOMcunabV5M24ekTR2qcuS333rjsotkq9GULEr1h1M+KNlsryHw69lPppvv3FJV5FI
wiVIQVTs9ieebMmb65QavKem34hYdT7zs6NGiE70zcz7YLvb2xq0kvMzSYmONWL00TxZ9nDxgovB
8nPplONpjPkynrXsR1Euas+qeEb+8PLh1OHX/nEC9ecicxKmIeTBVSvN+lIgX6kjXdkWi2uj3zm2
lc6gkhNNQwJf3w9yWEAkZIrbazY2Z6ktC+M9v7oZR29PQoF+YesEQDUKL2KV6KzpjdTgZPKs8wZZ
ArGniplj1xhp383h0KH0A4vyC+dogct7RXaYUUKB/2CveMMN2ET+/+nbUwApne+nHaJ3Frg79Xl3
8ANlqpyWmhGYV6tdAwCJaBdkGqGuNiUN8WUu4Eklk72bpKTs7RL3x68c6Vum/DpdMdzcV8hkLAF2
7ydH2vRYLcgUwKyZyOmgvQQJUkTUXCjTnLJvIfQVgu7jPuKN1vQNsHhYkncDcVSj0z2rWetgG+K+
NDGYUll3kE8AL/GdRFzRsJ3+EeuesoQ/pIfp9GmLFMWJGDlHgJs8P7PQmU5V59qYWUT4DYUNbZaV
YcCZQxZ+2TzNVioJs/5e9FZUq65s2/UjwQkFd3CyFFws7B0eb+CMF/b9huDvZjQ8t0LKSw1Ffiga
pzbW15vSr+meFXYoMZP7HokSl118gTQPyUGN+qKaoENzJdPhfnRlL0bW334tfHpeUfDpYJciszTJ
TgSNewWg27+e+iq3Slze8O28XpDhPHzHV1m6cVV8ORM9aOA9QDncRygFwyniPazlrn+Qkj/sZjHv
iYdsxyOK7vvC/PNn4H/3AJFT6zIq5FVmcXwYxcjHtPv4H6UDt1Id5XIVaC21jIbkWQVIcv0lAJUC
DZOy4GcYF5wBGMDr59c7EyrIpLk0vv1JGkGW4ndrpvyVGkZlNd5Ngz26BprgqVU3XdfN1T1/KVEq
runL66cFyOZNj+MlcTQR5o2Ks7YJIR336te6gArbIZ3J26RSy9cswrUJ94oemobfwF2v395zd7CF
+1Nk8sOLjQJ4c3LzFSyqPviBhJTeLZr06hx4Zr8O9UjOiaPJM2LYbu4l7/kdWk8gDlB2NygapGqr
sn3OiwDiO1npHN1mTft7Cq+RWwodYN6XOqf664t5r6nRTktuuCnv41hFAF9u+p5gezq0wvAXH1Ax
juynUtajH2aQ6PPMn2/cro1GBiiGpWdIUKl6OrghOL7lkK7IdfNemdaujQKwa3UOJ0118Jp7RXuH
GxNoKLFF2E4YY6yDBz59rjYZ4kP9hSuRIjlhOG1g7j0Pqj0aTdYcQbbGOju1db2aj7SZAavt8P+l
NaGxd/iPaEsUCLJDJcVu7QchDJ0b1mdpkbrSrfR6HOZwQ2ItDTQTXDxrMBJE1qJKAJbImHGMwVER
3Y0ESUL5G77xcpjwGmOhMzDcQnseEXngBs8F5u9nKXhKnoCfxawnp4znyoAF7cTC9FVuwLmR/y1t
bn/9QjJwjBs7oqhATSwUnyu0VeRFWbd+L4UKBPg9N01/o08SP5JYipth6iFzh0SOxedG7nlHfK6v
zmD6FiYR2xVF0nZBLM4ra3LBg9o1SiaC9HyWkxmWSTe53TtrEzG8bL9L0FSMibvq2vYZMeIc3d9t
JqOW5JI9Lw5pACdDcdNCoFwTjMlbUJ+ZOeCrt6sWvkAI7kj2/W/KWOr5rwbgO1li5AbFD9/e9lwT
xj2rfzWPwKtwXYDWdzVyjF1PLVmKfnHhM6AT78TgEXlWkTfuAsahkCDhnQr9H98Q6P2CbyihUKqP
N4GFD8OfDP4N3TWGM3hPhfZOvB55HLlr/gVmRbacZz8bL8dtxYwuk4N9yf9s9P2HQc7H7IHIja36
J5J3bLSk7eIbwaRNa6Kk9L+WwtVXiR/hGCsghNiTCJ2csbXURsyLYk471Za/Fv2J6MvPerIiI082
ATjeCXA9VHRyKS49ZI7SxFY5PTFbpXnydCk1fysusHIU8CJ6uBOizDxGe33dyfRPT9hzEyUXdzyB
CbSLwLtjQgV+QBI0ylHKctIGDE8qNLjcpYPQrqbdyXRITP2kSSBbvlrLssnIlS68ELyfVvKk2Z9G
AGhbcDhAkc3QYFzaDP+IOI3kPRfpz0+RQznxu6hrOsKPzY8EtKNs/rCaACfGGQd3fDry1B67T5ia
4Clnxd+yk2ZrpYeE93FelcaFBLZhzbJnqkIqTtdcl5yjq4WjnoQUunSosL6nsS+vqKBxYx1c8N+0
nbxvkhhH7fpJfCuMsxk9CNHfZfVyKhfxsEIVu1jeQDDeK9xt5fzjnvzJmqQRmCB4T3UY6FPdtAZp
MDXvx19STyhHsCErG6fve2BJuihUedAUnXcDJYTJn9pZZU8+MzZeQMKMRrAeKB3bvBlwajji8T1B
yhxTDQGqmhthDHSs7k5EeoFSKq9k+wQupswStPDfjeq2gy68cQiWky1ptvI4QDr7OBT+jkrkrZZe
Vm6amghfp1XyBLERb5b8asG3lFq/NoLhpzzE0EFP1xldJ2XyOLdc6XACUlxBTFpVFF10oa3frPfw
LZaWUqanNbVT3AubmMLb2Whu6IxMiJmRIwiNt5EPWP1tSX5w3YARX2zpIM4UInAXUYSwdI3kG6Fu
4Uc3cpbD2RPlQoXfaDHsbQrZPnk5fn/79PXu469bK6oDno197vtHt4Rea/1E1YxfhRl1+vKydiWR
lLWrraGxnsyGwlVz0iue7JnLeME+UVEG/8Na2t4w1406h679XrL1ld+gsdh4PujTPKHn/P53Blz6
5fT37hxj2WYpC7dFToIzhg2dWUPEOyBFlNF8iADrju1P8FIROyu7JGD4FsojtZ7N5Z9JslhJ/N+f
Cu4E4REpbUHyYMuhKXJVy3NxgKUYZdQEybwFZv+h5JtOQa9bZ+pdNeWdBza1xr0/cF0v9HgpLw++
lL7d+7GI8wroeo8h2Qrv/y0TQP7n6sVKMjfqOJC1icgBIVC9m2PmIc6yKIePnXhEVKnlfbf1FH5P
ciTrobGAdsm9CyZkEoCIlG/rfhhMDxlMgB6f06E+WSTvtt+kGbXWdsKo/lGbD/lIiJ8BOFC9O67Q
5GGRHlq2Y0UTVYfIAv/InAN/W0OMChTPrkmSfpHiQq+4kZwdmYGcnQKO80S0mRqGJP2ADGOvcc1N
cGMRNqDCe2Wo97hj/5G/loUm8Hocpm/iqN0jIAWKl6NP089eMbI5lWXm4aUkAjxv9PB3Hcy1D8+d
yvRDhvqMgCcigccs6hWUR25d72iA+Lbt8tGKRbnz9/wDvbtDrTqTCjr7q/s/YBh5j+5OMtmLpVjC
ajwwWfcBJOLoOl5vrRvmJRRDChfHtpX8p1XNOoFaBowKcvhCwlZ4FKJwnrx3qNUcDL7WyLihfe+j
o9NqUjJNwyv5STv/MC8o5cAiIeMjj/xil/1Z2jQqjMNTWBLCZd4WOw8JAQFY0zy6X4h0oTbD94Mt
72nc4fNEJKdR+70uW9r+ZOKIS/gDQ7oEqQKj9hFSptV2lKFWOwGg2EKajviwvWBCzx7xnZLny/pe
vJUEC/8VNyLhl7RZHn11AHR/07Zsy3V6jrzqBKXYyLSbJUZGnbJYbXXEfHvv9gYHaKHIz48MLL3I
bGshRTVpd2sVmfzlNVuHHrRQQi572BufljUXuYCxkLNEicW/jBwEotWOQiM0Z+Ond+OBI1T9mSAG
QEfK84g3R04x49S6n8tmliUQYM6Q6Xcp+x9YnY+3+Rjk9kQ7CAuyBlQNKHfqg5+aXrdWfzrkMXEx
uHej1+JjJ7mktxissJRprYJRS1GvvIYrC57chH4W35h2hr6VCGOmqtESdujoTTTaJ1IU1zBfnxk8
RuDOyBwo0Jf1eIFNztOwExXt9viBOhOGs8FfVvBqtAFX/y+2K6H2V+HCoZ218HUeGZjgZ+KGR84R
/Y2ax45bmoYUHL3SVZu1e/mU45+8iD6ga3LQsgReV3huWNdKaTo0/gb/WT9T4AoYCtaXIvkGcAW6
M2tZTqZHI54z8isDa6bKcx4Y9NN0uaWXLhkkmm536kvralX0dTKms3gJeuFqgT05I89mIz6E/gev
p4R6/UmDojICXpw9XNB/D3EdEPyVdGp7sGePKP+uyLBPHsVqvxDvwP7u/KGqnMj2XBzNNn0AOmAm
ein+2Gn65PPcp9tRHgrE0qATv9+dv1/kSPFLvfByeG0XwOOl2A7DBTs5H5Igb+hU8XKnsic69mCK
2Peqdem+kiFwmf1EGGn9DrKvCWQNNTdFZCOMM1IMbUU771GYVDxa/p4ca91D7wIEtMrTG58qSGIR
vLXHX7LN1dMPlCrZ0GVItgZrwH2KXqrVpyj/FlbbxoXBamls5XKMe1h7xxXipDVMcu+WnOI9yP84
2A0E9SKXUkh4idTjSAONKep28a6wxqzYZgRWavSVI7Itp7HT/Uks2Z6zEmU6bd8dVUfNmg92Pa0+
DLBlPVCVQHKnVONY40xmcpzJcrYxkKBA/trOh3Zi5TE+uKuuoXU++jBPI7ws30XMeC68qU/Md5J2
mQntNOjw0msyq/CX6kdIu+KJaxl+NEqR4M0s5EknZiBfcT6Yv5OPaopVcVuoAZcgp3Ah0GUoXRoF
eysj6YeskyNGheR4XbZVOfjmeQTSWlRzku2ChaehIL4ua5CF0mz+ej42FHYRKsu7czcd+6X1ku9m
7xtFUusM+zdAai6eZBw1CwREpg1u6xPxzQASkcI0gGeezXQQCm1UGHv2WVgB+JmftjD2mivP+C4q
24Jiof8oNFUW62tJW0DWFmdCnB/e4qylb2D9uLebHdus23AGGnyjbCJxv3b5vkuCG3S+QbzJnzaC
YI92lYGwEiNOqHFfXmEPtGI8Dy0NlXBp33XvSWxnAm4BU4ZFkfH90cDoHrRRuJMBm44eVJLsh7h4
O8RmOgPPHsae8KmVeVJjOtNuSkFxyIxyRyWzQclNM1pa7M4PZEvvQn3esnvOIEhOSIJPZf18CVrK
4bFJuRe1c2TH8vfiRobdUpCLkUAqFuktiDY0o9YLv/Eap+RqmpIyMYs2TypTrdDOsV3CLvra6jMA
VsO3zIViqOtdr1RsrLiE0s9r9B+gILhGxoYnAUgwmaxXia22FVXK6eJg7KXtYOHrb5m3fhNmMaGD
Bh+TiNJJEI+CW1sape/+rLOBG30VrUwUlVbWZTI/1JFKsBp8McsTIyBLob8e8cNKGvCiAxqhtm/t
5afH6/4E626yKnn6e5w55WJ/2qF2xo9LQAYaB174OIBYkTSJCuO6N1+M32kedVxFDze6p/ZcFqjx
w9YY2lqp62Q2DmmfI0ZWEjsefbOwG9vEOxyagML6aQeZy4Xi34qiktpSCXu4cMXDA/DbvEa9r3Hq
PUaITwW7DXu2pGs2nE2nZm/YnVMj3/zvFnWOKkM0yzj4nfPbBrpsrndl2hux0USvo89jxgClq9Eq
6M1tRZUpPA+6YhyMqNFmA5wrXWTVL0+ke8iBrBdaR9wgVeDl9l3yLShwXSpFtZ22CJGFSQSzWijv
8LKIVG09EdR4kH4s88yYYuyBKP7NxhP9T6GjcmKOEcG/YC10rl4h+WHRgr/KjxZF4ibAHAre6Ogv
LFjzcwG8quuK6EKkUUCwZi9DDYN36GsY+bPTRYyPDlF8G8V917/Vy7CQeybaoRdmD1u009tj7wzt
1m5JB1oOg76968NTC33cEfOofdBIoPCGQvhBT1rUkTkcMaCULpLpRoVbq870+N+LI4Q77ufu3Eqm
jL2bbtCqiXK621ru7sIqrpafQ6oC+LXaV8Y+PAUZEBHdWqrRVPlPFpfPfVyoPoGLbIBU6F2sHgM0
nT+4SLw0dJ6aKEi2/CZkKCHgDqscp+sbCWo+IMvQEGvnUZFxwjYQCoLBbw5dalZQZUbCV3R2KPYR
Q7X/LwPJg/QffaizjM6XWoZNwxNsDhEWuXuPTV4ItTqy74oZViOmV6JzXaqOyGbrTRA66om6dQZI
9cMk3A6rdzGm53Unspax/Qaug/OxeknqY413GP4rM8otgMJeliUSedoQdEEvKBYfGRJr0U+i/ov+
oBTqrVa8kaXu9Dy/clC+kftj10iAhqMfda00FmOftNuGJmWoX2nD14bf86p17Owc9zQpvHwCzFJf
pSHE0RU9sdUPkB8bwNvgjmYSGeZzIQnzZPv7pVglb3k5bR68LAhkSFtEkepgjot1CrfbMF5We65h
shH+cfIoJLcyJUVlCW7/N4VLNhigOJkYxAG/IR+12GUGM0oIRjN2+j2DvWmbuWpIAuF840YI4vH4
bn1z15QMjVcOv6YeygUd5saJvin2tBCE2X+wUAonYG+neAPwD7HE2BN49/ophs7s3RbgI/ndBybw
N4QRSuMhd2uM1t/bMmuLJzoff+/FCPDFxl9Uzdkcbx1AoXTRflX4U7GvgP3evys3irc2UQSC8kqG
HD0exqGcPuxTAsqYLITOM9lj9fULj3JDjPhsKM6l5u4zWSIKWtg4xvZ8f6QjLpoGdnMo0hMWJE3S
nBNZm3l9h/LZacKxRI7zdmDJLc5BL678jBh4fqd9BMA5/BXz4RW4oOv/c0TdzDERzIlV3SIfHZKO
MBgBHsYZVSyZ0my62S9eDir9P1/FqU7kx2f8ElkvPrTbCl/Gd+mppKfeQdOfj26oLkHlbsNRQfzy
ZrITfi4OoEvNeIN/21YRkfTRNGZJaonMLUlBrYu34feo6VDbRnV1RxWKNNFfRFEKzvRr+I5GbdvI
/1V27M4pvUeo37ur0maxWEX4MH2m0ntc57b7tziWvtb+o+KMy72wHrlzW8JD1R4ecdJaJ3v0D0+6
sNWzRVoI6dlp6DwzaLtukoWdfA5dSPxpcEg9K1zFoxpe/nnhphWVdxYEIsTD7lYPwk6p4abyLFwi
0kAXD1yhSwRgmX2r9P/uSJ1+i3yAUd4STMjOahxyF0ttYaZuCAYaP8jKZjVyXZvB32de3FmpAP1H
hIlrSK+zogIziDUUizfOnTY6foUjhLrFU6yvH09zivyqkEi1bcK9n8ZhzBFT9jqi5XhWX1BEh/uU
k1eJhTspPYdt9nvuc6JYobjGRQGeCpqPcVwZ5YIH/0EKEWqB2CDL145wz6Vx6JICaos+y53xeogM
u4PlQFcxUUiYD4vWilpxo4pSWhQhVVRsRU6iQecKlnEaWoCTmv0jDoPaoa2TSl+dlUZzrjDSI0uo
BItkDTrkNXQx8f2OEI1l7hXg7l50JfqjKinqM6+ftEvA1jHxFWDLDrvhfI6IatLBoxm5Z+yK1+IO
CwAU8b2CsUZoPSjXa9q55HjyJgwWzyxdq2Fgf8jXuQ6doyOhgqxXIZeoOOeCTtZbbGta6BnyqP20
2e7ipwIukJPAdA5GgPj8LLcN/dtaSflIElu2TJgn6mhbHs16CtPL0+24sBnaeA/u5LUYO4xvSjVw
IZKigtLvzu4O/gPwUaay58NopzvqNZ4IKWIJPVqTZFGktuVxk6zoGq4n6rrZY4j1J7KMLvBsJgYj
4sBAF7yd0+czCNqlCiJZf1zFhKJZKQ6iozQ8Q0oqeA8t4X9+Ma5Oj73dPqilj8VWNeH7KHky8pCQ
LJbvdJL5/lwmzm97Akg71fZ5ukLM8JlCKh2+t7daKcVhVm39xxTfMMx4CfZsjoozupqvd22A03mQ
XSLeLGVC5cj9MD1Czz09ZKJF3pTIjaJFmKHdIdyy3jn47xhkzilWEaGQqSi+DEmhw/tPxjondkME
8KM/KLaQOAYYeh/bPPOQShKgLx6lbzb3KUcDp+dtkpqj/ck46CbVc8XBNcM8nCh7+9e+HLdu1jWe
fuuxZSj/fhmJAXXEnT7uQBG14+/or1+Qs5oempyOFkVHc+IT3lD1VyXloiE0vx2FEO25lZG3sbE1
Nk0TWkPcQ9PZMUyOVkbb91y+BoU4zNtX+GnOMxDDRIjNCk0PgiqkzAxQXppZSG6x2TPDJn71zm5T
PvQxzB6pnzHM+r/LWaiAzx44a1WJMtB+RujTHJ5lO62mYX7es3wcK6jxUGDaD9D7twSgmhXrcQPy
dmfL5AVAYc/17I5B6KLph3gibx1ogk+KS+9MO7b61Q41yspLU2PO7/dMbTlRg0FcUE3LEvSxOLNP
Dqihuxhpz16T29VmpyuL0P2ASqmk0a0PskUI6ZbraBwRu0uDxEv8Y/UHqVQkom9eRvDyd8osn5yC
YbtwtCmSX/6v1esJICexOOehJlZVVj+lQGmU2XqblBANo1RS1nW8h0T8vzDzssCQMN8HiWx1QUAa
7lQ/qEcSSlgfJwNzSL/3+rM1LLuKwN/j+VSJD0IOAlgwJ5LuT02hSDcP+PrFAgOD8T35QzxBqTaZ
wawAmBIo+4up0WKchGnfub/yvec3RPwaMzqcU6cIrGnOJq8uoBhwSOzUb3rjwR2jrEI3mmI2xV6c
jRNgklIAFs5y/CIPhS8EDxVP1Lhl8Cf/gpqrltriT3J2txorwFSZnpOL/umWrf9XanibufX28lGm
wyK98lqs125FDTrdt8fgRWrSrvtaXN90AWoXYj0vXolkxDXS0rMdYn9sFfQH74sSTAe+JdMxyd5o
ZcmJr8abCtfjnRyvfTb146ShYKbH3mgRH72uXth5mA4pkNMNvEw1t2pHv2fd7wO0cbQNqZXvKpb7
xrmSFgCUPqQ6bt+nO4y2i9qPnWw3guT2NMTlm4ejl5No1t19AUCWyMNwWOQFkblaXHqaH7NYgJIo
fXI/sjKpO1h3t419XXAlpgupMkrGH7HXUJZmNPXaIi+ZVuKRwJgg4EW29cEBaHVVebpIWtwX/3q1
tqRu/6tzsbqYhWX/7JJ9C99I4f2hkaWLcd7iMGKLyS6qenIV4lvxqcnXMfp0quaqqjezVqsWw/kR
JdADXKkE80l+7Ykwn+Or7+MyBxCiMwIwQFgvuGT+LgKrKx7Zc28xKLPeGPFJhjLG6GGZxrTWjlmS
juGzPm22LkbW+tHViy7m7TcJMRDik5p2OQVBrAg41WPu5iMMNxNB1oQZzMfLvFd9V2Yz5tDrnJ0W
Do6FSIvaWcDxnsFmnTcOdwm7LoVZVTdEh/IC7J/soJQKEeFccqVWK5OKZ2+z+NReBTiKqp5RKqGz
gBbcFAHZvYdMcZkCPWMCB0BjEtgMjqPK/lQ1n5quCgcW4IxxXrwndH/Pgz6zAVxDfZoq5Ug/e8OS
aZqaoWLCJJ7kADF3i0E6dAXSMpfcT5fj8gF5zqCfHRlkxcJcz/0qAJ7eb9GTj/z1GXLlutBQSW5I
4YSBp1+aVF8t84n7B+IViHfGEJU5jzkIzIDEddWzhyWo1o9bhC7UX6Afr+ZTH1NLUgztSyd/bbrT
Z1Rwc0BQyoj6RBT7LHBjayM8sdSIw1bumWJ0JcJTsDrkYDZTdIAG5YzuvBnmGWPDW+UEFlTkNNYK
DCdZr9/hnJa3KSb5qIUjMZIcClanmYBnkfrhFW+C0TmolSmn+6RCaL9XwY4R8ceBGJyaYpa1nrJa
AjzlFQu6vMXYs7taQ17TNZxaqo7VK+vgneBE9cSi0mYEzozxc4Z5zAWK5lKM657xHntUFAh5DClx
E1YIsFM2OMNxJh7nra6vV0dNcM+0gK8z4xuOy3tE94JzsFRjSWdwCbUDLlEQeUUDGjcxF9fb5KHN
A/zUyFDwxKOK29tEX/ImBgV9TeA52NTUhPiydgqB44Outka9WWZeR262IP+WTQI4m+NnCa+CT1d3
0mLSsMhtix6ASXqtWFM2E0jYNrY7WS5PgdIth7zd9Z3hZ87LgqQQ3pWRpvBqSwnvYhISjHIq0Zqc
sKEd2fXHyUfR0tabjgy9VnFMSCCoP+f9GMEWlvFaNN3PseRqvwfeZMEJBAMBTc5hcn2yvDgKXjMY
3VnbPMZ89lXNkow6mgYB/uHiZQUt60zWiI7k6aQh+9orppfzGUcPG6nnrhzyWfa3dSHd/UW2z/9j
9UxY4H7ilrxXQ7668DFNXZLGLC2yEpuikn2hRuuxOGJ9jvQyj7JCRpPjQerX9KNDg4a0lS93ckNA
H7lXtj1mZMGIDnbxdPVg7psTZzy3VNnFrxJpONud8udBHfnSHRyshAyrGFYB46zS5rji1dIKQ15C
BkHftoNHRyw4u3yiunJPEaTA+sg60dzcn/ibHwniqEHJSEqztmjvcAX1fjdBdMhUZQpDunNVgmJh
vtWwFRfTQR82myDuSJtTtQX/RPYQatV8OeNjrdKPpy38tlzTTGuBAc4Bb93RFIE+2OR2lwEEXWSJ
uMLDZCdyK2vYYh0rPWxKZDtudrf3etpYfk7ZiObdlS6fPB3eVktXFqRMrnMaPguzzqiGsdcTHWV8
2JBNFEiEY8dH+Yw87Eo2X+fie1vZx4ubTTf+wj2Ramh/uoGTqlFh0o+4HTw5OBq0D7zVUNi4XcdJ
s7vWiXWlgpuzqEkP4JBVeJeLBtokKBi04cbfcDR6k4bqTqKZ2hIrw7O6NOHjxCViJapWx9keYAWk
oBae5hj1/j+ZFJkSvIpCnJFKCc4pdRtN/05oJg9gGIaUmL3rhPPQQWIPY0rGkeHq+jOn3ozslavl
DXVKQSx+XqOrXLgP2HMbtxRjNall8rKSDZz+7BXB8aT29rAT/BFzdxEuPOjToW6KTmNjl/LAg8H3
E+Nk5XaKQAY+lHJyvMVD5FkGUlpBdrl3iuNJS07o7sDu4Tp7IxGyT/CTnWQrVsNRikFs73d3XW53
GxxWDW3IH8VODhLAqm60RsU0eEUWELRGPMIoVfyB+TpyNwTr2ZeHoIndT9YgjEkmPDiDYOZEawdV
frHYd9aimYreynQVujKLD3t6PgWshwMPCVO9qpzykcMdypoEBuNu4WscZ1s/ZcCi9NhTxH470JSV
/x5Af2LlJwP5HCVNSwc0JQ8l5ojW13O1D79rbBfx7VtBTJE7YmHoL8awZ+ZTCmCWUYiSXaM9aqIb
dbqEfBC+uGS2tq5c7FCfwNDv29a3+aPZRRpYMRNr9GVNC10nCs0mcnvHDQezErM2MtGzWkimHmm9
AkZPscB9/sopmn2zFibRDQfwsRuLjgPyhiXBoyNqKSR/5Dt5019FnQSa5vbvo9xmqC2Z2EBmVHwr
WSYdv73p9hXjPQnmSclhbA4Vf2fmEW0jxqa9/Mhd3wMwwj0jwaKM1dZ4U6X6V5ZdRngA0V1stUn5
zHlSsG4TMvR5ZSIiMbO/SqH+vCGuECLB+W180hkETkGrDBGiqq2989zFf7QQVDYYEc7ihMbYpeMA
s8SQ0R8qtDJOq/osPXuYFW6ENTKmSEhI4xBNiw61GVNMEAZNLPMug7+YQ9WFQj/C9uJGlhOeHWzO
TbLDD+8kQO13nA2OrqkLOwuEuDf+D8lzAI5Oh/I9SsAA7uvgKEvNw/6dqRx6JnQWc/hDb1L7Xzeu
QyOStdv62JIpEzXX9b4KEE2O4uVZls63Gs27Y4SEM+KKXZbkI2x5hVmb7kcvivn6Md7+MMQoxT6v
0Cb8f0bemLucbhzW7fm5DS6mi6dakNRazW7LCpJCNJSO6uuapqweM+QbDT6UoGhLHdk1ZWDXslI3
j/FJbGpX9wle+7N8uLbEOGSRtbGWeExDYtOUuAD3nIEwMaHVLFGbnPPTzUq2UuUW17qG3o0sUPHN
EkrcEa5JnQsf6L5kAydUX6f3/sQtaF8KTKQTARRDi9Fbw96GMNk8lSKjQ4Cv3mtDEVIkWz1MH5oz
R0jYnsramgBQM0wr7w18Df660bbo5KB8TgNH1WvP3x0CZqdlghSTmVo9ffUDpL8wRZqbjNTdeAUL
ACWj5rsE1ijFYjImOEYMhsuusFh0rDSmisuAl1Wj1xROCqK9DRxhN5dxnbUk/2IVrgPcLkDctDoN
PHCl7HX6sxXNEcyVSmNQdNbAecECELYk126FAxh1TjBn1Fp6jz5RSuECyiLA0ow9UKQDBuR3Cvir
90EpIfO0lJF6B5pOcH6htv+lcL5miXJyTMmirJdYYs+KFYoqA4YlZJRroeq/jMzieah13drPfXVL
VvZj/eysYTJAkTZXgUui9W2eriSI7TDjevf2sU5YCBb1Dy9ueqvBDHwAAriQHCKyoARMW2oIfdnf
Rp7um8Rq2Yt0fRB882YPBhuZJMIN1MO+bMBKXMeJ0LTF8KVwV4+0yb5kdyOEhkc6rsx28QbrUw+i
aWYX988NV5Y6I1+sLVRqc7Rr1xGnbRoFnFwS9np6oCmM7NPERce4kwYuG7PEGOQvOo2KnSraZyMV
hUjAOxKEAyOJOSuu29n2za9i4GgKfh8B2I1r+UQIpbStpACG95J/TV5WhwDmcNBzqp9BP0/kYXQj
8K8i3nP4ri3CpaMHXWVbzER/haCl1anKlygPUgCYHvFHbSPhtpTswh26ZAG8dPzX6p/DzqRemXru
Axl6G2tZWb1u8cS7OAmQnl+4SVowV7LCz46j5iAcjSnydJ2vI3+EHGa3BcG/3V7ZHW2DePSaqV0B
NCSphmqbG9ehAZwGm2QV7Yb+CIyfVBBfiHTCvKVFwHkUqq0R7KFEf6GsPbfbTBNMzBOEP/2xekns
1MLveUs0rrra77KAxXproTdtpWx1qyAXWsxJJ0hgMepRm7rNRWMNk4Nh2KL/lQrSJ+qW31RvS/z1
g7sXMEhF/3OkqiWlUwO23eOfOmPdse704quo9G2UisR8LHH382p+B97OhEorNpRwOupK2jezTCom
vAMhNlqlJYEzQOxQn/ZazKPXoHVBDi+1fZ/KATZZR6Ojhl/RiEwkxPHLna9Az+1lLXDRccIjBLLI
zhiI926hwv4s87jog/teXCeDpP6C3loERFHrpUIHe3ro3icCEDdMipqSfppwG9ZwOzxGd3p6HMrZ
54Bm3z6a7ombD+hEnjq1i8PTe8e8PVU+xoz5uocCJrrxE7/rMFwGap5+OAtvGqcGrg9GYu2XOUar
l1dXlR+BJAp91jVjNWflrj+sjobjesXzuB3KLPU7gCOvsnxsj29NgFRDsYOAj/2TvAZTR00xIYLs
WR7iEpa66tsXuYWXdzog6RivCivE1CYjINENtxpniudvAOT1xu2TeeCcCZS/3zY9H5antSnXYXQp
IdRRs3EIXs5blw5PWj2kpmvjcWjEGZYQ9ZCy4giLqPUk+Nl5jzS0cHj8EJVF5B1aavkY8lZDx4Mp
2G/gX6LwIfSxOmAhPKzLk6ofj3hFNFVcVSV9P0cuBX6BMex7YRjG08yt6Px3hfgp5Wg/pSuHiC6U
F04eL+R+eiwuwaO4HzMN8vwOVQgv/xEJHkmRKUvozqDU1eoz8P0gdIcGKULj4KlChe3ZzXNr4NHu
MoF6Obk0FMvqg9nIu2OkBTkDEJS+eHiT6EbjeDwCP9EExcViPNMCAY7Ipe4FlpbyXBz33g7a5xnK
JTABH8J5VLpqUO1/whDEc2VrTKYpJt2ocWPNM824abDPr1cbGRPTw7Kkzf1YnHF/gbzEUceH7WzS
vhM94xcJ8j1JZV9/g8i2XmhEHOv+RJsVzec/5iD4OHk92qzBS+QdpSSof3zlAK12+eYf2Z/tDIxz
Q8IhWsNzEm+DPwjY+Oj8Z9qUiFUxlYFcwtaND+jea2yK5DQr1LcGDQOvuGV7jPtkCSlbVsClhzMn
HNUQ1SddyFQNRdgp75TJFOl6tgvGsm+JygFJKYMW/RHK4Gyike0EuVXuDdwvEq4KfW+fdHbSoAl0
aGC9cJFVLnqA943yYuR4WMQH6ZJWKhfzTeeh14JtCc4ejSe9A0UiK9a2UfCsTvEy4AdpqkCM8NRG
U8uSxJoSt42SIQYsWk6Ep0/N51laGkLyTESajDwKaEnBFVKmAHMqRb0yir8VF0mUvKfhojl2qMJe
w3Ohh07eFNnGOledwTP3HyfDC5ZgQhOCgBi0pXpE7PRVw2v5jAmIWLGXOA1UhayZd6gt3goxFY1A
ELhyuTopvBdrZpop056lqor0eJVz1rPd//VTPPNcRFvfzouxpvLfVEMrnTVB/pTCkhXBofDXFS/X
CGSo7CPbVZf+jhx2O56SJgswoRbhd7oL90L90r2i7B40imjWn/36UnC3T1UslHLQFbxcfjzugNXb
Rg2VSbr7tVluqSwf5iG4Nu4O2sVs6awYaZsDqq82eW6+PseDxUIt9ja2XSzw2HpseeOeNR7dqeG+
OK0yqD1T5+LV7fPuQow0+SEIBb2rFAWMr+KdooHb6fCzYcA7MS6KhrN2fGLl72Vzub/8XVVBTTn9
NG7evuFSySNHmBIZuJtG7LsldwOyGulPQwIcN2z9oug3x9FVOZUWQgpihdHvkKWmMaQxWZEJlH6B
hklZ/7w8o+AmjTP3GZzvTAMlHD6Eu/wYI/aIWUQI8cX/yZCDMeyfmlmgRfg07dhNDOIE6RGfVLFD
SbtAE7Kv1US6JovR2ReLicZMLXbNbpFtr8HSZ/roVeoDGv5+yRvPlYyh2Z3AqCetZQqtqmUnFj+p
x42o5V+09Rn0GdcblHUL/NHbh1QRpS0cMz+fC4nDXQFoCiTtx+t/gVQ0sIhL6PzxOLCSV+qXZxDH
CecK++g449oeWtWNK7kb5IYKuuXuQouAUoUJaadvDafHxwAy7Ih0PS6JQnQWcWbTi3JCNRsNwaQC
afz9Wlnrl4+HCLZx0WFzdbB43OqdY1K6cJdKh34GfUx2+nc2BihiQSOzx/nvS/0ASVpL2KaYcL0k
61p5OvCYl5ax0cgzEUJYNyEsI86WohCZjaOxeGfSOBHPYrTTyXS4lyWjFU42X15sPpfLBEtFPMfH
thtCK2QFxENE+fv0Lhfb9YIAX2jISTwZuaAFCI9Sr3Y0OfY2owYsu19IOqKQVzBdaIvToKELsYur
BhvYe8G0FriwKEopFhqJZqrwhKxUujkWaAVlt/xlPi0kCUMQF07sZA5BYIACbepPx+TTg71TXdyY
4RFX0XMLrwzgx18SLhvAXsYrijZqCq5GE5ERv+DO2joPtVJIeLtrxJ/GoKRSRD8fBwWMXJQMY6TL
DUKChStjFPlHidWNXheRFQ1/MhdiemHlOjrFD3UV79McVgMY0ABUiZ28bVBPRsYo8ecZKgBpZoiN
SQEKYlv9i/mj6EEutR/0b195fb7Ku14a2XixWoCiXFCbUXiBH/UFKMpqQkvBBwI1WJFqFK8mtNMH
ZVwLL/tKIpdnOr7mCjsX7qAdOtrZsIoxtZA93yuCU+yt5QtwwQtKrLOPfLrlRJNrxtIEufrxhlGm
VGy48wEycf5/ma8enlRWpfd857mYyUMmYm4sSkY88v0NSZiBAZlgrICuOTjZN3xQ/dn8nwgJIjkD
WuJyjZtX5kI6EY4VmFhb9hXGrMw3DVP1tpz8ff3NKC+36KnToYhaS286yteNdZirhixMiopB7azQ
C8YM7SiIAxnpuvKeI0LVmIfZj3/h8ni+JI1uP0tsWZQgxDydInj3mYgmoPCRzQiPpIWJDcyxgPet
1wyrhGE1tvgabcb5wsW/hSfQu4mBLHtP4BrRsNeE8w1ukZw6g0H544OUpb3sDEpWOM96mKBbcmse
XnzHHhYdpSUbewXX15kKb7qvOhVjy9n4Xx0xxfrkaC7esARPwtVPPGa6JPyqziAciPsSLbgVtVcU
1CMWsmQQPL7VQ0g/Noe25p/tLFbwERrB3A+wB28n/4plSmR+Z+8/tuZ4miT1VkMC96vyybmqXkDu
VmcWrWY4ukh5DbyAy0Sb37yv33CxsBC8X2V9qXOZSyte7c+xpCyvz0Rvzunh3NfR6AwQAaeQHjDx
WZg0sGBP8bXE7Om4FrzDUg7nufQWzea99oQ1Q6i5enU+FFkFPu7CcwIbsTpYzvcfO4D9wWZ4njlp
TM1mjwxDrgwLtV7nGngMERNhM+A3fEOywHC3gX1Le59gthfstpJHYFeNeK9WuS3NAEjqdlfvJa0P
095PwBx7gU5JSBWprOAzpGnLC/L5pZKZyVAjUtU0jZWyCzPBxRRxrtplp8EkACYRrV4+ozKcYm5j
iaYu8uO2iEEdDPJ0V7xoYtVV/msNo95R2swhcXMk9lxBx7VgI35S2g6lcp67JV+FOsbjP9G/VCJC
76TXvZ5XM0La7rFDdDYMxBu2TcV7dWvtRKvPuwnliCL8IZbVTbW8Py/hOr8dIpDHmUYWjsyqs/C0
p00S3qQwZHjY5G9b37PhhyXnRX31mGFb2nCk8QfLU4JAyFUo41Xc+BPfjIUnBpWfGV9aTG4wiS6z
7M8rqdZYEQBM+H6wphNZYhNeWZ1NVCd+iq43tMNm9cBteL8uLk9Xe4+tJpAyZiZpRWkZPRNJIkCA
cUWnaIVo5d6MM1ojOGjuP7XYyb1f6bK7fCPkTss9h0mRG0MVPpd+Ex2tYZjpbU96etXfDP8UIzDt
aJqjfcB3ctMKx6hww6s9mohAWOSmCVoylB8HtrYaU5hFuDG7OrKEiILcpRb/nrtvtygqInqN482a
sSbSMaG3L180UrZDZepzQs6bCckLholE3DIHvLk7HDFLDzP0JcHB2fCQin2NqOaaAi87XkZZPr6f
sW1kL9FX1pKALnwkdqgEu88nHSa8QYM+ma0Nct+t/KRKkNeWDZglfAfBaoBwXpLmtHxep6vVAluc
FDrJOCZS3X4mLDkJOI9tfdMm+hsdqg38Xir/4cAsw8h122AAF+lxUBxVjpAuurFpXE0+R2s2Mk/p
8c0KY1eqcp6iPY7sOcvSKfJpE7i6I5gnHVLS3x68QP25t+7pghwSQu9jDFbouG1BMZ80uBAk7WjU
Dq6FADAHwF1ciQuVFMWVU3y3+vh2X4OpamzUfgT7P4ZlH5XXpXqEd8YZEV75LhtuRxdIJdBVrW4O
zUkK/OjpNv0zZml+6ItsiwF89JkJmmXGKYRk0TYSXLP0vcNI/V3N/fWVV7NqLLm8vZIf/3VjFZuA
AFahmeEYTBCYBNe/nhXQn0Y3JoeiZqp6gxSRInCk3m00QdlWKA/480KhZc277P5ArwAQsRivHKbS
l8r+ASLO3xaUfe/QG5q0Pkwg7a+XzCcSfSpMTY2cysZpZnV+OEB1tps2h1zh+Z//+gsQhjNKmzWZ
/sjEbPTgDwwCbHfTGuRilKs0zQqISxgfvHgUkOvzec5W79VbpUiFx6no9CYFmpz1yc6vv0NTw6Z1
yw4UgE5lej24Y/naM7NBA4Q0EFDjxsWWgtZHgZfYcZsdvsPJjbgKy1f27zaflqnolxiKzT8yXaCj
HWV0JskW+99NFggWaUl/QjrbAzkIZRyT1dEQuteCAcUuAt7UjI7oNOL/luNlYhygwaXT0H67L0x9
Vn1aLu/mXawGIHYhtmHbBnC3zlgoAWRpQ6PYVWA0LYFmPrtV8fJj0TKW0+JkDK4W9VhGyuISTByo
rowQHI08uHbdwdOGdKZfHvSzmivUMUWMdROU+gWfcm4EWXnRIUcAaSEmYcgJyrnM3Mtx4XU1lBAp
lP0QLZF7WAPSFtVJigSxceBC0xp04p+pZiKt3tixC/ia59z212gjORboWZvtDHKTFeWZcEjsp/0I
eT2n+tiRZCFXRqk3DxfE8zWtG4I0QiAx7mJfk+bxWiY/6ZvKDUPbhxwwFd03pn4iq3xe1PQQtXyj
m8KiUg13d+hg0YAf8jI+923w7f/5DDq23WstwKBHJ953Uhm8E3A9wgionN19W3H8rc7CfVZ9/G/8
3R7VE4au1sn+X4SzY52nlOUc6IqdqLwn5GwdxYI6Kbjgg7X0pM9c06Hw8KsARMk4+nx3413oIww/
PG2F4Q9bAQoI2NekJPcvvARqdUsL0czVgftq+vOTALErdPq+UOppDNlyGKn+ZVOoQT/Yk3m8Fs2c
fFYunE/K4p+MVQuXFyk/b/SC4srtWaM1t3ghivY/selcj3yTmUCdp/PaVwHVnVPVS5IqhomQNxz5
OiLYrspqoI5g1h/AmQnxlj+IuldwIE7hj+sVHyJorwan1CdVFRMkf1qMCO3Fju9bdWOkI/ARXkDn
5Qw7AGLZVhcgFjo7L/44mJqiuDyKVPJ7U3ZEMc8x7spHkB7fKx1Uad2twf3OvscjGeXOchOTvOS/
b8EK/ayMyf1Cq7qJ2+zieenbOEsGbjUD/l2SHx2DIS9Ue8JudC6/OoS/Po8ngg1n7bZE4RExkjXf
yoVQ6pFxYcA4wjt9cIBjgaTsGeA+9kqKb9N9d+TSUZEErLcq4r8tS+9K/IN3ULOoYexxn8LRI2Z2
gToVwtKHDvN9TGawowghmTpIQX4BL/KeUiApo2MH3aY0vq0yxdto1AILHmYMhve/9UVTogxBOSgS
D4M5bxNuSBfv26mTlOm9y2p/0MQcqNEmNkIeH0ZnPBGhWl9SxWdincjb95+s0oFN1I6U5De4mUjU
ZU8ibNegHWplZN2Pamcr3fsvn5DbcaLz/rqlCIjjs7AM/XRkztRLi7A12YJVEN8k3o/rcf2mmaYa
rKwj0hQvQwO+kTAWasF7lSvcZm8WYvQMhqYVtDiAjoD7iMeMg2hhBoxpkFO52BDUJban05up7EGf
J7kRDoJEWQ/p1M/860yFmbXgPtH2fy+CuXscVFPy3kS/aIB/MhNdEFBkKcp5+KmYojVDb9fCQQZp
XfrLer4XNekZhWVTMi6y18PLyjQGmSkB0zn/rSVWwMpDPxZMGD3KwcfdSyMmZwKXk80lR0SRKisE
hfp0eKv8P1R8CN3lHJ9SjBQQVQwkepJszQqBq1YW4lZSgl/+NAgGcFVcxs11yTzpN06mxt0iYtu7
owQ53L5MO9+l32dvNDHw74b8JgpOCjl9Uc+jQSssgP1ez2fpoIHRGdYZPUGTR2CMQ5JjqCn5LwyF
nI26qunVoB9vUiUWmiZppGCsct6351wVps0wqwpNFlh9Ufe77vMaVfHRkTKCxMLYxN0R2vLGG1gN
TEjQS7Z8UG41H1/m+Sl+wGL5r/tnuffsYdM+dAiJeptVSUfh/PVK/V75tpRjnTfyMA+1cNIitnkL
Zz8FQlvqpMT73EaA2guhjuixG+y4ZaiunisM+wgScetFRcL/Zmt0U2+3vCf9WgiemWuw8LVT1kRK
Pgbot3Ag4CW4+20u9d18wekNYWnITXBC4LoAJU8+1CE6DAncsnNX5YBshpg9gCq4b8KfovJLKxsB
2fQUQTMeOrEdfA50IIFqUznLZ55ZVAv+j4VP+aCgaNbckX02ykTxOC44/jkG7FL5PcHGUgHvbc0P
LhWlGrtv0ELY24d56OK+90RDNtIg6HLHIvnGwFVFbnTBNTvbHyK4aia03+FUxxZKVl2OuIZ16Qsy
9avbE1RN2v9z65HNJp1n3KyLokeyhfF3A52ljyeQs+oE+2HMO9MjKTi4D/TDjEqJ1PIbPbJnedbX
ZYcBhBcJZKjBYPNcoJAQ7UDKMvNt2udAEVMBN5lGI14mcnNjPjA7t40Op4SwDWBex0HCaDd1COkH
GRG6iWUeFqMr9biaSt4l4yYG97BsM54Y2ctZEQ9849zHrbEGLgGI7C24G8PkuAG0hHFia2tLtISb
SoR395/k9cvUEhV/ydMvTq9TpINBDs3+qzTCKPZnGAgvv3qLam+9vliF0DjyuczMefMAlxjdrwZh
QugUE9nKl/7HDohTH353XXUUnAhyGaEAQ2A3S8jfu++sRox4ipJkbeY/S/a2ACyqj30xdxZT1UOB
Fq0lp0HOD2QblI35uPtgK980iALLpBmLADDdKRvyVNy5GRikNsA5R/8j2yDov71jKBhohwc+q8My
DMhkVylEtuAmr9CQgUtWnDrfchsnjCkem5srpUvXWy8SfeptBPpT332AuBtqXF7y8Ax1TiL+rvWD
wDXG5Iu5DqpCCpoPReLO5+Lkdmalf/H98MCLxOMGgvVqG7+11MhOq8ZZATL55I0C7qUSizYaOFJj
jNIG0C7THin0pmzhfK7HULLFoq9oLg9L1NvonJk8a5cVc6ZIUaAAYUWY9Rt1LHgKDZcHD5xwbxTr
nKYxvGpJduCEokzOEYp5twHQUpG+Ij4+0wasSJTGoNcWQrAwxQuaotpgKKfTljFsJuDaNxALeVkG
0L/UpmRb0Wd6yC854HOl2Oq6OH+sfqMOItOxv6AhT2Ckv44XW7uccfqCCH4arHZvMrZiIFLXwKXy
U5rVks3LECiJQ+CLegIT0+pzGFRCC6giWzKP82YMgstaULtczZznJMK0fvrUlGh+2xrtbCYoBXZF
tpUkNbc2aNjh97VkGiEX/3Pp+9s2K7aGjrwbaiSVmIe6/5+hCEptdesErHCF+RsnNh3GzN9MZrAW
fodil6rmRYedKPYwCxHI3m67qcY4cZHYl+RiyQwFcIEVmpLPFWyXQKh6X8NWaxT2NVkFoaZYgttg
mUN1iXAFPkxMxrjqUlRT1DrZUO5L8J4REs3+ShKwPz0Jhxb//hH5V8tM4EcC5aO+J6ho/Lc+I2fd
REfHfKnsQ0d1B3Q04KEQyyI1paQ8FWfdsBnZtYu7vAbKsBJe1MGKVpAIZ2NWDpT+blD0Fbt4K1Yj
8j7ht1CLTS68Ol0/shwbpj/xcArrN0NlbgwGpUn1OPl6cTOypnLbpwF8y1Mvhd15ibI7Bm4dcroK
eVJMgkszMr6XYWJPAa1u2dbeem0cP9KoelPdL/UTLpMOeVTG2NQUsbYU3cbjzZQp9xKYGV9GdDQV
bOjUNKuBwPI0qNitcgiGmhoiFuoJoXQOeCul+r97mg4g6ARHP90uKnNqq3H61XrBfJjCPgup2JyL
JhTpVz2pu5Y/jvVSvTxaE84AC/2Tz51k3gj76Ngvz2IR9O+ti6lOsRxA/RaKjB/mkEEwcGc1IM5P
5gcNm+lph2vbpr6qMEwsZYwfc0Z6xevBd6XruRFZoU2aIIJk0bHx9ulUvkqLdV0oln5Ws/pX5Oo1
6/Op8PAiBq/GZDYPLeKLbSti4irrK4FQntXw2RBMj4kRnb/puWdrYd5WbTa8e4221y1eSuCeMJdg
JSu3cUrF3Mlu4hkb5eQPmbTQ4EboajrmG5c4OvfeGiqJtWyEls77oX9lo0BiVDE2YrpFt78P0LBZ
qLfT2NOdHeTPQPfRsUcKgC75KR8QAQpqUmBwa4N6c9ct/CZC4aveLebRRxsQIrVytNV8D9/FxtQG
BD0qs+XeXH8RiD9qHEdM6W7Y6YQ5CARw7W6eRPg8VYZ58G402x0wzSDHtFIWpDD+Qg6WcSkFH5iJ
FzC+XDBEx4IifF7Ao/zym4y1oSgC+U0i5eg0HfBJ0ebczBEUfgMIqh06XtnIWvJ7uT9cnYH4dYH4
lb0YJ3FHQriCAtsV08wiSSTpiF2BKtaFsiblaKRQhqCBktWw7ZIg1uCz83KjYF88Yr/B7YNOWWP4
UraN4pdgEUbEcQ9Tf3464CNJtpDGeBNbZZr5t9yNkAAjUtHhJksxIkLDVRjIRd4JCWCEvXEMk8zD
auG0tclog9by6XzMT7zmoAEozV1DZytGCTwGvsFzqgc/iMgQImbx2b+E2ApZYfFrptJvtQFNMgxL
m0V8fhmmgGifwkzL8H4eZ/VO/70mv1MyG+vloOyXtV2AJvYeGCAisnjI0m60lfSKCXykfce5Anlc
PMwRagyST+uMRjmTqt3c6Bf/d2raiRBWKmxe8nCFytyxP3p+0nj9TOCReRKBedyVNdO5x0BC1z+w
ENm4cneiX4L2ksXyYgBo9OEY0JPU7SGFnm/NIVCwVPrZSnpTHyZbGSLE1x1J2bOZe8hjSXS/QnNe
HwTLa6cgd0EPy/Im+qULn7qoTAH0J5vekEguolWU7Pqkj/fha9MSa+XnSDoz2/obAM0AuxecwLpn
WmEU3gaggYtmmMoQExPQIRH3FjCi9CtT0b6/PvNVBOmRiYsuIU26je62xek0lLVuIqCyNE4Zs+XF
NkF/CwbrDEYx9gY1yfraAYbw+5o1yrFFHRsfQVpfmPdOcpEo0DbUgYW2mPb7DBw0VdiUWhKUKaRY
2COe9laqArtJQuieln2WsVTpJGlnn5KSUeTZETRJpUH07Okf1mY7y08HPey88dddbA6ZV+yQEzE4
DNauJsF68UI6wtAyZ2SQg/uKXlEjhWeJYriTgEpks5B/057fQjooZ01FAxSxFnihcnGnVWsz2Lnl
XI30UQ46QCsisGhGEZtW6XifxTEbd9DqLPkdXdFHIi+A0/pl+VFRL6SV002u4ZEInFzMeLo/I2LG
zXVLfLVWEW9nYLTAXTNw7PQsMzP3ViqdBSriY1P8kguRjdzmADN3DEm7tsf7gI/0UlJLRknVfCkm
4H0wXmeg/lkcUT8NFdm0hTajM97ufR5/lUO2e4OVyByTkg7BjBRDvOGcr3CLhuky/R/P9ZqfMv3D
powM/FQ498vC6yJZqwtF8QO25RurWD3R2jJk3XliXjUeokI57tjGegHJbKrktEm7eM/f7b3JaPbM
IDxA9fAsfdES5zn4jQnnnudo1FA//Rr4u81ji6cde0A0IFmMjmjAxyhYLjbe3bpCUAVNdkhz4KCP
DXTgJeYq2E1LiZD7xmnBPLAjxiaL9YajP0e1qOkmq3sf5PdJi7PlVb3DChZPaAitWGhiC+Z5UfBw
pzA9TWVajqZt8L4E6+U2/juk62TfNz0/kvJeZ/jZnPSOylkxte3o6UE5wyS/pd19cTeS+3IDWzRp
hqZ4hMNH2vQa7+JZyllrYUxTWF4d8w4mlX/DxF9QjGa3IdLrrETmW4E5c2SZxw9ZnMMAL7+hHvPf
P2IoKteEbPPQyHrUaxqBHg+MYNJzDO5GffBdheanu3rC2aiTk3OeT/LBVe5/Jh4SjOYs3ukmJ3dY
vAj83YJXwHGgGmiO64fktS7Tbra3Sudg/o5BpmEVjI5CtPD4z9VmDXLs2FVhJLxRSFuq1Db+V09t
Spvso85eeS0R/Wh/ibPQuIf7jyMEbcpyIXuCuLuFhROVzxRrBDNMJOETe/0ca0TIa7C1HjPIJzoE
nyd+h+qiVrBGhltAe670q+HDfyXx3Bh8zi/lEqzS9Xej94oDWoG2S0Ehxay0oPoZBc3VQOYY7EiY
ZAolbmn8ZQOnLI+hlwgHMHRfWQTa+vZDrIwf3Bpvgiit7H+qHu5HBoITKURLk4c7NB+0OpjarB/B
Xsy7qJRR0qdfskt0lpeG/jZHs7DSc96tiCpWozIq6j/6d4vOeNUrFNTatx1By2PHGC6spzhcAEkF
S4Hry2LrXjM/BUsjrz4C+ulrs+li+Wiv6pfYIMUDwFn5pnEBgRj0d3GSWBLZjKyFa8DYKVd6JCTX
TlOuqyvmV7bB5tUORtdoZO4La2I04oDsp4WHuKYPiS72o0JmRalGX5v9BB6A8ZuogUgYXsyDkNMW
hkQQywaRhEdUTAxxJeVcjQ+cm9BTi/roIn2A6epMXEqye8hCA1d/O9s1E+147MSpgAqosL2+n2o2
mZMoQRuQadoU+iMKxzlqWt4e2J9SUU9zvZnwt0jIrCQEymD+t+7JMj8ML8QqsoGkaGe/wgBh/FeI
KPbR9bIdW+qwwO/zTZG3GoA2JGKusD0dh2Ss2fOKSCSdbSBf30Mw3RfnckF6z9GR//hRPa59tAoo
WimhskeVUJY6SNE4snaK8M82xhaq8aFYRWhRogRHfIpIYEeu2WKZM2Ljwn016yTYASexrGBztBxu
kE+La7FIXd58pGyXmjzGGhbUVVRg4cRjed+FWCe34BRu6yjUznJ7JWZgTx9zDtP9JgVfl4cS9PYY
QotmPm1TGXseE/A++gxMIE6wpVaUNwKYW0vvJgA6YbmNW+9HxNYwkma6GAoL2RSyoAKrVx02uUav
VYBGgWetL/gz2GRYjLGu5LTAgpry9XAjdZeK5bFqWy5M5tMOUJZAZ9t8WstsGxYdcq4fLJpCgbin
1iZ7mm+KymYeHe6nn7LDc0LDzrKXYmdAmKWUhizHpfFX7loO2Gdkup6meMwtY8kzKW1fXPjc9mcz
ujwX2bgu0U712m+5mxvOd7jwlkBkhUnynDIfUvVi474hRxCUA8uA7FSDpEGBHMdM2A8qIxHRUMmk
tlqzSQtdF/zjC9Q0Cm1bTiPUH4Pw9oyZJuAEceg+1vw4qMMAOplOlaamSAkaTenLgsPCkymDAXld
yH7ol81pa9kOxP28KvYF9lVB1/xhrFWgZ8WYCAUc+joy4jcSdo9mB8rArNr8cOcM6sbUMr1qh76w
9SKw2RS4fqF/yCpwaFSvL/BjQpxb+JPMH+pcft/G+bkHw5ktFGeNJSP0flSZ9Ye0GNu7OayhJbab
sjYcSXfZUwEK1/ilVocXPLYk0xLblSdb/y3oSf4LNjkBHcbyqMxRj4h0HpwmCqmuof8jV5MK/pCO
r5I8Vf6abDDNZcbE+SDeHluf/B2cQvcOoPvcEFRjFaphGjDY3KkNwJZljjrMI7ZOs+FK8e9gN3F3
hByVdGqfb7i3aBZsCS0wwrSzYFWy4X7VFrcIQ6iWxEIHP0LMmFv1cr8688vJTt1Nv5TTFij+fl+H
F2ysRpkHerATgh34vQ5H6cDMcXexiD0/nK3R32ypun0daoNx59DBBjXVP3fAkDKho1UtRaz/MZEY
4gY4LLJtUAcDzwBqyjldZfEcihY/RvCYvPPE353zFj/6L/5i3WbnBFD2NHlykTKhSiXSXn7PENdo
oImj/+yG8eGf0JV6Pzng1F+YdM3HgOFLiivMz6qVSKrKKENC3FmznfWl8l9bRFVu8LTDEsuYaLEk
XtmSkKMi3gcafsk9wC6XVWYUpT3PZvrGBkOWDpTxto3U0+mvXfmsU6KsEhdy3SpvmCJDrd0qaJUm
/22vhLxqolWS4q2Nlw4IryQTRZchYdmvxz0TxAzSS1kb3EShsxUsOCaRbMFSKndOXZTOww0BDD4B
+JQHyz0C0Jx1uCpBd9dfhaXMt85iKt1doW1mndc/vXS6psdmyV+FRAyzzT+44PST3YriWazx99eF
gCwYzimBRzXin38XLUCdOMUR+ZY+uFeeVYKneNqTYeYBkCWLBKwk2lh4NuPEkr8U8HOQiYzZGlqq
MFgNdbyrzj3STvKSUnpFnpGh6lHl5kpJYnqfcf/vSqndSmpuXpHSut42Y0NLJY+ZSQZZyzDemIRb
yEZ/KSPgLggHtUQuOEaOdmNsnIwfHIPZfxEuarGqSXPTp0T1RNr12dPmqAivQwgxy3LqurBN9lLC
Hl8VafPu25VlSdygOZsKgjUA2GHsswXriHrENRtNp40Gpi9MVD2aqP6GZBlznJp6Us14san40doV
H+flshjUQ6CYae2VGG0TkUYFr72tgg5LDoSLgL9h9SP6sni/v7BCF2Rfkbdzyfz55TmK+BG5f6rm
7wA3ftuDZqsyiNSnLmJL46Vud/kOyAlmoSQDPd6tWG7VdAB7ufNZ5V4BXEcouGI4/ETfsJNIK2A0
Fd+tr8knftjlU14bnt8nGIJDNoKx0obaqvRT2M7IuMGoa8BscrcHKG9EYJG+HxGTT/mcmNrd1az4
LSjU6DAn0ozMd5rnLk4gHfIsBkROipMsjsWZ+IFrJFSYzFMHFtQczwCmQPI0cKmdavY2PRmRo/v4
PZk9ko2imUPJT8UJUMaquxaM0/uy+K9vzHYByQL0hoE+lflwyRfJqj/mpaQm4xsCeD9MQscfQfgv
iFKxECkjLKdAXyc/6Vdwv3GP+7pp5tzLA1hUohuuOqheeuYoFdnVqtFERLXudk+aTw2C43frx20G
E+JQoDhomcUkw1EWFcvRV3j0+9Mitw07SqHRLjO74p2zYP7ONoIVGUQYPhJ0YD8hhkY2/95jK2wj
06Gpsb4qMBcUCoB5lxtjnHR7sogodIZlG47u2tOTovdS+Zad/xVjFfi9A8mdIBcsq8eLbIVH/wzf
fnIcRMAMJ5YyYWqgP7KlYL7gv9wReiKbBc6SwFyRXn/pbKOu7AJrUIHWtPxyz85Kiq8XNEYCjoe9
7hO4rHUkOem3AoPpUr+tCvhKosWKE2LU74wQd67Ee85+5eKG0Bh230Z6gbkCkCubVvtNNS+Iv0mP
slukFBE2ujJSu3ZCVoVcqZ9yCoahfqEyu3WTFKmS78CS3Y/w3fvRw6xQe316p8o0Obtc7nMXn4nJ
mzVuhWXNk93aks5kJxdtlZBr5BzSmWjXGssq2MFYYWWo233mZps2UhNqzViHrFpnLnvkhi/U2ZI5
kB0SlpjnNW/KfTVj2prh9elE+BuRWWCD9LHmeBeHksj238opVSjayBDTq4BC4K1761GNX7BVtQ3f
dUCAblzBRKcIEvi3cqG5a3YaDJL+ZMXtr9NUXbqp3sEzSZPAdK5r2ke+mYDxHkOX3ajpxXhRLWLx
hR2rjQE7g19oH9/tW7QFV9rc3P8d6XMMH7MZm+N0BBHxfa3KRcp3n+ApfdpnS8tdPuaKO8F2Nnhs
qya4rAZlKSny7V7y4/zMcEEeniQNg6VCe/x1/DI6z9s1wR9d+RER31ouEFN7Jbo5lHllVli8dT2i
ahR8HEvhU3YE1GsLsqhn8ChkGndem//dB1W/tXc9DnZruDEuo5dLV1abXUzj+u5l34qLYM6Yus2S
Fkv9gVYrsYxxK5DHoQ20azGJwX53noyIto9ZuMlYetxCjPpmQ9CwatZram3r29+qXOx+zc+gvniC
94eu+ZWL+Jlpe4O4AhqIpailY06xmtMTdFoUziqgzb1iDEjwBlb2472UdpfZCtPMxBkySk20CMAJ
iuDcITMK6q6iPvFjbt2HcIJYIakT7GZM4Ggu5Enq7ALk6kec+Vkt+iFF20Wufe45pR0oE3jGnhp7
gzArQ4yZKZ3bUXjs2z7aEk28o2QAUZ+XaabwShAOzyz6ksIpPSYAyDPvFIbmHwj4h9u9eiQkZAVG
ya4/fm/0H01mo5iLYU43wrT7e77qFDMDrW8G8O4LXZuSzj3N6f/xr4cIgr9oX4AaJ+eb6WlIZUt7
RKd1qfAMqwJbzF0VB9neAUbuahoBP4H2muudK0E1x9a4gp+9Gpnk9jfT/AUmXPh8W6nH9QsTPhff
uEATSwFCAePRDMwS0b4CIv4wkcHnLjbjIXQ+Fc58R6am0p72mx+JMJSlvCyfdDigrgMGfJuayY6A
Cpyj6Y9V+yVCSK/KumjILAiNwGxxzuiwrPfb4UaUllF6A88S/q9Ff8jBfPDCbx9lHzZAoBivAgvP
O8UmeeB2RHAAx/T2b4yk3BU2cibKZBz+03XpEzkAjEvb75tirdXsVh9z6o+XxHEo7tXbx1Q4y3Di
Ycr4Dewc6JfINDO/vSV6AuimU5fGTn8KKfu0Eu+slJlcfYi4lNNvb5/hNbWq3oEYlr/yqV3q5LGK
aub40oD16GnTeOWuAB/z6ALlQn2jQYrjtYrea0ngZhnuDcgR9bqEOEinIE7UFRst7mqy/5nbnJlF
mwdA+qA1jxEDzzJ5VmTrv6aQhggym1AfjnUG3UV3Zx6GSdVORejWfI9f/OPfSj1L7RM7nZjaP4qO
Vfv0Z6qDSxkwIWvq1hqOVSDG6IrP7zclVd4iVB3ORaQidrA7K/HN2Oa+0Q8XHPIcYs27ChsBgw1J
e7hrTyi/F6favEUsgLu2Ggu8esC8XqnJUzt6QbX71LJs9TEkoCfp8LTteWKfYsESYFtPTdByIgWK
26sxGBD3jlf/mULITaxgcnEJK7wlnH5ZKIE0EgSUDBq/ZLbu4B+4+HltPu8ypMdd61vZBwBmoWxG
8QArnMOGFz8OfqaPvPoD7z2HjixhSneoPJaDiWDJO6T2f8rpC70Tc/lXFNlWvNleIxsbBQTmByUe
AGaSCZGmf2xf0R0aL/OF+vukdbfn/ivRrxbhGqBaiTBnZhtWSHDBl2icHydQv/wHapIIXMcgAGsD
MhbSSpLCtQX8L8g6hZ/wPEeqSWxEdX6a2h3qVF7ucw48kiScUL9Kb2loZp3UzLXFpgDHKDdPGPg2
uIjZFUmckdXlGN5VPI3H3RhkFcPIGszXdNiHeWkcKixNTklS2zyRGqVks7wycbvSmWS+a2gvZyRS
Cq7KlbBzC4C5asTRadRivxmCakBO6gM5mbBp2x1V3zvDL8JZ7YQ68cdyCgjcKSbXSw44dNUVViph
+KNvjHbSfzYzPgm6IID8bStynbpcDY3Znqb7cN3zdECiV8V2iDlZhdOg4CTCdbnp8L/BR60zy7z8
KnE9yVBzmg9DSbkhQm2jwZ8kT3G2FQwz4x3V/VqzfjXEc7hj4qt8zx73aSLATSOPfIAwnyltj+Sg
+UaXSfzXzGTd2c3x1oSi1+zEUFz8Is9jHru9JjfF1FuDmF8gyJNou6iolrXRp5o1qN4reo3QFiPo
iDqWSl5snmE66ZxChFzNN+mCTtlAKStjhXMhL9JQtoNnMoCVHdoqx6GE6fu56g9BEsoGWxrEolVf
xWkbqDse1n8BfV8SJ8SwuA6Tegp5x/hv5tWwfk/X+AQZR8f4ZRbS3PQBtqyHsHkx9K1TV0KvJAr9
xhliTvxeoBkkullTG0nXH/5VXDjERSKSY96UVyakCvx1iNNMWnSeqTYNhs70Pivrlxx1Wq2gAXXJ
vxIz5Z445/k3q2Nva6X/e4J0S5Z6caV6KFcgF+MK7e9S2qSGYmFDPXC/5ytK3tXFYb3VuIQyRORd
bMueymWxRG2k+KUoPdq5zZWKjFmNvCRJz9kdfcYF8FoL4nCvCK/neb7A9x7xQ3nIA/F6WS2o4m4i
moqHkEil0mO5R2LaHv7LfzPIcLBJ5zuyFOAAawEZ/3Orv9NRtnsosk7VTV5Y3qiHseU9JrU9pOF8
yGG1O2Q0qbkxlgQO7yXNW5RXvoDN9QRLfauF+8fWda+4w1ZBnXtWxzDE5X5FMFVgw1XC+ILgf1MG
m4+pPnVgnpIaQH4pDmD3fu3iDBJtWrVXQOuXGO9T7a2vDMUK+sGCgLsRTyjTtd3kZ2xDPzq+pQId
SyPHF69EqlVnbKdG04T+awX26YbsUkUnxZi4lhN7kfIsuRzE1/bk05rWxh6SIzTyk70OCN4x2K4v
cZgJjaSn6yUAJNURgqCf5zlcur2NYHi530RALMj9CWY2MvkezylzOxbVOw0HJKPF4SrciHX1b+GJ
YvFpo4XvGaeLFMB6zjjrmf9oWmG7US4nwst+mtxsQ7Ne/k1amvxK2eraxqkhG6EIM5l6b3LsdY5Q
NCMgwyLCfRuod1++SqS0PsmFAOaGkIiRDQld8ty10MbjHKT/bZFnoI83u6251BbHuYqPr4CHMVr7
cqw0EGVwmJhmHR23M1TALdTlLLq4hUbFHv1XCId/Hp1Ik/7Pk6dTSLwFYVl4Qn6vHCmig5VGE+6I
UlfpP9YNXaJeOnDydINYUhUD05bM3OH0DviS7+RfnOqcD1VsyNEdiNMuEIx7oTUHpZ9qB/KgYQE6
SAbl8JgGxZvr7GbCLROvIf6kf8SrlW6B3QtdEd48TFo2HF/ej7SvHsMUvCJxMFBv0mlugKCQWnIA
jB77XzbNFfpKFwWui0iOHE50/aTMh2V3AQmrPSYGRwT711UqTezH6ETxrGikF8D+xG14cgszyrp6
s7+LoZ2S3s8NibSz2I9jNsRnoR5spUslcF+ywSLVq13oZWpad9A8SOKjHq3t73tPYHn6TDOP2U2/
q8qD1Ucy8gxuxZ6bqpCuxBqwEG/FwhGrjlgHu3cxk1eW066eIirqyO90GYUFLF4iqM6c/Wfy/QNA
gBOLxsQW+gvxHSxEUypWnYf78pg7wE3fQxVvcRv7VLRCyzVFTNnQ2eHwN0JkjUkAwOTen5vycWIr
5u+uQI8e5Mgy4er/doBjYYR/VC4KpxGdAGE9yyTqiZZsvowUqkrdknZrdBrE7kE+9uvv3sDxlclE
wk73oWqfMSoJ1d04ZfbdRgzSgn/U/ZyZyJBBGGhC1KF3y5nb2hgehbI1DkyvvaBKOrrtW/8T2aK5
7DAstqOIQYsfSVOnnoAgWnAld0LW4T7QWg/X2f8YY+HeE6kY+PRi9fW9gLefdRy04U+jnwT2FY0t
YvRkoBD2eCvNZ74UAKwBIZi2sHx/C5tdomk3Aopea3E+UxW2r5tpgSYKhT3uWA+oxquyu93VM2ZN
jGu/yjab2kZmNhBuY9u/b4iwGBpRG7kUXa67BMF+uZ/defYLIebBxzEiIWDInL5D6JDpwo5Faamj
0EGBXXI6NGav7icYbhWxHhuIfGBncAqzZD/r8SO7a4h+G0hws6N/TZcEMiffTmDE6GCK83PKZ55Q
YylSMSSm7g5CUHH+sQg79V9qLts5uqICCpB9gd2aoBjv6EL6lDym5973B+KdVWUCrWOLQENItIWw
OrhnjveOktvE6xUKq7cSO/IaKoH8J8pksPKvmHOuHEuZl3zUoaQFTWNaCC0/D8QJgFJEwE3aD8gY
T9SbFqVHCBGaEBYdgbiRbQJLJImghR1gxA7shtnwZ61meRwMoMHKT3/KXtO1aFTDGyv81Hnrf993
UofwdonHRT69AM7qc/YZmctJVskv8Wl4/KMzRr4EXSScKVPEMgQ7KAaAPUPdtxHPgRJ0e1fDkrBh
30Ni6ZiICkdxFmoX6qVrBI6s+tXRp3eWiqNA5MDHm2a/rXCPxag3y9F0yUdKqv51QGWUcRvxjP+N
1vXdMd6pZFWdm2m/SIDEqug4aqTv7VCe0bz+HlJ0/Wae/QKqPb2Cd1doqcrkT73RqcDs1kEqD5oN
kmJlcMoMO337cvWNK2l5+wi+UfcGAOuKuwH0ZgHYweyY+fgaV/qI+O0gOq82lSRhDtH6lnoB2dhX
pk/AtvWy9fc8z/kUT78Oy7+hR0d8G0mczCZlJCTBbIUY+/xi2QVpmVcRM1UDTm5km4XIyzhMNqx7
Xhyh+0NQT1lG2ZFhO1prMAMLxprza6xBWKPLPocYWpYxs8hDM9Ps2lUaawlTOhuQRh2u3HBZnnBE
qoQjQfoVpxeOLqI7dByYt82cewgMbJUKrS5sidipOehXHQltAAM/gE49iy5KjMP3VgMBvX0wMBsL
WbdWmLnHwYWoX0GWt/qtW+UREeHAPkYfs5iN3k03QEwuYzYO1WXWwsyVoQsKr0rLmKJSRGi5uihi
AMYL1VGVHZTxNYtCjPFueaOZkkIQaZ2G5NBZflra4bk7Kbaxf1B3jk0lrWu8LvbXa95SnfWo9ZFW
fGe/Ua7CtCcIgFI7JqofNblxdyuR4XU++p9NECpDprBnWk33nVfqT0XuEPsVPKIw8UkKWAp8YIt4
7YxlHN0J3V1nH/DDsagX3KX6Nl5r9b6tgM1brEMlf+VfRuDiCUHFVjh6BCdz4Ux7O97NDyKjVaeG
RnSczx6iBae9wbbgO3sv2G1WUT7d+xzQoayShXBn6qZqiwBN8jh41KAovTcGL6mlPgzhERIGHoCg
d0UinBtZhipWZwGle1jA/y/ZogArXPH1QRRRWgokbSPgZx9t6wKMvErhw5A44s1hhK63r/esh/yF
TYjIWbkYvchmzMZkG8RAzn/Us7+psC4tEPtJdUjlBS5kSnFe3nEskN5A8E2s7Slc5PuP5uPj1seL
rz9EqUGp3k+L5OppgLOKs1gpD50jeIVaJW7bfD1kgPpncl+vK63nihPsq2mImqy8fKLQ+BIjsknA
CmfU4cxB/CDNn58ejH46klRtUT3NFHxWI+5AYPIIqK30oDvmK+ai/DyJxAmq9RqHtRSMAekdJ38N
8zbI4+ctTtIRwGqB9cPcFNCihz0uG78gTVhsn1JAOwkKg3MdY1aT4oMgNIVgmC/KnpxQ6pdqYxqE
Bn7V4roIDOLmRwqxXwgZMyItYvPkSANS14xHJm9GL4Vges2MtJXgmr0zswEX255OeL5G7+QY/j7V
EgN6aeuPhgOuIg0AHxNU+ok2b/lBfhlexViYYMKK8ugfXNiFqrUWYJCK7aAXq3256GKJFifrMVdK
wAlplIXJWxZy6OmeaYpgrQsHUAFRUvMmyqk/AI8EgwrFQ3nrvcDNUAOR7upoK9GxEVnrKCH0Y+EN
CAa3rEvqYet6cO/H1Jbt0gIXzvWAwbsF8fq2KeauHhqoOIYxfZDLK1qv7VlemDzjmslMHR9fkEY6
OrEaSr+WZmYERgjt/1i1QlkJLP96t+hpEIVDyiDnMn5o8NkrbjJr9fYmikbnZEgFO7pzif4O3Stp
UmvHZx1h+18y1dFnm5mLExswcw1ogQRO7jsF9cio8xFcGFygvOwm1sQDPE+UuF/IN88yr/AlsFuN
nPkl7vL5akVaGGB40HesqzdDar8Il4KLuJQv3hP+DSuuT+mYMOGT90IhXzkcqjezoxQcNdgKdyba
+mYw9V9TGJ9eH7BGUuq4BUkDLGDs709ILHQNTHB1hJhyDISs92G87FOZ2EULP0vz6QF+rLJTEjCH
LIa1ubJFwqHPylJdBI18GUZU0PM9YTyAjzxccAHs/GbDKb+HVFY2cGr5XK/bS5HJlFlZjmULpEXs
6JTITtnyDxak0lTwDmZ3Ey8S3HzU2eBGwGAcHpLxwqO9Ldci0bMIChy4BiJ0segbeo/7Zk3ka64e
Q/j/a2rZuOUjE96zZEqa4Q9AEykimvESVL8rZd0OK34djiSQ5SzA47380nMPGEilS6xEPnXUpQv9
NjpinvG8ToAtMIK40ZrRb6vcfh2XNytC8ZcZO8c35nDpKEVdyxz0GfCDiXSIkZ9OZM/yqkNHLmpo
a1gUGTvvp1dxWo3Cjj6vhj2V74aVfFosLvgVXRib7UU+ivBUsOUikrwmCSkT5u3/GPRYHJMwzUvW
pqAmeCYUUEUwsKNy9J/WucguHK1g2vn3+vIUFFtG3sOC6lNHJ1Yp95nM9GjFvyBXaicC0M0cN50h
jMSuAelRSZ4dhMcX2J+zU86asQ5LHYvtC1N3dmYdzQzN7/TZk2F+nN2unLygUMSHyZYPiTNt9QFc
cfJFFOKgEsRWGiiReXMH4tbT69uUiuQkcfxIVYf5r3sJVFBK8RIf3bonWSOM1HLFj+BFQ1jRZOPI
wWfsYHT29c4jyBycH931shakTAH797/Qjb4YcORIm78bT4kWQymjXZkOBPYcyziSWVzm8ax+qrxT
3Ud/YnLy3TuJljbBfmYqnK/SGvehyc3LvgItCT4ZojQq6xW4diI0UPkWtj0nXDZNH0wH4R0JefM3
a+klpMu0g4/Kk5jYEueb4MQUffoovIB8qxLTrzoM/XR9/1PORHGrf8a0lBJs6YN4DLYlYdDSxGfn
VeS6QIBANbF48/BTmPCDGMvJsMN5cv17NTFLyg7asyU47JfJCyV7VpxmXDkxlNmqAt2PtY6ZWRgE
v7VlogPzttDuEqjtiE6W3vat+IBDhnDDrQjky6JfoJSSwONU698tpvdQduwMsS8DZRYsfVIh/xcd
/geD001o4i+AYdvAHrk97oNuNj+nwklrWPBCe+0DB0Ujhj/60bTuIpDcLYhiJfHC5YKMGsiMcUP0
1J8pCmUEmyd7sWe/s/br67wjVAit0WpiQaLGtUyNIufjqt8+qive4FR3uRkv6LjfYyZHL3AldARZ
p5aiN+HHy5CInzJtSd9ayL3XjH9MHEjpCI+7DalRyUqyQ1XNEROMGbxNi/3bSJAkMBkn+JMRNIHc
JYNc5vzHBa241cb2cPDSybc7xShAtWYLCJvzmDXz17X4eafv5+D1JkZZF+GPYyz9xv+e5YZ/nmrg
7vD/4v/Ar0vc+6T7pAhbnp0NVc5gJHVnF4OeNXanQ+coMIz42+iSixouZCt3DRIFskAlDklOPlMw
cvJhG/s/HRkIz5/ZPdaCGPoveLDTSXLi5FPeooLFnpgmZNk1lZl2nNockMMlAadODkXxfENsr+aW
AEJIBDP2FpJ7MQ4naj0Fown6PX09Bzrl4xgm4gSWzCxbjW3CemklzmCAgM5nL3u3tp3JyhRd5REU
7V/eHnr067PoscfjjxSrmPVwoqEnQLNswre3k9hxvl9bxMaQBTVQ3ZP1zigaQDsa38osnlCy3jig
2PY4wqbckJXr+ipuvjiAoDqWeMOO4GUZFLTevIJMgPpD4WUTomxtkM2FeetEbPnoTk1asUxr2j7f
aAWxN7tLMnizes4M+5GYRqIqWE4s3nX5L/m8M7oGhJcxCRfRAy8WB2jxNMNV+t0z6MsNaEpGwQC/
W9eUJJaO0yES61uksw0e/moiqPU2pLDU0t+E4U/TcKjvYuHAj08133Jhxpvd7nMVaMuUk6ysG/Vw
RRnfDPnoODhPh8EEwPvBpQzAHuV6h9ObEfF5bMlRRODr4/ln1VfGCdhzDFM8DGnuycYM0veFsvYz
v95gFo4iAWItMPucicIkIoh2xmU4EObEv3j8q3fmF25z8fLRwWGUnVSr6KXA8yj8OlVX37W9YtkM
zQ3l16Zm0J1PvhsJDbmeKwSnsviorQxYISZ+VTvnLLhWwh+5MyVuKi97AjlDKnDMMXk3OKNfT+g7
TU9ggJd2MDAYMnscqE0uT1iTJ+DrzWaqOUUzi8zBMNukNY7T/7Y30L7E/7Q+ePT85qo1qv9b8zvz
BE6FbHQiRwKKHnnpJFx04HBXbMHs2Q0R2i91M3VRBwXy09zFeeXN2q+dKdFuD7NPpN0PwkBZ25Ww
8TnWPFUBO//IcPn77miRC4TbqrGkKDlohw7O6J4M1adM5m16ZooPFUg9uw4AQ5cBlRHvRce5rS0F
VgVQ5kkPkYrG7T4dchdFtLtMJQ37fKckvXlRzuBknCKlPLxz46Tm840JRckRs9lwewTQKmAlE+8C
PS85IGY+bErr1Dr6uqLGhgBD+M4AUmLfyML9+HtpQ9vWchtcNVjp4SHEue9ZuMOMKnf7r7b5ZMos
crN5L+mcFr9yv6d+Kz2DbvU9l+rwISA+DMIsRpzXw01LY09pj67qqd6hNSYRRSLACft/nk9fuGOO
7pAHVf6lhG8o48sCPTd4F5vG3ylk1dRS7CruQYpiVdkMjrzet8C5SDkusGgVuiR5tpROWgufgh8g
Zp/eRf+oKhkNpX4hYfsHYmDdJFbLpQJRLuyF07trr2jbJK8cZqMxwXj3fFJTHLFi1Wa4yCEYT2C2
R7nlfkU6KdmiTCmjzPBTi8i9QTYhrnkNvRgOfwCzNID3u+eBMxlzOjjgqfKCwhWsMIZIaW3/tre4
EJj6sWxQXV1lKh59ry2IasSre9pQhsigLKGbcKFwg7MRlqpP3dRWFUocWByyppK7lAPJwdtriX8Z
YJ/8RFx3putT0pO+B16/kkngLUVrbniSOa+w4kYhMSZsPGCoo6Q09cfWg5aTXuHH9SjcM7yZzr3r
L4B4RiaHRp/EiRhbAeePfeCBtcPFLWSMylrHr73hgA/9yPXj+s6Gx602cuhGtDYloOvtyG6PyQo6
0A0H3PjLJ0W8qxaqAqOL0McnH1Pvmvk467rIlET62NJQKWspT+3NwVfcxxh/Okl3mK8bgRXapuIo
D6tBRzzKKnAlsDvAdRtkJHSQmi2tnDzk4lE4NzvdmtNTK0nldJgLYv5UMKKnC8UB6SoxBWbqjHcd
xtK7W/5a373nPOKtp2j2BaZy+cfAQVXY0xBCGuBPA/IyaUBUZssA7qtvGRrfAFNXMDOYW2v9MsNB
JN3TNjaa3JqtYhlWhpdJf4AQwds1SDIpV3PpP+4/IkYVeSY9DFmtSXj7h6CFZvSTvrm6mnfb6LDl
cM5tKcLF6Ed8+CzAPGTzDC8b5kyefI1s+7mRHMHPkYvFiWlV6qQrME2FqHikIQuaU3MlXpQ95JS8
R2LlvMuprgtOpxGncOr1vhKuD81BG4/0vxojC6cle4+L7lFIU0tPjuPAMa+xb5/BLZLfva7+d43C
iv3DbTHovBMFOid2eWf8JHG4r0dxJcJ5uZYpsmTn0TG3wJT4lV9IvSzwI67fA+jkZ6lMsoMUWTRV
elKuxCvR6qeRkwHQOPu+EgzP0xe5L28t8qo1I+vNxKIO8x0TsBtuGRBeRk7w1BhJfbP7qsHMvnaZ
3/vrQeehoppP4J2KFM8fxzk1A/7w0WF2mehaiQyP63gQR1yrRDauFFDDqNEFOM3ankF2lkanPh3T
v/LXQjr5ro6UBjlBsHi+Z73cwwk4fUYZ0IJX5rMirQB29tNocrsS1fMatZw85z5ohyWYqEaVmGEU
CmN534W9/ANfGk+1OwrVEv/Gij/12XeOnDVTMHcrlJ6aO0YSv9XgzFmQdoVAjc3Pb54ribhsPFiQ
msY+HwSqlIvehGL2iMwnyZ+SdnCT2vira3sYgx7IDyRHWLwCLna4H0GKxijMPIaMBV5pZgsxLUFL
23o5jMWcC8vwH8v88bksgdITc3bTkPn3Z8soEmKi+KShBZeyrmu+ou+pDVY1TkuPaxY+0Gy4czLo
pbGNoDMIwyMFUtiDKsL3gNTbW93zitpkoNBmRLN10mxdLzQvfldgBx4vWi1hjTUsEpY+Yk2stRdy
3caaBoKzZHBii6EFFT9OmK5++HDbkJ9v5AShnteP7dqIzGXAezmLd9gUOGboWd/KRPVMMYIsKtRX
ZacH1R8Nm48+05to031e9/J6jlw87/YtM7L93Tj2d+7YZvIZrmZEtDpX0f3drsQV8EB7qKD1HjLP
fE/VKCsILMbY2mlG0HZ3uJsn01+lvOtHfoq575CPhIUcFS6kOvW0rcKmXv4jsUbKD0DIeb3ZnJ6a
m4ejlQT8u5BZrDfs7hlohMs5tqSmmQsByIHDvDvFfki68ul0ltUsBHI4aBhGeSJE1Ckz8Xku0/WK
S4FAjN32BIJRwqdJ5g561BqYdHLmhjEBQ3odh5uiy/W9A4npR2286pBYppfzlxIFX1YOZZiMn92d
jNDRi1Q+sY9YTWzwY+XInccUt1hGfFxrWActh6bnz4rj69WcM4dxv3+wmkZW7bmkuDQBFh8cD1K5
kMGoG3cyeRbx0GL9y6VKFaL6xTgMN1qMDrIgMqwh9JJtZXY6lJlD9gALYciqYnGrD21+xbh1ZgeC
WR5LfMkKuar8neH02lBaZpUc1tw7AQDfY1PE+mOBVPOIeVYK3iWeUcCepGA1KBR0kHSZVzRVu4OG
LCCi3dOc/R0hmU0IUwWE4wOAHTwbUPrYyu19Mbv5lbdh8kFcpBHlGvO74C3RLQXiSwhlxewcoSZt
9WW0Uwm+jVOu2pyqbKvYNxNn0MF+nKkFoZt78UBA+XNvV8W3tc0Azsd2vuCtD8YNF+mdRCUr6gS+
18rLGnpC7K62nEkHpsIpj51d85E5DJydgwulppDHQbjSpSLnCSOjbox1Z4/AvXtSTBssEFAtJTsm
cCK/2+MkBmYvcOO4L9PA+9wuCWj5XsozWd78ycegnMpv2ZbmJIM8v/lkCLtKKjkqiFt5NwPhhzyg
dLaULIEQULDEGB2SsqLkeoo9IgZRMpgJIXuoEkVkzgszq3yaPVCSTO1+tBukXraEdOJ14a22r1qY
1HItQ2X+guEWBLDPh8IKqQo+6g+hy+elU3hNQuKKX8gc4SeEV9t0/0shOipsuaduG0/MvHkmm0b5
M42QbUywipHemURwdKDl+zWfKhzOXtPZaVFOApjO+fzEbHPb00IASfSI+IGj1hFgwjLHzZmu7HiI
6+nN2HXQMZeTp8cykn3g+ZQEOq1Mzn7CxZGkydkZwZYEfYsvh63u2b+RDtXKWMGsVJBk7ThSS5Hu
g0NQiLhrUvxQXfMPaa9ylfQqKtkk7EyNaQaxI+kNRbi5Es/Zq/D8931Jyc9mO40rekyjKIVRVaUl
xcGl8gcQAtHqJSsRkqu6LJAWAjF6t0F0l4KT5YlDFN3Ksbgp+d+918OPE/cTAkW+B7t7XzHkq2cw
qxon0xAwvtmZEyhITMUzU7WaUMCJa6MxTv1w2rnToHLrSmzLz21TlLnSk/d7izS2uKywPGAR8GNO
iZtoB2IkFcNVk8AKlIgfGpqrU6gezPzBJEBEhbX/c+w4Fln0CP/o6spaAgQoLEsYaolUGvVFgfx3
hWGF5/MkYUDBskc3DW9BetEnOuiLbVnygwVqfFsSoCXg1YnImZbyRwEwk3GkHH0N2O4U1YdkgYVw
d5ykJgEq7skCRh7AnksQfvbtgvNZ+FxRN6kAEtCOfefoRa4hiJ1G35fuIFF+opg5JiJ/+5WkadqL
+XnYLQvU415lxZ0sn1w1kX5kRy5AqtuJ5sPuDiSRU2nJ9kBYeoOeHThQSgpmUuFkWQX2GxiYz/az
OxPGmaYph2dheMKt0Lf2qBrgK45XxuW0HzNufoJItejksDxSAY3nMGSdTA1zIkFVG+Ks2BvbrYSO
VWMXtrluRMT9H7FuHv9L5xgdUy9k+ei+uFXdeLyzrZpJ1aGmJAPt48nK6nfg9l4Luu5cPYyJ2x5u
V+XXYvk7v2EecvldezqaTuWgNy1ECmxVqMI4e1GOZMcd2A/RMqVvRkFYg5thTju9uOqt5fOPV7oS
vOULJqMNAzALexE3kmWpsVL+qL8ylTStds45OJa72ejsaEIW5AZFYouqdZT/I8zO47VFHg9YYZte
T9wsG/hYglbBP08S5/DhadK0hlG3jAgvYqCVXavMzp04i6wD+Evqb14kWRHUhFHmytQcjJ3ZR1zJ
NSFY9gRqrVZuZNzR6jS4pEoabwQz18NAaWxvtIs+Ci6FqmQWLzicdjUu2RY7RgfyjV+JdjVhHaJe
GIcohLQ4Ef015ofMDsCT8QTGBQ2wLh+rVfvGTeUQjkQ2yLKvlxht7sM+u9v8d4qM8NIv+bO1th7s
khoi0q45EuJKFh/ijP4rIwTC4CbrHll7oRoP+8UpKen+dco/K+v8TZRgoTAI9u1Wqu28aQeODpaB
tFS54DUz2PcB5uHm+qcqSCERu4dIihwrx2xjZE73lRFPhGtaTEcGdDtA+y15svyw3fx0axDtC1m3
IGowIcfkUtygTnN7BUWqFy4kq0DhGN4jaeh7wO5OsdFqgXIceRP0WPCFZ1+Xpm93rQeK+d3yD3MB
0m0a1EHi67oWxX8plCO1TMyHOBsikODtloOe6bKKbJTPVUdfvrni/HOVS7qvA0Mj6Vb+4XikfhFg
KDJB7WIZqY4f9SvDmCxRrDaOQhAUSea3v0iDRqn52gB4c67kQ0v3L7nTybmMRgh4dgWQj6JGTszQ
Lz6KmCjd4Jx7adiUrQOnTL+1JKRTs3nf/LomNjvUoyTfYHkOHQpYsNyNTeWyOL7VhJ+1hxJWnEgi
SH1LLIi6wJ9Fe2YrP6XaEGYdCghCG8B76V1lGN1iEDmj++negMh/oMyymeTkpeDBfhpjyMKif8H8
nR9dCfs9xlhueqniq/CeDiszw4HgfiVSNfGO8+jNjpbJ9pb/SkvEA84PRqBqrKnm9By9SPB8O1x9
hrekDwWF0xK8JBVocYbgkYTa4SBVGKbwCXfL4XkwwVHdq/WHcXm4FUmfpPg6LufYPT+BaiqsJqir
K4plNuIppOdtWOw7NAwtfh+FJ6s0scrcoe1ggmo5MqzGlaGzZeaYxHS8AJ32ok0ObF59Swn5wI1g
sub5Wu3NAa12NGxjZVLvtOx0IuVrpzQiRBKMSp8SVeGkjx4tFFT8mgcR2OWc3BOiSV7opkzmENA/
BXmNG0v8WbN+j9y+Vr1OLjRm4ZHYRH5Ro/XHaNEqYuf+VJXBSciRKH44jQiFWS75zXjHYwp1xHtZ
qCZhBaamkqetalZhikMcNxXGRjxZkgwoiqwkrXSpPBPX/S1ShMMSuLjpzqgpI+6jBUd75wMwIhBI
dMr2zvfluBxFZbwqZKnrLjbWDl16+YVgZoX2tYPS33yl5qcwA/i0rAZKSyLx3EI65iPz7WSjwOE/
V2hViSCCLZXEnlDmcJgO9F/hALeAiXEs7IlMVfM3DaYfL3yPTQe6E2972EoPwZe2cZNNkDWwAITV
8/4tyTWR449GzeizT/DxkvuQYFypOXXvYp0s9CgtWx/2couI8QbiEH2gyvzgQJErshPFl6NQUJNj
sPTulZw8TCOIfQWIc20GYm/r/+B5kjtPb3ZxeO56ecPEHZlqB1x+oFdAJIaeBya1sjvO7G14+hgJ
egS3TgvB5WZvNqPW2p/iRVpDlfSatuWwK9t41UUA0uiN5d9ZFCYKgn/Ejsjol0If7K1OUpMcdaB1
A0eqsN1YtJwGj5inI/2MnicUxNDplIwl/pywQSUPJrcG4XLK3zZDXQyt+Ymdi8Slw46WSDEHdsYB
xVkruMyugn+BJfHOCnDCOQrGrQQihK94fQbFPuBsCmPl4SdyglOq0mHrRTq4EFelnbK/3R6ly/+a
WU3mu5aJ7CtpLxKvMvevtd+cStzt6jCv4WX/Iu3Oux+5/HNuV0PPsQszBUz+qD2z82HdUkts98JK
nt4Oz93/dXCZ1Ve5fO2Y/USBKhU2b144ho2lh61XffGqTXv1DzYEcj75zVaKfZ4QdLeWBsR0eW9M
cclOfHqJeUCRGSwrGaiuYbvHF0CZRCmOUPk3qy5PVAtDspO4LhaZuCM1O30PablSewfjwfjacnD5
KIztRnNajWAWGv3oE9BTEymq5Xaj7dbfCrxpwTyqOF1BNy5N1K1dVVNB1F23MbrDwlMXI9G+tB3U
YBoOey/IIOCCR06bhaJA6yUmdxwz5DSgIxzOVD+7f9qQvAFJgW/bm9v2HlSSsegzA9FbgD0edEbG
9CcDtSRRlJH7SQKVyLsQWf4JRULzSyBGvGoJjrQDdovYrc/OezTwcHqoFw8wYxVtx41cAY+KxTgq
+h8TkI/z9vtRGIYArk/RKUuz/NIoIZqug54VFwKkz4SvvW3ia9/TzLiltkWPgbX/NGT09zzE/ZwS
/oHM598/mS8z2RWJCFRZqjFSZInre7y4fdOkZImywhERYIy9DB6BPTqnig94SJpZq7Ydvfvq3ScK
+9ADiNJ2pCpKmhk5B5ElsBj8pyGgdxBm35XujonJ1WA41NNkFX0T3n4nsYkIPSgq68aPMtwxxMwE
C1cywN2v3hclJgF0DuMiefJJRIDndd4Jui+oNOV/JPMqHbA4qXjqHfw4ferKvsTa+ZJDwDHgkhGg
cFR///7rn9eFWBjTbY4mSNhGzy3szXRhzA5bEAjh3xSeTI44zgsTU99X4G8FtbvtOvJVtJwRH1Rb
CVKP4jAjVyRIP6cTxNr1XkJgr0QR/5CnBr7sYc15kAqF4gHegY/7ncGiqMvvjNpazmi55mNt7H6v
Sq8xB885Xq5dj9+OCZ8okB+zFm8oz64odSW/9XVmsXXjI1cw1K00f5JO7oIZHHo7uTX4E1pUtWZH
XeQ53gOkwhKJDB2IWh2MQgDu4baK/YUVJKkIsfKhbI1K30wojSNJS7WE8XjKfRgv742+isAOm6Fk
IcrZqEdoxSpryh76mICU0wIRGFa2Le8BQPVsNdCPm2Jd9SJvNV7LrRg9d3TaI8rnFxtxce5+Puoj
BSl6hG5VjRjNWRIDzfdHAlfois66PHjODm4YS7sQeeE3iEHc60yfMmTGbIAa5e0YKRQB/8KPU+kq
2N8/1jhtyTlKbhKj0Jl8WWQ81+K9fmZ7E+d1Ag0HcUdp2XbRI0xsQY/QLLCaRLf+sqftU9ADqPFI
FdvAsTSPzIhqc4h5sdK/IbHPdgQuDDng/O1JA5dadt0hZIL6Pw42kaUvQhWHk63eeNUyB8dpaPPm
0VYmQKToXnecn1q0JxnPrn3gQC69up+5ummWRTS6tphctuPF3Q4fxo/eVsJGhAVKbrwwo3+jhiG0
ifHnxaUKIIUROh1ofsRU4a2J/tyDIL9VGs9ZZE5UxODRflsJdlhN0ziGQ+NWstK0LVznQlJBq6Dv
KwVIkc/psVtX2Nnqj+1UWwVtdr3b7kI5OVJQ+YhY890d6QJYsTKLzHx7xc5DDGExy4V3KrszwR7R
j0Pv0W/mNv4G9SvRzHqtt5LhrNV9NJv4jYw4eA4eKnn6otdtiJ8FolEp57stx8ai+ex0KVgYoFUM
0V6MYxCFNSWr82lGMOHb3h4StSwC25kKVhP399/EzId707duKopSp47di0vI7EsKsi/PevwZuXnK
7SAhV3jqFOwl6KdtR9aQKb3d8UxAbeGeofZJJ4Z2uVA9qR+lmHqDZ+yzMQyuvU9F8GWi4Fq4z2Vu
mT9czDIAB1qbXDvvpvkYLVTBeik/owD3mYSRaSEncTawRebzEuHgLbAEpH1jb+sE9SIolTCKDUzl
e2voUdmJZZw7Wz7r/EZ05ChLdljvnBz5Z7RwD2hPebHcDztdCxiUdh8HqTO/2wecfrS9j1Yej0Po
2PyFYkXnAChwmivr5aVdEFaQY2KAe8n3pjgbWCFlwvrRuDZ8uAFipuyLe7mOqKSfOm09wJgk5YPE
HjV86ZwnascrwcEnaGEEaj/4KV3v+x8Ss9CV9VWVtQ4jzzsng38YB/2YPDUOD+kwrSk0gVJTibcp
5rvGg0tvcS/d7zp3vjI0Bqnd8eaAgLqueK7m6hfkkEM1cQrSiqohZ7vYhKfINqHif9M9YqNtj4ia
wWLTQ2vL5Q2IKiymL8I9IYXr+EEfBmORxiCQhTEgD7ta08vHJnSiB51umtM+rPtXSOqlsQzz0ots
kAgM3kVC1YAAS5YCpyRWGdNd4LhVjzYOX2q4VEsAsBF5rkphUOB/BSC6BT88Hcv+nvQGoQBDqxOh
DATt4+MLx+QQxOb7p7qVgS5T+OqmcChF1FgHBoQZbrXDMFEKLw6UgN6vsl/ACmy8fnO0JFOIu7fj
dSS4xGCVUAdREzAHGRMkdErXVKIBTg0ZW3KJ9M87O3Suw3r1beV3N1rma0ko2PLCkjhvgDszT+4S
aFGra73+yUnSlThrOSMdm4JWa/snJuCcg4Td3WS+dEz34weP2USMAhHS1jN4LCIf7tHkbBtsBxdO
7pZZ6dUnpV2LTEQpHSZEeoPNooTd7NHhPhkNrk8caT2ja/GbASl2lDWbkx4lqdJJE4ncfr1b3bJx
p/mjdawkogxpdu3f/d+4fFqg88hB/cspOsvB3y1+Dr1bNmfw5EfbiRUzciU7HfWMq4L9qj9r0WmC
ntFqEWM1Wp8zXRovJ50ho6AyF4SeCjNg5s/iOGljQZaiszx5YS87ABN9i7K1v+dobo/6g92Zuxcu
an96gq4HMkC39P7GIujckCZ1ttyh1H1PCAOZpNee5HwcCtVbnBvxeF5yKuB3YgD5wP8cjEcIJtAX
xpPrzNKERgox/fM5sSp0ReW7hIQoXuvd0nV+wTS/lQeBM2atf25FKmiIBpEDPffTRsnq2DE/2JU1
1spIU9R5CMHwgQrTVq2V0faUoVko73Zu9DSawGyG9N+yIHk1bDLMXa4HIgNpxcroJ12qJWh/f23l
uKdpcgNDGM3A7xVe3kWIqTrN9FWQvQuNzRLK0JfPRDnlV+RnQabuTCcfrwRWEFwsakGYmjfoJzSN
yKBLLwkvK3arvDkcl8SFEtugY7TBgZFMpxJTNRVXTc9tQ09pJdVy9ibGIfSu+VrbqD7fFw1ZeMZ/
fKdufy+ZrFSkXDi7AAFlpRMC8x5b2t2+maaP+jzqNM0wo4+0WGH0opEZVkxqNNRcSSCwzvBmy82K
UfA1oQqGn96bbvL+HLjh1bRjxTD+j4+mBYr1s/Z46vzg5FdD9SUQS9D/0vHas9RdQSZluDJrD7LO
RfQSF5OFjSmCkzrpxMtCXXNUWBbrZiF8qr0LAeCXIvkAbVaDFcOGFkicnNgkBVp+qfsEe+2rh8PL
rxx67ybF/n9Az0qm7LdIOfURoBSpgDbk5YaetSVs9jxdstm7d83exd55VnPjD5g+oewEXZ8Cp5iZ
I+Ve8tdKtTGHIaZbODMJx1pwnoO9mA4sJ5YHzm413QWiU0oENNLtdPKhyirsOj9+yFvn69wZuZY7
kVa2wuCBW3xRJpTg2FszhkaWPG5SJ3GKPqkeqhqnPOS3//2azW6kpfROKkyWfjqBsGTnCoE8jsvw
AZZAi3v1rYLyyqgzWaSfqu1q9QfjIIJ9u9ZgfJtSnwMsWwdJYEm3QxwVqItDTCE+f+XZLNo38JYN
3wC+XmqJ4cpwM6ZjJGfqrupvLO8UE8sfyNLDP6nXLyjybBMSemefRAKoa/h3SywioqQOY8UxuBCa
3y406JzGdQe5DcqREw9U3z07OjuEi4s6SJBLyWubh5+fUQ3633AdYjNRJ91cy98NlzQDzvgt9mhQ
RGet7jtw5yfJdA6jCcQns72ZgfUoAwb3fAD0baGJaS3l6Z/oh72JsAxlGzllHIeHyfMdOgvuuKpG
/lvDUdYv18CNsI4W/1Qc5QqIjjkBbYlpxiP6ArlnFm+0aNmc1YUBbBGk65AJOCyqassGRhEfrvie
h3rwq8rK0Xkeg2lManwtidAc7PcxcJtyP2hoKYW9ENqZIUBFpzmaAqYUNOKUlxPuk2kB3p07nxGt
KIg2/2siF10hU/RrMJb/laNr4PnJm79YVOd6/Ax/DWfkezbFiRgUgL+RGUcK34ZUHkz0evusQgzf
8EnP1kLhURHoDOsETyd4f/Xy4MnZEfsw/AqopwRKMnlsSavM7jsu1DiyEnMVk5uvrT2FY9Yx7PCs
kXDdLpi555eNeY/Fcvz8W2hh2IEeyfK+LEWLlfpg2Kh8tTQpQKMGKGFrtWdkOJLEwNWL11TXueVJ
0RVDaH4D6GAgqp413SLfDalA6HuAHrxwolGey7nR2iZN8HqVQ7f3Uv7NGQfmX1Pc+Eb5aaXUMHxo
e4GH3GRL+gQHjGpBjSSiR9pA0RGHINMU+WvnKLGWsN1UvHH/FQZfodXaNgN6S8qBrhMp1BWJ87MU
OfcHBy7IPQJTKHzdAmEwhPcFn0aVCWWznyiygtlevElX28T/CuiAYVlD4EUySlCoD3t0QgG7WnNe
TdLy7+iVy7C3mkfbV2a+TpMtn06LFxda2eVINw1gBCzLQhrTazApRI2q33rPcExjQ5QANNm0p8vE
JbNI1NlfHWumCI/5MRN3D4M+kj/jXTm3JOsKd37Clr/+wc9dqALRv4mbAqUzlgikraJlZphrt4Vu
7SldZtYUJ8i+NjM8lDywl2+jBas460Ui6rYr5GIAQ4O8+5gTqguFtViadDfCBrZ2rMp5ngKO4km9
PFUjDTR2GMIVotgmVEqGR3o6gHBkZ3GIJLCqbFAkMujFSrKZXg+1eXoL+nYd0WP7enIaZYDN/GvM
CaqAaRxPeC45A19Szi0eBCuZSl0fBXeTlGTL9x+lcN0fJvuHXv3wgpRwxGpTA31+uZc3xiIxtEOO
OOZBtut4Y9Xy02mjeJ406sQP3O0Ln/GClMpEmc1Ex68SkFzqlYk5ZrcLo5OP9+vsD/fiQB6NaFom
Y+R1ZWrHu1ys8RGXCwDk6ufr9dgIqFLMRb6cZSu6HOo+GGdpnIaciDGMZluRCa8cliwYrHWQfNgW
/6VwSte1hgZqz/U4rqhCF1BZuOUaC7zhKrYcJBHU7RRc/vuLOCU7kyQoKXFXnRYYVHF9cyCeKZ1j
/y0en6TK190G+tQBgF8UY0a6eOrs83zPKOeXt/gPLXSXrdsr5qBSW8KRm1aBKlTROS9P+ndqFn20
0nvri/+eNilwW8Q616SdMjiJl8dGLCeQL2tP682eRvoYglVAL7+iPZUdI+eyylgUIlhjzuH/Gwby
8iABS2xNPixmHv0Sr/CoTXQJzgdEhi1ORpaMj823fF57MT1mZQbd9UT3SmAwtY/XTVQK3U2s0iOO
tkxwtjOPocBuwyzBKFSy8VTz7PTzuI08ZHKHpBM/wHpkxj8OblJ4V38gVSDzY3ijtptjkrn/RS46
V4/NoknzoO4n4RT6zPnICcA+C7nWsyhwJlA5HlIkV7sm/mu9QyXg0yQ6WaWLQq5WaTR5GYNdw2wC
T4QgF4lJSAnQjJoZMDUWM5pRURh2vjT8KPIXYKJx5OSZ9CtgMvaLpBbWlhtf266qQydv0IiOxg64
7tk/imrMwImaoUuD+xlHzdIhyYMPNxFGhCopNL5qgHll20CLrR5TWWAQheKHnQr1n08X0XvGJVW6
uLez8qjbFMnH9XXkFuYYmbjOBPrYhnRUFv4pbb21iMYi33ydO8kOIf3FdB6IVIYu6fqOg6eRb4g9
N34kvAgDXNLonU92mTiZHJhiOdHrC/FsTJ0QUtoQUYdwofU5oq/oe/i2+1Ls+lSwQoYBieHYcX5d
3rCqLIi5DJbbSVw6d0p6b+hUZa643620i8SRIR+sOnOdouT9bWd8A6hi6lQDcrGRu4tPf3DXQL9D
dq4PppJeJkTbc2qcPUddmEktO6G+rwctTNO5W82hFLa2VZ2DuUYeJona8z7WKIAWZSp7w9V2gimm
m7mNC6fXw02NYMm1duIhOPREmulLoPpFKD+lrxGJ1r/w0XGYZM8oIxPed+Al2oRFuZTjS2JWq8lA
SrCc7778op886T47rzYMT2sHGiOAZ7Xcj3DEUCzAO3RVJ/CjdjUpuAUJCJPVYtd+Q+ognpKWrLUB
AOjif/KanJWtS2jnYzmj4gKfam8j4LAnQEOyYxbr+7c7QvYuXWmepD0c/4JSx/FQ5TdGDH9OMnRD
Li59WOuadnI4Q9yRlZl6eRgsK+SvVMjBlYzGcKFdE6R1Rwd3ZB6sBpaOQN6tq0r6Z5kA3kCqQ255
QtnA9+zu/OlwFdiL7nTMezI5OiCh3eJRFPyNo3gsyreRgwUfUGUxdLltACtzXszmBpPRdrl4qbqo
TjVCZ9uTJtvaZ5tjkTushv0jP8iHIYm1DGcSdlT2e9iJF4NWjyGWqqVoj1RrYIibt+Vfyvou4ATj
yyg2idTYkC6eeOnoLalMB5RrHpef1JR9CsgJTkJ50y5DoIwyN9fEFqjHbuuHQMSHXcgBD7ho1IhB
SttHwYAcFV65aDuqhcqIojnykDkTgb5aXIeGbncx/2EU9IweOpsC5NXR3GPpWJO1yC+vyiS8H1CV
VGyyrfBpvolcMFSNoDkCHSdjxebcmwOmYEmStRSMP43vSZEe9Xq3x83FaaQWfr+dP31H6mhPn0LE
7H2UcCPPh2Mnc8hmF37TRDH1mdihJdunKEV97hIPO32FM5TMqPV/BO9nttFpEujJzmjsF2NOvYvl
9zHkNCvUQD1TVS9vIXt6qv9LDuXsrEmU+Z0tlyxkm0Wbeb+JEEnY3+NlGvpTsP8PY60F/ayS2j2T
mmf+oeiu6x1MQNHvkcw3EXEoC6IaXOTnCGZgikQNipLgwZg//4fMtCeEmutVeKrc79VRh4vNZspn
ng61/FH71X2QwlnZ8v8g1oc09/KRFa5knY35N6l/gt4F+cgtUP26Fb8tjp51DxN3Sff3pStw+lKz
lIkFcEWxNaXcFO4fSFbbXzmKoGKM1UKUzLEQMGgZE8hiXKMx9VPE7VwXlvGVpcg7/T9aRJxahHzF
3GHgnj+XnVEunhE7dQzRBRbX9Nw/37jmhEeNx9iBjmj0kRaucXQkFuERyBv7OsC4qjk9R6MUZ0UF
G271TwHWxwNy7xDl2LSTMAusio010NZGaq5amTyh84oTpQ9wp/LIxU4bLH0rforzjUB2olH0yuDq
nS2Y52nmjDVdlt0dpOF51K04hYDeewnpJrSfdF9t1LRzCPdQ9DLHHOj4jO/TRZe78+jhhCcCavi9
DNL8EsMDs/4FGxYoyZQsscP1+Te/Y5iasEQUtcjlL6mShje4EGY4aD4+nJvjvLSbIM0swBSVMZUN
IoiGur0qqD5+/VKYJ5btGZ0i19PBHSHC2jeFn/FpSnbC2gMLgyvwDLxN7iq2u047C/mcBaOOq2WA
reoVmpaq0CqooXDdKlG5q6rACcEM+myDyw839k5QNOqFcG2J2u6srjTQzrfmp76nypAzpklDCySP
POtf3D05pg6UncG/HvrZr/uFWzIdZKMoW2jr5LJUkpJ3jta0hiPNsRJoLH1Xhsy/c14V4bUhbGcq
cyaiG3YEZxMI/UmL73/7/W2U8v/ydCYFnTbbFFlhOxZkRFV+lcLYDLv8qcEgjCylbHiiiFWAQ3Me
uapZjvCcwDEcm7aLtL3pBNov+KO66Yqn4uZ/8KCNO1LGigXk8x/psE79uovsRzcQS1RYzCcgUOHX
PCU3zITQAhrT6j1VTGl1/ZY3IYX6XPPn84WAKly5p7H9nbxGi5gPxOUo8TBl/vKWdO26VwTrnJuH
IV2muwrZEJWrYfylSYNK7ceZq6Bj4pij4SEbsJePTaYdQvUVLzCcDQ6ml/N0lGUVI2FCycQnSTgx
ttcJwYi2vz0P9rcD6Bzurk4h3ykmBWSxZbIefjfVI5hYqhHy099yOSaF4BpBsP8FvQkLGlSDUmQG
5BZg419/NxeuGhVto+D2SPOoJ7d+8Pkm5cXXgYiwdqgJsi6FjUhaENHBT5e7ocnU/3qBTMwLLkAS
hWQSLPxbjOXWabbf0Gepx22CaNjNZc85Cg0AI45o1wZqtmpY6o1UnCbL0CJ+9jptxcuDk6DTAfsP
Qy41xHJutwlbUrDVWAhhdf4y0dipsHvm/93tu7TptMz4lOggJ5QcRrtBpq9NR/rb2yyxSuvR+eHi
r552Ukd4MQCu79/4KvoTo5jszQCx0LjOSjqklt1Ds2mwVGh5ofp9GknhHPa4vVD8haAj93lsqnVW
XdwU/iFcWfGeumS67Uwrq2GI4YG/RH1A0daQCApRYY3t8WGXDbUbqdL+3r0MsaCz+Ym0xMl6znpx
8KxLLnpHz885AvGEWKhOfYeNbGD4trfngbvUfA7Et8m+xMmUzxns4EAzMwc9Yb05OrpJN4M89bDz
iwm9jlyXrNs2iX0bgU4Gn9mfkQp4eggWdiFFXhqyV0Mjvt5uUhChA0RozVhzrjr27ydexxNtkhJk
ro6x0Gl8kDrzB16By1SF+O2s/QMfh6v8wOiYz4YdbTovin0+I1Sb2favi29AuD2CAlGxuKYcaJxD
3u8nqUZ2HlL6p0ye/IFm6pF3j/jdQuP7BnuNd2TYsQ+1WG0pjz0vwrBQ1ghEh4eV6bMQ1oimDVKP
yshOXuj2yAjg7yYYmhp+Dqbmhm0E8wtHwk0Gd/uyfQYADt4MNZ2uXbwo7zbDadgUbP6wpEujTnPa
8sqhZ4jbzxxWzBDKtjNSRy3Fl6/48pR0Xq7lKovrYORfmQZP0+ngSnk6Cx3eeWFYAX8wOv2V8Q+m
r98PYtkL3X1hCNRii/du9A7QhrWT340u1R5E295ysV3Utv18MeNcKkj+dHBaVVdhR/qt8+YQM86d
D/HCZN5qZ9RdHUxKaB0tuevyeWmLRcmQv0N2l8ooUxS2bNGCmheCzdG1tRL7LgBsRX9VZusKnVxo
eblr+WPpl1RHu8k2CRIf6+ENnGscyoT8/dVdfycGGEPPwG0uqf7u0Hl/PI+epVoeEp+0WE1gfBxk
wV08eFUsUgLIfu0/F0CMB7LNU/K5jQVUYtl3qkQskDRG+oezY5ISR/sarBuTycw5Jh4k2wkMHQlv
kwtfUNGRF+XTlWgGEkmElAcIp9ULq+dXdNhJ6Y2m1iEIpQ/qcdFInhY4ypJC5C5GxEpfiYLaPsXR
Qa/AULOYHMMQaIfBhvTUUtaJh7QuccqnGLGQnAYBCFQvTkBgnWmZ6SVrCkMUg/pAjYUKZmOZ+2ZF
W/R4BIZhD2kBsVc/6xw+9s1yi/8Lbb3jKfWnxx9m3MHkrHNuZkl6O+b5uX42KL0k6WXrfCTezXDi
XXm5j+6ykLJ/trE3Rqdtj/P7h86QQKGEhJgzd3O/URAMMztuicbCDJcEGUHF0J41LVYxMxFCmtGZ
nEj22JgCO/W8jB+DJcUQO4e/M8+5bhXOmsu7oyZYBejTwwjhkTUq9OzjPfzMROyNl6E9GYiJxscH
/tFWm72qBQ4m64IbuWbVNK4fvZZZb42YixfUGETjiwPc7BgD3mty6H/iHT7HNkVjIbKF5OOU+JpG
JqBRhCJy5zjKYMwPJBxuC/rCx9lQmwK0qCtXisn00GueE9qDTpAnXzWUvBv9KO+SYAOre2d6idFQ
xFKAechahn6rOI8TMt18PwzCqAE1OVHHjPNYUwWzAOstH7uRE6ubCOpIPY86Rk2oE3GHV7Z8dR6Z
TsDHqpbgTTInbId6JPHkiF7kcWJXcKCw8px2TcsynfrchU0+FbJxl0hR1hcYXKwB1WAYyQL1ICfL
0YUqx17zGMcRoH7EHi2P/78FZWvsEWpoFK+GIK7cgYlXrh1ADeiphGlqf8P6/QcSsa7lQdi6ZAkq
yLwvkcsm6Oc5HeVfWxu9yY7F6lGN6PtXDyspUiMnBYNmc1M0w85N+AWci/VgyikbTAspTwnV8C+W
TqVQadV2UN9UujGuTTqNQ6xKr+WvOaQwuD8XHKrmS4lT2sVAjBrzz0WbdB4tR47Okkwv+7JJdLVv
vPY5VMBCULws9+WK8qQOSqGCzNzUwpwT7ANz0m0Dd6tPxj6j4fYv5Pul1nTh+PiQT+l8LREP7th3
d7btvu6ofnhUS+t2vLQZ9ZXwLZJ599yAxO1PdVqpUYsE9LzHLn4FJSoW0ROFYUnjFmVXgrc7l++E
xwNk97/uFGF4LdxJxl26fSKLh01ZfVkmScWdqoKARdZ6y61tHoO1llF59aujaqznnI2Sh3z/DgN1
HJW6fy28jGaDXDNYhGjH8S8680SAO3oKXnVtSOe7VKbWvCy2RdG7vxojIJAkjjMTUWor3ZzKcuWN
8c7a2bKT0248gbtsUodeIpi5e2oXBT6QH2l197C4IHyUbARTvgrX0Of5JDBwpvB2u2fIc01FsL/K
ZTmZ8u4rs5XyDHJkFveUAl7bP0OxHX7+Y5Mt2BGCA6h1uGZ4MnK1myf3coNAA6yffhHYMaZWPPPP
+HOkLA+xpIkEtvoEQGtGg6VsQMuXwPx/VyTdD+urGzCjD9NK3BmyByRg+Bm6JfwXPGF0dWWZCTiA
J2w8JW/E6jb2o/Pdr5yj4N7WaQ7QQyT10Ho4NUAzAFNiL5OrU91hs+T9tI9WbEtQbukYGnZhHku9
B9hjhegk6hUIOyJCT26E3wnep3r1M/AkfV1e0MZdSz/1JmxCmR7U6UO8zGK0fb+6CXkC+ivavLAa
mmo4UWl/Ns/N1DGqSLF1jFDaKCUNryAxVLRTit7I2NBZsiFWZOOcONt2C9d5GDWJ5Vej4r1o6V/M
DpAEalV1qsCRcCwwd8UpHmfZdYxYhPMa3K+E5xDpDz9fD/J9gRbeVr5aBOvn/xMg3lBP4Ihnwr6v
6WSDjmpp67kSHv6+4tfhUM12ZwHjOimY2cGozJd0FcZHKoOMNFBAg/GXSYgtcf+kSLm/KrgOu0PU
ROGRSv3Q99YiEZphGSHo+gmJAt4JbaS1hsHxyvDMK+XJEt/0S6Roz5YwNkcknHLHxPAjCkqGmnL1
AB4z4D7BXtW8XFHGHunu0IWQ6j3jmVCyEdPYyKIs4IprP9nJW7aG5aoDFveakfidzymwDPBDt3DS
/m5ch1R/2TGUGHjvt3nTyuIJ9yjlKvUemFvxuXx7mVrb21XChXs9qoKEVJs5J4MsBVARRQx/8VtY
3lYtFNQAKlkpLrIxVRtQUOw/Ud1gI6sfj/s2RzlKYYtXXo/kWXp1KoQignm21CnY0EAzEjmwN9jh
gesk13kS+KjSFV94QeZYa+X7nYRj3UNstZLFNKs8+MW9TFP9c8wjRdVoE0V1sN4vkEDtyYZy1Kys
YdxaCkcDWu17DWlZjYLzjq7L+X0JIF2oJn1ggYXRkMKWUBfAfE/7wuux8i6A+V3BBf6jf3/wYd1N
vmQ8lYtuTuQeaiGY9sWUov2FGN7xpHYgR4GgmAfvqoExljzKd4XXeHSSnzOfjOyRJncV+tsa1sPp
9DKw/+0GM/QaWQXM5KZ+jNku3DVryJIAE1jQbALbn9S9RuryQSjNSbwRpeIVid356GMGlUqAEhXS
LXils2oUKQItltM98FSTaPlTUQhDdveeYNnYHkPkUPjrc0afZJvFq61GCdNZjFZKH+iXocEuMrFi
EE4QOS5CTvzWzm2dBAuKfV07VWbBjmZQN3i/TzooxNktns7g/0sIcx7R/kigVWcnsBHdCZm78WJi
qavKTvIJ05sCLHwKzsh9eQcoYWjQ03vUZAqeU+DxaIHfPCLwbblNiN0sS00kngUDEq4ZDwsXOUVG
P7LqsnbLK4BlOnJYVMDL8M+mw64ad79cbRlHQs/bBTal8/dY1RS0g+1JFCWWdFF2Gmsz9B+AKquu
FU8GfU4QptoO/J9rB0uiucj/vuOx0qfaNyBr3EPDSDXbrJS5DhQTVdSgGRDPHYZii/MfAIGVbQpG
H0cxvfJhqHdmA5ZF+ai1a6P92weqbicvYXs+ibqd/AM1WyTY64d9W503Xn5J2TY++89vyMAEineb
EQpBoEx7zN+RyYYvTPBGiSsfgf2n1fZWYoHXL6oRApXGPhmewEwm+uoXowQ1t4uk98eYUV+ncqkc
DKNFYPW6mfHtQRQh4OuzVkTRppVbkPy6CM95i93243u1EV0Oq0AGw86o95e5DgJRu2Jgu3Y6PmPq
RXJEC9KruGUCgN7oSByxyezLLbqmV62Blr/Y0Fn+BJVuQovooC7W5DgXD6t3a+FQUU2wuI0ENhjs
OLHRkldwmfjwo+MzpaWc4TGchsjXPOVQnsKHmh1kdnmW25F0fmOIUOhWcUlJv2L6zuz8f6vKNJ3D
QSUgyy2aSFdlT4EuvzNZM7ej3iKiKGbtWmIOy32mILJhacT4910/bwMN0wWTDX2gdwxcbXIdRSRj
Ha4cYJjeKHj+KtVsd1vAExar3fyqM24zEgJRcC4NLUlOKkSzs7vGl5e6V15ZNXSv5hO84kj0Kxbc
8mMPne/QDIqHWU4TT7MHGPxQeQjD0Jw5ad5b7Z6J55ExVIufRQaN+AAHJSRxdRxeiKBSJiaPup7k
dwe+zASadCEJyJFYhEPO8E4mE3KQ07twWmqzkPp4N3HfAb9q+pDUl+9FhqDbHEedlTtAoowsTjzy
UXaGiUqGTiQ87Qy7TMNx6M9uz2nv3wJSMx5KzhTP0r9GichtzL3mtfafVzaIsNjZnjoTQzd6/IU+
tVD3Itnw6iVxgtQ6ENW+zH09Rj4VgW4OpznVRT4XFr7/x4NfoKqsbpwhqC2a/aQLtD5mr7Nn2EP5
Tz5SGkj9hN8JYQGwJgsv4TC5l/X45nTs6BCAmpFUvLuECMphifMn7E1ot6J4EjaK5apv5RQEMKNB
QYkYsSb6lwoV7Epl63ab+EvvBEMjYe7BSkJsmPzqWRY19tktoZVlRC8e85Fr6D7gfarxLQEQehxt
btaqoiDY+MfJAn/eDALdIuQjQ+WNh4Lg+U8SCIHYKoM+pRo5x5dpyfKYSIXN19qSGTBtfjzDx9TS
0fqqMu7CWuAycbw8KfFSolooC3rcHBCra80ANMy8WGyl5RxQkrWHZpcx4dQTBlqvtCP4gHPH/PlP
qeoZppJphfzBWPE0vQFDwhRqY7rVG1oZH46IBnMFTQIU1VVV1rXT1kGDr7vOL3D55ui0eh3XzWEk
KdX6IDJulNwTUSIzvMf6X+d6Z7zdIYDw9ti0lSirFVxDWRKP6mHcDDYrkf1lO9kXcs97p/3/3oaL
Jxlh3MKmm40vrWpbnlDvegTKRi4TsVG3yrUUlGHWZ+y4QyxvhAfSSqphSVdElj84GmKB4VobJ/OU
meJXUccOBVpmCQeZH9PROZeuxmZ550fok/mwEMYqN963HUgNIRzKGBx2BdykSWIbvbvrA/uXxs1T
JJP0C46wIc8g7QuRPYMFgEhTWIxOrXfT0l8Q0GwRn++AYEYTHT1usz8sfznkPiAzDeHg95NGdy6Y
DWU3pVzGpMq06MWD2RHaMSOvkQ7X4dICoRUAWmHn3uov3cEKbkjKiQT3jRDCsXy0Ugj4pqXRpz/v
89o15oq5C5w7+bjb5eRI0zVkZut5JGyrUj8nase1sjIhz60UbA5RCUfOg/YKMq19gnX8IUWNpsaZ
dBfWxP/C3COf3DabrHIoziALtPBsjTdA7rftaMNwjAxWSNXcKtwLPDN2NAaoX6s4hYImbk+RLDmD
3aXzybwjRFbpcZSjIG2gUxwckQ9vSfWSp9vnvO5mc4H0XuPlliRi8/Ec5K8AOte06Y6p6Z+8DVHR
/iE6Xfu72Jt/J3ZR6/JOVnwNnwUI5Q7SANqglEeevFbK2UdSsEqamr0FI7KlxrJR0MHlhbXXblhD
3GXX3DmDaV8C3wCv6qNwoGeXwdwVlBT2fy8lzc/8Coae+BMuaB9JvIvMile7b62oPhv7+VsId7gP
1yzogmiqbswMMs+6KxHL5Rz3XKyIqg4SyeQ3axeWmRil+54ErNeGgSpQWPhUs9RpuUjd+w2QClzt
Qf/3D0UAlk20SGXLsrHCCOyXa7F3OcG0Tp/APcmPda2k0+g0Ezq5Jux2x6+zMPcIMJyD8Ss2mcLj
7D1S289KTPtprj8YdmVnXmWU2A22uTcArMOANbeCLfvqX1goEnu1XuB64YSAYbboxVokBany7DjA
tV/TBJwjzhuETT6mCU+lsOneYnpzvBQLMjzQ+VsDTHOMjeDXjHh9caILfqMeuzcgzSkeM0Q5IrbI
7c+n7RTCJjzyd4uJhMwsZtf1kj/SvhNDdlUKZW2BLrLR1s2dLOge9pJdz1IbeYWf9ap9P20cp+IL
GRBLAOqLzT7BqqX9v6N5wAvPk8towKOp5k+ET4M3Kp2pexrZwjpL/tyNqqih0FXRL3NlB9G9JFS2
gLEDDOD13zZhIfAOb99ptfY35VvOWgzMsal/dDyNqavZQkNJ+BPM5fqjFrcZ1ihtYp01eOjLnMi3
vjJMDJSWOGq67iJ9KXkdHKeirzMXa4FwX9xlWOhjUFnOInGPIQygeFGiVoWhk50hWvvi4ln5mcU9
758W/FTRdtdieo7fVwOo6p337XTt7VTMSaYM01x9gu9dDsHqnjport5rjlYJvOKmjaQ7+Oz+aPrW
SL0l1Y3rFSi+9uyTbfa0TgP67Q7iqq24Rg6YTSa6TxfDGtJG3WE46uqDyzhI2StPagMxA379g+Dc
dy9Vf1X/GI0XplOdb6VuJGqtzlrnY0jGS9q3g33g+wo4HtxyQBNQXk+z+Ol4Ub+BxijOpCxGEvVc
eHWUt8QxCmFuELNqS/gj8CgoStdTL4rwisHMFDh62zisxBZFeE7waXVCcppWiryq2kpY3xvgy/O4
n+QbQSCpFK1XdGXesYfD7FUPTEX7MLpq2NuJVT0LPnrswRRWQijjh2S9kpiknVWE2Eg1MuFSYUT1
oDk6FHqOcITY/ma/CJ8Oz3m9bM/sD86c+Tk4BAs0oc4saVr2IyTedYmqJb4Jl8GZWfZlDQUAe7yh
uhRUAGN+TAJN3sNW4MIoCqaffHmNDobrmKf0CXxsHxOY8eVTv/Vb0e9WbwoaPzVJfdzInlTGSqfG
HM6qAQtgapnywpROV++UPOoGltwYASVt1bU5DW8T0mJ+vZ2exgvWTy6qPk2ho6sv7MOFudy42Y8H
m/zwzQxhP3oxf6EA/TL3o+Z9wvDI/XNw4nkAgV01C2/mGOsWpTehw8Ye/1LSNf9yv7HJzpHuxw0W
ouybnZ1ejLDm8bUH01NjzbntOcBCkNHQJ1s7Ukd6aFtpHMkf5kSVvnhnOwRT0gvg5AexAJL7xq1v
t53rhurPFkW9mVA4Y4f+YdQYzKeFQv099XCHZG/ga9OfuthfQ9Iu68NhrCKqFfeCPjjdH4tvPsSs
T+lpZ5+9j+mJj2tekJQMDBaNoeVBZjHsfQ+qJ5fN/kyaVpSbvTZJ5NP6BUc6F+bJst9kv3wGDcyE
AduUo14vuGkWq6hJby6ggKVJU38J0Dvn3lg//1HL1dvW6F9r2ZsECN0CdOKAvk7rVRGE8TMFIKFP
LSbyEF/9Gm0peRfsAU6wg1p+ktDF0WZnta2fDtZKvKeQUHOxIE7xVcOJpWudllr3EvEvsvEYWLpE
1/CB9lsMHMrYQgcL6I9Tu+zuZun79AGueQ56K0FGbpIkWXnfKkCLdJKtYL5N60W3X2kfhDIMPuj4
7ArNLYnGB5kgq3h9GiA5HMyEs2Qr2fEzwskXD3fuLFdVUQ6qUdTbkTrbQBPyS4tjYzZ+DIqSohD4
LGWx/AOR876rrZ8IovbZvMABnCm7aa+HxkAylIs2TYOWUxsOgilsatFlYaemUAUCKOk32Qdudg9t
dMbKoe+sHTz3BI3ROnvrrDesf82JwQF0tQlvpfu53FvJWmoDFNJxfDsRPzRqM65BHMHF09ixcYyR
32UgLUgWqM/XF4FYotHNalfTwNhQv+DuZoJh+lH1fCPuV35ZmupYvNjESoufpVGXBbZCmq9ZqrMU
iB08EGt0Q70wMqNfeD/4j4uyLp0ikPQ/2Il17fJfgIFdGeQU6ZW98XD7we+s7Mc3c1Glfjfkbbcy
XsdOtAFslLZvf+KmIhj4GWCep+vd7G8kWrU0xHvkpqTh0+Q+D1FqMmtqfi3dPoMMkhBuiIRbH8TI
C/y4+5JIZ4cTEBbklCHCb8ZOiZxalJlXtmupbxDjvscldEKu/0YHQsk6Ody+pFt5ExEy+1iD29je
Xxuckett7V8c+ZshxNfXy/1pTMLfOmu4yrR2FWC8cZ4G0YOT2CYY8DJrqsjNzQC5tuOuL7H2sWOp
nZuMf/InOBGnZkgRCZ3vC0KNh/wD1VPCeRtyvpqcAE/JhLVXOQkpYiF6sm4yQOs6ovFR3ppvn6CC
vZ7Z2rWkVueU8B1EgBuo3gg6oQjis7R7nXwB/w8aqKHept2+j9KWp/JgOu+8bOj339tpBZutvkMK
9FcbahTs0O20sVoYHykC1tJHtaC/+0KOEKgHFfYCEGrVt8aNgPdgF0v3h1u7pCJt86M7G07BRtIq
vQteAsZ9bSiihMjMGW93C7R7mtce/w6e94DHlvo8RQv3looHA0GfmtKsXHCvUfSEtUKchBAFcwbc
RbEenJj1U4xbOE0CJ/7npTZcMJ64XlI84lawUVubv5fZ29y2EHDSxkG2JJ8y6IS+gWVRUy8qeMtT
gHjBc+Nm7mKr/fa/mYbJeOgXt7Y06VjNLtmFxVr81DKoIjaB8X8C5+/kwTn7czNe4N1xNG5WD1Ld
xhzzzp/l55+0HVYpMtFfhjvRcIRjXEZ8o8s5MDKcVdKx9vfWP4aDTq+BEdUmXPykebblyTyaw8VN
UzyEKzAxTJM2D6d7sHoQEgw7uMmKhsEQqSFi2OddrvtjyPtkdWP9FG06FIXVsrCREOBSFC1Uvimz
tktjkRKUSc4ifu9uTF8GXIGeR6QJiMwoO/c1HfGUFpadJkCkHSEqKFy6KVgZ/VjR1tvPeTz5sA4I
VL5Nx9vkB2bxvZxaA5SNJQ7O0qjhQvZMuXnnTGL7P5SPoph81yc6emMrRDM6dKdJQhDAGghTdUvb
qquI4cyyjR1HdfL0UNg4Z/h+fhNdR7i5AQMfs+CeYlbEY77rIIXZg3Gyp9C1iXqLolbwIXKtB25Q
FVZLBswimUynGnvK9x91tGZoeWYz2h6sly4RBNA/5kE3Dx755dHSIJnH2zBWTZQHETdamfdIrdDS
Z0q1Wd8wXxIUKOD/wWYQdRq9UX2n/JeMV0x9gAmAsYfUv3zclBDfGVnpS+XuZ92f0Uhugq059xXO
AgbMJ7a3pJsQulNZ5FA6EvGuj1Xp9tpMKk90+pCQ7biwsPv9C7t0ec8+dORMRDk8FE2aKWxkiDnM
wmT6M/jnSNPiBiHLYqAlKTa4aOvDJADm5b2U9OTG8yn3gZUi1ghgw3m64/YV0m7T500pZxv/3fkp
2n6apew5Kjz47Yhqg2vO73yf+OWshSITGhPcXh19xgHNR9pexAixCnX2aKhtzmZKPHav5zRJlAHT
PDNiBmfB4eL7VJ9Dw4Z4JJ+QPezGlS8Fn2MzY0+LN/x+JzbLENQEFDaANVNa/NeBrhRoZjb9GdmC
Kk3POzMG5vnPEV/ITwg0UDiSQQoFhOQ060Vc5IwNy6FiNXSEO3q62yr3eD/AMskIvBeMPN0v5zWE
dipjv1H9xpfkUveCnZNTAI1jyaawGvGuYc5ggnobRD7U6WBfIPm6FWTr6EuLSsWfA2MLKaEmTRaw
cVTdchv6cgZ/OsYnjO56svGl1eEqq1RYcGN0McJdsruvEc6enr4QJJjQ0wWm91GPGQh2IEVnxMmQ
fKQdzGUyHMJ5ST/5liJ2XqdEFUGuKeDrW4pui8rEY7FKb8MrCBYuaIhBXwAjaK4A5k9K25z91fVA
BX4RgKUPceQ4bwE51AzG694CtfscISDsE54w3WwPaIGt1Md9yOjvkX+Al884aK9xKYxgFRemKJcX
yTuXT1/P95eDE8UeIIdsWjiaxDXaNz8CNcXqlQ2RkXKAZMpXebbOLDVIGtd4ghpkqcrysB6rXAU3
jjnv5K2R3GT5U2euTZ1KrleOKAuhpEaoh5Xns1XxjZ0Uj2sx3uroi8x+0Kco80nx+D7ly77eAwVI
HoO8xxW2DA1WczfsmzFZ0teFP6evaRMqT68DDDw218J70KmLtTVyaiTDOn0r/6dNQmxb/h4XvBgb
oPEKmYG8F00gxoCUX86bTQdifQlXWj+cj+DdwxLUeZLdPFBov0BUFfFEqPN3PYPmUwjemeu+vkP5
yY5OphvLHEryRWNM9F+oMBgM/EkM9qyajrT2OvXUGoVwPdJQ3dEJxiycs+OfGtnfUSvNaLh2XLuE
LwEQ7eh52iIGjAZjHGOL17BqfKJqRHO6lbtRRACCOmV2A6wO/oxGaMxtQX17bNZUcpg2LVCsHU0c
/HjVIW4sl2vTYbwCvuixy6WSIozmr9WarjAa720SNqldCNo3BC0JnkaDsp5/10jjF00chhjeAaDO
m5sE3DySmC9y++g1L7NVDBd1iTjX9JHhdONNIfP2auQmKdjvmpY/0KvXhblM42amueiApvtXM8km
UvoNQzXR+nJSjxjlHqzTC+VcHVYXEauenklPFlZEc1Q/9HAoBoumW3jiauM/w1RgVPCXX+3Z+77s
LQGWh3dGmkcBPgk0tKRFrJOXHYgT43FWADQVDlafWppL7brINh6JCEO0kXiQzKh9rif6Kxt/7Uzl
wOJZFHvQzJE3/r68vq1qGKRUMD6xfdHlHGrbCZqcZkM35sEo6jSwusXL2LLApZVVNo1fAcShNay8
1nFVSAopy7tSzkHWKI5abNUdXiOizx7Ahri54ZhX7pm7ofEGuW+QyLSACdOzy7AAzMrFYYOtGxqI
lihoaRYF9ksJCoAiMenhz9Jc5NZ1GICPXKsoCfsOLSSBdPhAa5FZA00PtcgHS3NwoilsJTKM0dL3
BnETW1BNqrnV9tcx0bYPqJaJBIEsjnLsJ5or12Y7KZ/5YAwV6XwBhz/ApCjk2nKav+jIa9/kfPkH
iSvTcAq55rH5ZeGmdrogiVA7FX6fcuvbiHktSCyr6mZN2UDVeJod5xOoBOKzII4d95kjwFPkL2LQ
CbDJbvTkgOodFC4y4V48zozbO/uIEP8hnly8irHdP0iMPHM9dWJsvp2ka45Ew1QAw4/glWgv0NFQ
00V8VX+P9DgUzczsLYFuQMo0nWeUIZSO4ZcT8mtsY4BZg6a7yuo98Vipdk6Wrtd0blOS5mDxBw5E
eEXjGQhjQzg+xU/trCgRwA/0Up1JLruoGlEgs8gw1QgRqVrU4y5hlkpGw/7jfQnF0GJdTmReCkTJ
zN9oaCH1uKNnTBFS5TFWPLrlfKroBmsP8ndpE0bD64fxQ2mjynvuOpaaWA6q6IdAn2KvbqWkvgJg
4Ocfj6b5JPtbEMwTN3u95VsGC4SZ2WVasQg49VAIaJxKoXq71nrIXLT4YO/EEzOmrW9Pj20KqdO9
PR+9gt5INsVNn8Vcerht1bSYAphTKNDfxvuE1oTIOZ5I9oVu0AZNJtj0kJD95l9QNaRiYjKOzjzf
8ySMB48xtYryZw8g9vQfchPCqxkZRiF4AjX1kQZLA1bw4W2uvzTc1TtbtH4LRzQ8IcdHW2pEBp1z
X6BHx8KaTNH5uNlPBIgvizDwM5U1frtG91KqAT/0BKphXlEPTJXNq4ZpbKk41uQOEA2oZ6peW20W
4ZdThfYwglkuKJ37q6uZePx4BSWv5VD8XVtsgqfzEu87gLXAYFmmirUCUYLErFu6KniiCyG8Md3m
dmOYFzIoeZIJBmNq7h++8syfGw7jI0Ef99qcMEYDw4VCG8OMv8bSRaA2v6bTZGueohuius3cWyxY
AEdbQdblZt2qjad6BwOj0eQj4sXl8o17sIvaLZFfmEjUBIGmSNrzVc6F4g5jk2jxEe/mWsj40GT7
AMSc0pp9O/r/rVfnp9aZWtk54go/ZyIvw6ux0sWV8sNbr2ju318KiA0a7Ko6mLcPzJseHdgU/eHk
TMUWm4CpYClQml8Tw4ELWAvYwunFAJt/8XVjc8b5Ok9D2BbGXd4dmU25ziDBB5u38eB5mkA6tPqH
8CKkKkxnvWItm5I8TAaML8nJ5pBD1ITcuDsLPHZSrrs8Cqv1tpUSU7HupGQtRnHgWCaPMmm9ULae
xzPzth4zKekA9CVYzTttj2fD65gODWs9D5d83HDA7umxnQjWHxxPXF8iaQdQb3wsXFuzQAnhdx2h
UhfXLcUu5OxMhEdDerzY9VleO8uXB2Wg7WeJQE0l6m0RtSJNEmFLRpD6M2m2fBNy44F/TYzNoAbb
4WLbTfarl2tLZq15tMphT/H/VRyZderr5tvjLBVO31VGTJzusyXRVGVyLisuiiPmY5yK5YU1rjm1
KyqKO/nRftIjWV0wX1+u2vhGlmsnX7fDho5MBoMnURrFyIa9DaGQOwA+74zwS6BAnZ+upJbIc43C
SFYu+kANHxk4DCshjpJ3lXOmeMezDOp/AdU1S8oSb/6Bs4bh8Sn82z/ZVnJt4UhsscnT79iT6zd4
bqP2tLQQL7VrbhJ8jNh3+GKLJM+4I2VxjJsONSZpelx4DgNTwQipNMiCsgLYZR0X38Nw2eE+Uyy4
JW9px2xEYassWLpG+izk5kvaARy57XN1b0e/BxSJKExBdgR74WUVizTNDYaLTUeHWv0JCGT8K6iO
2Wm7xjfqCDIm/faOGcdZF6qvZx2pUtISYC1oOFBDMfHjsrERpawdoCM6iw3un+4TXts3HMhHtbdK
KtG6HyI3PIYiFufRY+5Ui545f+9EYeDZsHG0m1/RS0Kb5veRCbjkHruOGVWnuTgcDRR4ZWy7TXW9
JrcI02PpdmVQFHy5motaO9Lo7EFquSLVhzXBQLBSkk4xfg10YdCM7Vx2KBSBQWRWfRFOCtLMBMJg
XM3AyEQsccuxzXfNf8Hiz9bd395rtGrByeqY+GphrgTcV0b42jr6e1Msr1RtH/nppxfCMg3k+KEm
55EUlmLeCS7kdK9KVJw5d9Dw4Ox7HHseedvW/pL9PEwI9I+3qG0SuYsQtc4GwreJGSsUlTxrpDCG
tGUFNTTIi0nJIE+BMzO7mIxvdxQwnEE0G1cVLS6230o4w7YXikXyzeASQrxK1YI0+17kbniWB8j2
WbxemmFjxjzwxGbe9XacYv6sjPKSVZ3iSoqXOZB6K37/mj4eExINfamR9bqMGOvXymNeM2MyerjH
OTXXSMkIa0d5aBEGUj5AjTYQHzyDQC068SZOp5Kk5/I/lYuny4UNs6GYWFd4Co77B3Y7UjD8VliA
z6oqbCHUn2xBl5QELjHlUX26cP7hWWHeTpmjTmEkZvx510NayXoYH5GDBSnqTkVRAbBbw3Up/c5o
IhTtpLsBYzRtc6Ob4u5z03BiMOfQ4Y6mHxoYJyHau0PYzlxgCN3/nVUn48oI8ww4FwSojlyAeCSk
M0c0454W1qdXuaBrO+Igqt0GOHVuBo1iav/EZV4ymmgkFrCfxG5JKxXF/I6rf3B4Qdwqzj0kTosU
h2RLb22BCGFYj4/qjoD/nS+QRg0581aNLSHfFq2L49e6FoyTaFQ3bRJMoa18BDfHQnlFqx5RGw5k
lDvuwfL7ps1ncDVyPYmU0DSTJIWeq1ibjSFmja9FMhzKOItVi9dmICnktn4536IQ2yYAalc3lvDF
mWfmjiZmkcuHXs90zA1AapvaKIHPbNDQnxHIfFLmYfot/8K7d4NnyFyuZBuPqGNyVPsZicDAlWTj
S1bqtL03t88luRA2l1ufNBnhNkSlu2SUHh+MMHmouSxp9/r9XjeMg0h3FUIqQ5l3pPZmC97A+TxS
I+wvBefif6qwVvf2vlk+0UMZzYz86Kz+IDg2UO1jVCu6DRX3FbhE0hiSxuNYYTjwCBQGRVFcTOVY
s+B3iXDZMZG/fJm7Pt0TFKMbkmZYszFy22FF3ws9lprc7vaPuvtVAAPxBxJJ2cGTXU5XihiA6mKE
CVPaQd7wn0ZtovfsYX+piabjZ4WF0FPBp38vBvqXh5Aw4BvexuGw0TjMld3tw3cZH0AZrgrCzixs
T8kKJrUfCnmILbmelR8RJxtyW6KRvBqvtEAW6BSsVcThndOBrlatB2d3/ob9iyl5JaEPowpf7bF0
oheqZTqMa4ZnnbwOXRVLa+lIe0eJUKZUtMk94iyrdiY41nxhjGOkdfIsZznwimvOZxExZfOH/9OB
xI89CHyz9TdTbB9eCXYybGSFcbpBzFEuYm3Y0GfCnxPp4OZD0vLvzHBhJB7nX+LwTALrRKiQOyEf
JQiaDr2E3KvGyMFBk1MdCjXGSu/CliVVY/u0igSSWBhE/M4MkhL4BJFShn1wbHT82GCS11nlO4cf
YEcUQ2ZLZe5nXzV+RJcDwd9q+t4a9a6yHy7b+3n7mgiXDQLMmI+gxE1OV/qQqE1Q0+mmaLt5UldA
/xrE8vTrli3To6atlLXtYksZP5UHRpShe4MfnsnNOzO6xv7MbVP1XI2cnYAG5oaQJj7N1OzKKP1b
7Wfkt9H2BlMzbGwBtv9ev78lsRhMKbssH6sTtAE3iDHwz9zptAzMaB1TnFn6Ph4bD5bItF8KleQQ
0D89drUOwdk/kCYikoKyKkWCi+l5Z8EuMGwEZsXeOXEqif4PPvOUMubudnE6mV8uPYYaGk0dKLe6
vxGZ8uP33Sm9mmPMAtXjkw2IbyImgIgb1I0UMsJ4E8oVXjM9a+vf2Tusu74zH2I1gsz5uos1x30j
ykYB8IyeA/NliWz6G7Ypiz3GpeMmeG8reuiftPcm4b5Lzjhqa1SDj8IJILIjlOaeVI8VoZeNxQS0
PKicWHwOFKkw/0Rbpiwysa4yBsXh4n6J0XVH6tkk4JYsbrcicVv508u2UHqafmLsNkfu7XbEEJYh
BxCXQsefLulnA4scU9ne0BD635S126AgeXEk5gQpcByVDSWpREZExsaABVf80oZG2yFTWXp0bWNB
XtaHMNd5sIy9vlEox3Cfr2pymsuppCdxJcAyYclMQsLQ/NT5rhj4UtIW42AnfzvFtd3U4+9jF2xe
oQGi0NyxJPxgfNLzEm5gugAKa7iAgHFBRQfcb4Ac/3DGUp7m24frcaoyoBpc6cfSLGVScTo0faok
sC7VSxetnymmV0jUvW7H5H0yF/P6TVaSxwm2dn69ffsFDEgziLU31HSUz4wKW1l1E5cK8bIxEnwb
T5hSzsqCS5BRVccZ9EtZKXXpkoIbZEvZ4VmBJfAnPSRPMER0c2IYhqaOw/yyFlyDOXAWizmqMl93
qg5c07H6CBNMMfJlx1LcvquXIsNcr8JZzhkSq3YuV8VaC4e0KdhHyW1cg2gFXd9c8jr05hPa4w5/
l29R781Q1qYwpSh7LBZd+JWDLthUm1MX2gEokzH7yw4Z6YvLxNXWmevnfi9VZb6+BvthVCixijTd
DdCp9MMjwukkrnYoCbJRXE3m22evZ2KB2/bhL36ZA6eyaYn4WXLoiw4EPvzUyanNERYLX9/4BXdh
sw6p0BtQXOZl0WGjkfkVtGcaMdDOXcSawHJKu+Q1Vc4WVLdHdHeVGCIwefOBAgLMm/d16J0QLzvV
7F1JCLvVavNnklFX8cGykdtbGXigOQa+0SVTU0awAAgyRC9ySm9xUHnMnOYAwQIjpN0aE5KCONaa
Snbrs9PdxMCva2z4tOGd9Ge/bP0m2PnoSMJrhoHaPTQeHQwncutHT9nxvJvW3TVE5ywY+w75etNK
NK+OluIaMeDbh3ZSXz+X3lISoU7o9o/JeCiIM6bprZt058fLpp2HzgHHvX7cprgvOYvasOFDptZV
aOdYhXDbdDYgnFT7EflkQ117Yxe31ESmy7IDOtfd8icS5TIbqNrPcJam4isx88ISlOLXsomwP/Om
uU6tS4ACRSEVfaWUIVGAllidnA2C5/X/D+EbJiQWdD5IHNgXwVWJHDartJMbf5JXrxk89Hpd0U4d
MVtLsgC1Pih2yaJjk19DT9MqyVhGMC+BLlXHgVKHPN6smiXO3LpTjsvJqs/55nP1ttIvuKNBe678
tnkufb0z4/FjWfnSyPdoORbh6/J+jf11CJ7Fm9S6XHRPLmy7NHmpeMErrPDNPBl77m6GUwLWVKfq
QoBNFXR92tW/uVlEuukk3tfE3r1ou2c/ugiqXhdQ9+0hBDVy3J3Nva70RbIhkifO+0Poq8FkTCSg
WiDVcBfII5wo5eokO+2KSuIhQ1LOBKzHHtn7VwFpkPDE/5G1HPS+YYu1hGngII9FLh2eyCfQiE31
HArMFGKjlAZnjPwPuNCPwf7KiWLTeQxaydi2y1CVRwFU1xz2ybqA5+9/+99FYuBkrRWsnXQmUTLX
m259urI25xm9LQeOZE6Y8HnmtpW51UUEzvNoKHv5JplNeCwK3uFJWIs0qAHsn7HAMWXyKSL5oP73
5S7MtGDoE/d17beiaUEj7x6GKR0thI7h9R4IbLFjdYVxAf3VxqWoJ2jikofJU4HjDCATkkaa643T
8C5El81aRmLrul8zTpA1Dtq5jJQrDBfgdsZJ64xbICsc7mvvScQNO0b3tDqhplXQsIpPU+B6AJqK
upsuiGl7am84GkeApAYogzlZ/GPQfiePAgzPoYTOVTrtTbbWsxM8QvtdTn6omRqxmpPEeNQ/6qvW
ZOsl4oZ8AJhQ4u/cPrPtYkTgSxgWjWBbOKSMVADQe9h2XDphSPd9ddbXQFCtkDK6RosZxIHSohoR
iWEHVKdPWzmSZ8eS87yxM+f3fbYpMGilZEKniUonrRkUarunn7Hi8b8zU73Q0XW71GN1jkQS5MiN
DP1UkXG6j8JcH6rE5q0YDW/jWANq3blKETl0Y4SCuE2DvuHXjwnK+UOnduOpt4RbLh/JojVDQssO
S7xofUb4FhoKMOgYyAHb4Hgwmh2sVOsQVC0OwZMjVydOmel0ozIEiiXwoY9xyfpppJdxeasxZ2Kn
OA8wWivbxBrqYq3AKaspQ1PSyY1G15CjJrd0qehrp6xZ6uzX8qTRCX6hpUCzSwvEzqbXr9GWHusj
fIi7x2S1otSOyniqB6vun17DIUx5ULEe53+D8xMce1Nuxfw87GlnsiIJBkTEl2tPxBbL/4xIJjvv
lXtWruegbUvDtW5wJoA4ZzEJVo4x4XWSU3n/yEuRLAoWLVDrdBA5cDG/CFPj0nOHG3UF0aOPM8vO
W+cMfuh5T+vcNqDMMaO6SZHkYE/uHF7ZRyC5WnpftJ9dE32yENRxh8zkO/nq6A1CEK8lHKh5eOyB
McpF7xHUya2XCpLR3kzU6VgzrtLuS7pX71D+1g7PCm2nLjlZJhcZhG3anW+udm227BXUzRLto0YP
z0/n4qt7mu7NPFdhQsLSZAAu1848Eb7SHy24EPvpL5tFTcTSx5xKLbxvH1x3yTJuaS+viGyCx0ZG
ygMJUDgAMh7WCYAZ9TFcyriYUbDcFpFMKtbpdvTzgOCu5JMS7YlQiJX2+9vf4RKqlRha1mfKr6AQ
Dx9412TmQnWdcP1oZsipLmHcNv93Qqu4unJqyMR5KGFibsjijiUbj3/rEQlYxo0E3G+X89QsUxVP
bdiofe4s1nlEFeixSQZNaOl1cXvogrZ/Ms2bmeVUZI/k1owdgWSAOAs1U/Uws3f9TPT/If33+JUL
z6qsTjQALjaDJOqJPMrA/B7lirOK60jRoZOAtiHS6Mgsd5I53If3Y/lrXmu31W9s+C3ALpvmM64f
9kUhpczH8ZCGgFyh3275ubfLE1EWtciVZx5fhU3G6y1auYDhO9X7rj0K8+p7JesJhp0dCgkhOfBw
hyL3RBdbW+xARyHPMevQuiEKClTP/3xPpS60GEsp0YD1UQghYTHTjFLy4dyDOaYk0QG3WuSnS9p4
3fUmv4idAlVHTEPkw7M3jnJtaHRJkh8gVmdsoQXhs74ms/0k1MB8KOovVQWhsAPvvR/GBKjf7whB
5kRYoUCS/F8KoyN3PD2cHwJs9q5PpJoAU9+FpTbjWCPXgQalnBU0DSC6bx28nvPVZQYxMajQV+j1
j2scTXxaIz1drhxahEfLgDIqTSXT1Ky1YTif6Wef0eeQf89OHLSS7gbXiOnT5JwxvfLTrwwfqBEu
RShbCF5BQcQEp2nEJCdgwWu1zhmzi9iAiDnbNGx5+TaDsgl6vonGuHjiponuFAzbTfJtseFo8iCF
t64YEzB7XJf7qtsbVrHQ6mJ/MAYhJstUNfJX/FOJ4wHJKBj6MInsdBBC1oTnK00HU8LLYR1OIteD
z5RUmBiKjtZ98Vjb/hJKGX8MXF35KzSgVTcXESgJys+Eav97CnM0gdGxh7zfBzciF2sK0xJGPxMD
c2X1ApHhf7m16QfDYLBq7GXL3XUVoWyDHvi/R2Ja0EjhpYO6NyFX+bS5YLzTb4jjT6z0uZ3IhRWf
Y0Jv0W0/Bid6nIsoOwTknM1PSna/tJ5I0WESgCNge3JwEtDR76RAYrmJdd8k4FWJxNjF5y8b3SKT
ga7WoSwHzVzSfh9VY2HzEC0RurNhQ3Oap4ytjnvGINnDcn7GZeo124TB8aP4x9KVAxKyWaMd3PyX
eFRIe+lDliYWyZMBgxq4hr4cF2OlQ8XQL1xw3/yVoR0V2jNlN6o35xBF7JHWFpS8v6zJ/qofejlZ
ni8NlzDlhH6id4FaLsSb6JGzNzB9SEYdLaLejMu5mT71ZwRz7fV9aK1ezGh+PbMLUqWaYc3EEEIR
QxTHkzR32bOrxqeTOA4XQv00Ue5AbdcDPIwmv+J0PCXwktFmj0/itEI0Uvr+00EwQBM/Lw1/K0GY
qjbexG6pI7JpVm7eQubG7VIwVSmlY8b1hbar0UXBa1HyhLrMNl9IM0+bj63W+znZBEQU4A0iEJv1
x4jB1IPJXS48b6ElA76IIftwxaPB4M3vureeT0YvBh5SH1Oda2+1QUpxyDiWrPgx0mPpMmuJZ1Sw
/6oPIsj1A02LfEb6m40dAYE5GOj8XFRjtB1tR5G6bFh3WXsX4Uxfgt/uD3QEx/L9tO7s9f2cpivJ
HTc56ZKHUtskMFE6jKaH7LvZ2KVNxCoETUnWEHhl3zdt9I9Y4Kj/uOkagLmDcUXdUs4VWR8Viwcx
y476rQTCM9N4CQYp/ET0fgIqX0al21IBpn2ZnYV8i+GNgIWHwRGsPBCyM/IF7wS1YypvLWb/2fTm
HQqt0Ggf/FHxpHNRITm6euZdiiuyUHHTNwQuxUq8beJcVy9weeN14iMJK+CaTHBkK3TzMyj75TIv
eGmVn08l+8p8Q8FjgEOQL70IG4DAyLYM/ICU3clGXr0Df00mLfuwLYfJO3vPo78kTIn7blp7FDHD
d+dvZGC9PaSqsJv9a9ECkhd7qFUDRyyYHKF2MlhQJKZhzuLRjPsC2G5hre0OysneZDowvFx2CuxT
EUWLg0Z8MY+Fsg00fyLftOrP5E2L7ls6Q2DnQ9Ma5xvmW592dVSVwiaRZWoMIKUw9me6GPRca+OD
MQP3ta/qt25CaY2TQs4Mx3dieghnTmAdkL87FRAKfz4EBGf163GELJ9QGzgzSW4EzC6gnLSMQehM
JGxRyJG8wN0WsBKL5MgchuwzvSWlofLi8fYdqJ8uaexmsT615IrseOkoLqbgsjjltLfa9h/RwyLn
2Eb34Qffg7/VCn4RZTZOmHyC0X5gLfSxoo7k6luwaBgGvaUyvbvED4makNE79op9rfM4y4a0OTOy
UQit7RGB+qREFzyLi0AzMxEE6ruGUFHWf7VGFImswdNKa+MML20FpZsATyE81QyuouhCFOH58wj6
+e4H/WhHAE+HFTrMv+KZhRtlWemh++UbovwCY+TwElGbZ3EQU2RjpCrlsCPlY17qc0FLMVYU9MFo
Sv2A3D2LBIVINyNAKtVDEVFaLnKLFC8rm3GbU/PnbBx+in1NvZ20FoqMus9injRmRwBqMKaO/XxO
QxJIhqiqIaW6iVg19RtjQDMZq9lTS+KKDyBMSC0nYKwfFrsvb8n/fZe/XcC1G/AR6TtI9CUwKzub
jUISICyaIz154MMv5bxmeDqW4rq+cUuUMs4k9i6BWEZX5G0z8dQbo3QFe0qhDOLcd8pb0O7NjVb6
C4179GOPW+/Y5piicnTokmPlEKimhAuYBnjfGWvVIlldtSDBz/lKKkQr/eEw9OyXwpsDO8SIJ9s5
KoEeSwUiNrFOCzeKb52zXW+TQvD8Ueapts6Hk4g6tbX14YIfezO/Kctig3w/UI95X1zEyAs9jO64
DhIFzFmp+eyibZwOTx/9fWlIUuplM1jwhyEspFu32C/OzwbjAYrYvwsTKNiWea/pgCaBEn3laQ3v
HQAVMHG5hBVRiT4gcKnwoisPFrhGqszcGxLZRuaE6SQF+WrY9QZiPwQrJL0fUAiPhfDbSHRgRG8O
J2bx+9EawO3q7//UWWu6r3RCkvfZO5cWPYs3h/N8kcJdAltARt3Z6HxaJALxa8OeASqapTkYSvk0
wSnRDkJ4N2DVqniHxKPqU3ynwmZMvDmyk7o5lPO3qwIxbTAYKEZ4CpW/1A2M1sQbl3gpz0B1b0+B
MW3BC2M+ggyrJlF7sW7QL1jDv9TedyhT93CTTwa7OKbVubruyrIc8Jcsah4gD3nqg9cBS2ZnR9ct
aIzgIiOHQfjYI3+Ah5MuAOJ3IHWQ7W3Pdjw8jyUYPtvzuF9ElRpDFj62+yzO1kYzEg1beZ6coNU5
vuorQFC6ZNod4l+jMVPqNTj8wR0czI4UIAn0usZJdnkCbRfQxHlk7UW25Bs79vvM2YDScNauK6/K
ocR6g9DrwKYvbOlbw+9CDESvLx9ODFeqkvJ8p+6OX/Oj4V0sWN7eGtCHG6LbxSi/dbluRKmIU4u5
2u6jD4wBFT8bo+F6+P8FNiy/GkchQWQ1m5igDOIiYQ0RkMFTR0UfkAHBggQgdZfHeJtbjCHhvdCf
H6yaul0/5LghRq2DNMqSunBd8MZ1e4Y8m72XMqa59OgjZnEdfOpODVn1kNLdWiG55B60PuGZdZHj
f0sPW3JekYYJdZd5h73qrcE9HhXViW0VuaFZdKol9hjITuh4SJaJvj0Y0y31D5kuid90d9v03ytp
EAtSkgnKHYkP8c+TjalwKe7/33SDk3hMvOVYSHezKKH9x43VOb5oulq6EUv++HLVdonSOTDDPoAY
oqqeXepBzi3GBw5zMuyT/wR6k8h+qWZLgt8RJtNg6WbwNIN+kaWgCT4fa6g1rOxUqRwyzD1aWvsp
neqWSdPfAwufbA88gaDh9IJ4pB7dbIMb4Cscfhu1RFON4ci1JmnuTLc40cqg9wjcKAW3BhiBeo1S
08022Og4AgYZx7WXCHO2y++oISomVuPaw0ymDBalLJMeVzolIzCUOvQJxWe08BaRQUnf9l+VBMJi
H5JnMDWlYPJ8y+ImNxjh6/fGbYeQOJXXUaa4Cdc+Yqq4yu5/4Cizi1Ix9JK0UAr6nyqCOXrwWrFE
LHNKgmnGBybLCksV8n34mS5R4yeXi0U5OKrw7OHeaHeV0VsYxAV3tTIk0WPA4bviqNGOIjfJ54Xh
aIcy27z+47Eepgt9D0LxqOUJ/dQi5rs6ZXK2h4J6IrQswLKojii2w3w8O7iCyNvgTrO9uYlFTNPs
+Z0xK/wwCAzCFE1cSnEjQd8IfAK23ZGRnvWfQ9EqY2clSFQ57QTO1yfruEWzWENLdss3ZNqRrji3
KT58WdAacbvPr2Zi6Ig3II4iy4JM2WLs0NKvA/e+/mJQrukVnsJHqY72kFaO23/A4hPKR+uk7JfT
BqqZMbpxLdd2bMC9XEiJhKDCr2vB6aVeW9frfaKlQDhUeh9IuOU/M0eObFJXWhPga6tPz0Db2RhV
psQp5TWfaAiiFhdPosCpB2WKbdO0CGFbLeHl90ep638zkK8k9xYxmtOqO2I0F/HwhRKTsP6iZk4E
6004kEDCcj0RvlzkSxOKvE765c52lAUt/JQBddSjl+jKIiJT+chLm2IN4fTONrP0HPzHt6WY6Mc+
gNlJIOiKjwlUm6BgphGKcWIkICxAZ1LziZ8DiY1qdgd9KIu6Pi8SSLvvXpdiT12qhRq/Ld+M7g1O
+5wmKaJdjxWgFY2uR36aIKiWaFZQO5CH9pox1eNig4bV4bh6emUnE2c6IhVvfWrsR0X6NUekvwgW
zRHIkB/sguJph4k+kYiz5niqgiM9/cZVgqw7ynjG/idTW7djArCnP5YQDifKs0Opvb34R4E9bige
AGCXP/PFT9My+cxMHBIS6FISEKKuqh1uO1c9fzelWXVXttFEyKCmUEFVc43th7f106UR6J1RxXQd
78LhTrTXQlpsRP5kO2Prv6VMOB7ik30luhIAvnumoidDvvEsdGfeg2E4Egvtjol1SF28Qmsg6EgX
p7/nHM7fbA0M9CgNGitH0lJK2iDy7GtY6zT0LEV+7NrGxxqaJYdP0GZ6uoEMRYT/OVLdcPnyppec
6SJSaomCZjWTj/VZw4mwyDE7ro58F43Ah06ad6TF+66n0XSYP0fKo9vTlqh2ida545HVxFTYqdcs
YDji8cQX6+7fJl/Czh4LMisPsjPP3KC6G9/XGsd4hmGyDE5AfeqtBcoVXghWW4EeE+tSHTPct5e2
F/sEh6mEdEPo00ZgTfgMh0FV+EAQFkHQcrPrVGCeDZTHwIxIJF3bJ3g8V8wOTUP1+mjcjfKT8V2M
UCFOMHZmWyrpA6+tgbL9Aj2kCD3ZkIPuQ/X0S6l4doNIWVW9JyG1q9TjhK7WBliMLnycQLlZt0MZ
9hb+b+OtHxwFSLCqtFBWtflhOK16jLX9rflO3797wpmIcYqgBIoJKHPEFYKioo+grQ9iqsCw4Gtf
vLD/5ge/1jRPRuDIllVBWjFyENWY6eeQ6a/KEH9xB6bXfZnkAHj3bJuNA2i2kdVvENlXQ1t9saG5
b5+0e94OsAWN7NhVIDdsiet+BtDPuP7ki68dl+W8W0Y6DqQUD/yFicYC3a+5KoBSBM+T1BaLKguD
it3CYWaxkDSeBnrl6XFi6phrH0H1DcPlri4UDLNVcRzHqcVWIRjgPztiC9nBzVl9qWHkeYmpWi1L
TRa6JpmwqWg9OYmWllpV+M8ZRQ8ME6r2vxa2v+s7nzV9dp43+EAhg3UxcmG6XAhqokDxCpyr1GQV
jWYeTnaPNNzlu3hNP3HM/eug+FSNjZrBK3dyRSRsH9fAnTOV8BZIaujQaUI+ZlyUeDCQhv+aO5z/
/QEuhXw2oPDQzhojke1AoOoY63lvf+7J3FKvHdDzoBzt8KQBSebVbIacAvfxzFDgZMDesujcWZDd
1pexq/zceXP39thkWtK9ZCR3muoo1HCiHT2db2sHmWlbBwlGHPB+WNUijJRfjj8ffG9RxPFouYwn
QHlKv011azEHTjMq7WTKX1mx6N6FJGwPHipznTDSez+0tu7HPB1H3G7GaE+/1ZfP1m4SCMzM1HCs
2hik+wHr72bi+h9E6/u0LqRqCjVAcGJHdUMOxpO8QFg0S/R+gNGmDdLL8rH/WvpRLLGbkTvmYtV2
DQkD4XMioAlX9QaegHqlxXz11c9uUGwtjr/mZExTsG2bQ2yvNfYSc6IIWswuScE2Tsr55ud1d8/o
Tq+U96CNq4LPWwXgXxdgKvIv+DsxwzR9lLuK1HzOhA1Q4xBA2DXdmAqWcoPyoEQP50AJkJIMujbC
1FTNkdwPyrsdsBdglExLr9hK2YZ1SkG3KcuoOWucccI+aamv8d8cESZmAUR/yyXU52XCaI4u7ons
UFVoO+F7veu/jjUJa1op9/YeNDv7ROD2roRigbVCGsrTA7WkG1wO1mIzZy0KpIWPdD6vn76iJVES
NFdoLWg3Mu6xBHYsIJ9RShmrIr8IjDbwPA7gDr6B1S2Mpqfjp1vabmm4/0r2MvNPIXfCT2VL6S/m
qso4cGeW7PzWVY4rNVU8zZOVLCjsUZylwEM9+9LR1FpeDZ9zPtyQWRaN+MWu2vsLMYmhvH+lgTPo
O7UCqk1MvbZ3JTtA2m3Xh9zWe13jgSuBb8DXCMzGmvy61FCHTH+8wtctnaega+RVUxh3iFrUnQNo
i/4xoFjzPVqCCTjmFSNwGH3EuKTRGoNk7MbonRDMU8pUNhXhWVhGxdUgazfiN4GTzInLLQEqi067
QzVnjYgiM+QOd9jGH+uwyDARtRlediahn9k/wCkDlTxBuhxas0YTYTzjACbQ9PJ7297s56X/SPc4
sXO4eWX+/mZ0mh0CuZXoaGphE6Crrppd58cnx7lj8ac+vxuYrqQg6EKOxmCq40tgC4cfHMbSTGzm
dN6YZ78kqfwkrg55AAJ4BZrrIDK9cMbx4FCC5662Gt+/GW+q9dAkhwqomX1Q/H+zGptXwGSueZrg
/bBtnuuQ/WyZPYF9nEfAGwGQFtc8vX4n9TPRW7hZkx5VSCVr4+oGzwm1+0gNodZvkY11lgB6PnLW
tnKOSa1WlC/pmqLUMmQGNHgnTyH8e4VBv07vDESdsUGk7BuI5eYFsObDnInAO3EDIIIrK98HSywh
6vld6/rW4GB/+Ar7TFvBGkkotkwwCxvLSjhpqYV3GLmZznzkblSbVvX6LFV9PXY46WWkvbzVFgHX
jreKFltSo63X+kcrhZz665Z6ddWSKk9huFPfQspiCaM1Gtsa+d7wVbnjsesAfEiGBF8p6obJvNVm
Bg61eAvP5TbpkWzrMlKoADA43L6+OMm0KI1lIp+nsSjNKwpEaJZSzxWO66nHsHjlD+nRFVUA/fgQ
VctZPmlFP0CftzDP/GfzWDNK5ZTR9yJK2jX4tFse46Urs5Uf/RxB+ZjEyGUBSNhRPR2ZMtwiF2zV
fTl3oNfnPlTVldp43oTJDdnCgw9c44/iVTzs7Zddu5kMmlsOxveexC+tfyApJLzZXq6xsMGOh7UB
wv2Zz/Mz7cvACtSdZ1pS5r/9lVEIVpMqhuPM8EqrmgJDj3v6ogDfNYjadCPC5oLsnfvSAwWKsitA
eehIt7r9nytdpayoUEx2GIJ2DuMzAhYPS6BsaPxX4rt9c/j4NXGlf0kn3e2fb21rBH/W6+2stjUK
nMxEPCpS8IMftblNP3BHBnFds3LyKq9ho+hFCGhqJhUwSLA9aa6f8TMWGumJmk2htLyLmpQviWYa
P3gUhJgj/K8k+14QByGaI+C6LrlDqHEV3cB3ZuCh1YTelNLhUpilv8uITiEbfQSKvB0vHbsZKFv2
4lJOCdvY0VFXbMCCUEmCGajAda9tMIbh0OXf6wHC08rpvEcdKomv6QeQMpqSwy2/eW4lDk2ZXXCR
flpiT5aVb63vfZ5DH0iJRiN/AaylQmC+joGXPy5SH7Dj/6I74//eePyp7Yi9VQIdByuqf43XEY0h
ti4ZKYM5VC8s3MWtNYmiW+CvAyRgM6xOMnqWeIz0xWozAyn8wq2FAOdiUeHt0HIy9Hj+oDQ11BFj
UBeYiIoLM+7H8e1MvhoWVyiOwLTHfpFJD2Td8m4hsuwDmCBENla4g9I1mXUV5WTUmW/KK8/SSj+W
cNrn2O64GB6PyIkX56aqFbEGL0Nez170HI+hXJ2Do6cO0x0SoBep3eNYH0Akh2f1pXIyRugENcTY
rSmPBvJnY7UXFWZAPMKT6d29uvv56B1A1JvvUd65BbVtU76pe43UtU5b32ITMt7yuk2NLpYor8so
7O9AjtJGlA9ralMiK+/MX5E8+Zz/3yIDwuCsbFIyBuUTitvrpgpCSCmqI4ZSuWLYXu0z9FA17Vqf
0Do/mdDfkzh0Ye07Gt15T6tGHbPFHEYOFj+JLVjEiX2YPOsgcstAF80HGjjg1kbMWBWcjjU2lB7Y
25Z4hhTQV4jlaREWdTJy9w9yNO0PhELaftUsxjRNnJN7R4v8/iagV3lchEl2xrK8a7lZCHIodd8x
Na6wiVAUwnMmfKlOyeR/OsXqWHbf027c/wlEQme+uSnjnnQeFvvHjyhjHR8+5T05CAv3yThLpwy0
h2vWZXhLoS+Oufyvp5WdRxbOUUSdiEuOmu8nE7FAYxWGINwvorAHY5wvGFNnbJ/qNKfYLed36ExG
MkRsL9ZtSWuiDmAhHJMSFHXS5e4+cwfofH3oeoMYLu+x+J6UmcpjRIKBMa/9XP/jzeQ/KyvKenuD
9UMqP5i0YHQG3FuiB8sQab8pkRsUbCEwwUkK0OJdDwVzcL3sTJjlTBnjRCF4U5zt3yE2dxsMitTP
veV9dx+18pioQrfKaEjIEzVRYcKckWM6bol1IK8RN2iTTgpwZ79/7QKPowK3vpf22UoUjQ/+m73H
Cm8OwqXFDxD9zpxCztfRQkPg2WCa/BcR0XlKheErzuE+jcM7Wml+fa9eey9yI8EF2yI435wXyM26
SGvQPQs1hmPCtNhSst2CpWZPDC9YkjbUNtq7T8ZHJb+ZtRF5l5Ulw1cSJrK1vZaYkZVu7do00DCl
gT1HxDSvcU3ViAI9fx5lbaIyBBz4MJzaRGk9A2ayukJyVeBgbgkAUp+OJDHxrgliGVfRqFDp1NVk
TkhS/5CwZ4bPhhyKqdj++aBUqwb9Ek4Xstj67DlKwCgRVQnVnYgIuiI3SB8bboohz1dsMhLZT6mU
WH5jTtHapzrPDWnacYihaC7oemcWwH0wkgscGDqEllIPFGZT15W+XUZI3YPA3iVwpNRJwbCYY2Pv
9XtmDJ45TgT20KTU/Va23kcwFuAkD+DrimKLFaaxqEOxQId30ZJdF+SFT+4qo+fRRnX2+jx8O86y
sNMmC2z+Z8rn4SxSb4zz68+vf7WmVLPBN8MYoaFwi0B1GFYLHP2/G3mlybg1CR5m/nDTUKaMQfQn
xqTX/k2eGrlIEut21P/GWnJL7t0RsrbxS+FeyaDYkZJQh3KUXciu2/P2JlJn12rcQ3P94OnoRbpE
3m5etPYle36Bol1nkcy4pOCzrHLy/polsalX29Ep5U9tAFxMEYptwZjbMyrwQCCDlDTK1eDgtTA9
DFUcV6xnW1OKRjonlAkN5shIb5T18si+rS9O0BXQFmvP9mraEUIpImtDjctCLzzqNxW4x7kw+4dI
t+xIxC3GVQl+kGQ8NjGgwbKOPM/5hh6GY9J+ZeRepWUsjgSdcvsntsGaYZPOJCmK0l5jf3CRk/Nh
tyhP5NMy6ST9Au5a77Se1orme91XzDA8n+wWqOPqTMZt0L8WwQfXrAOGom/gwLxda1ovKPdcQVlY
XLikYY5mXjhM3HLQogbkBSjTUOOa1IKtPUrGbTGVZaebRyCE8W6j2Gn3MxJXa59xv3MrBS+P3h4a
VScqBkXLyVPQu2fOkxuGKuwsiP02F60SpGd/Wl4lBn41IixUcYaod40O3uj68dq6sUUJinUpd0Qr
Hn97wF4sGCOE/UhZkzbMIm3Cy9Ye4Ihui9zTu3Z4kC5R/jtrgtIcD4Rk+oMqbhCJ6jDp27f+yqKu
F1Cqk9HoFiWERCrxsknuGFr5tsf2IzwDstjt2NJLVDQJWTPFGEM6/TWrQ8xG+u2a6N8bb7LdSCeh
XE6SiLJCmDQv7oI+fzfWEe+ZwzPS/yu0HUMrXBfu6AmpRw5f5REABhySvDTY5++/uRgWrqDfaAS7
t92FbyvMjguBxJlqoszdpGC8Tt1jMNb3Vp/U+J6KyaGAB5U4WPGIXPwzIzXYQR6BLxwzPJMjPJnf
hwjGDLrzJOOQsPQo2W4iP5j1+S28Isox+JwF9tUStGj1zFg0eBl5slqv12huUbBKezL9sm12TWMR
QtOLoEzYEXyOw6RaylJK+426/3iwnQh22oTuE2Xcl2Tt9pjBSkcdQ74Lx2EZh1U1J5AvstX2Y4AP
JX9P4Abd2CoOoc4TsVD7FuF9kgjfDCbpUE7vgXvhzyp+lQ3qbihVpTQx51SoZMJSlrsGzcviKpLs
py6vkfTPrnomQmnzZ8oBlWgaR4rx0xzqY6+TC3rixHtZQ8crnTo3VANQQl4tyhAsz9PaDBcKss3c
4NkS2B3tM3r83E3njREa+46xXTxDEi3x3GWC9IcRmDv2ujR+snh8hFnQOCBhhGWKRiQK7wb1P0uf
5wphz8pgl8owi0IgfFzOZdAfSDvfD+zoaPjMmBMdm9FxV8lpjfXAJdRs0H2ZZ3aiJKoMyAkaFyo2
G7kBqCFBNDR+wXMxipUTF/ZQXZuTxmj7t/9MkzL9ip8CgjVZxvpDVrY4MjCjNlDi+51Z1bg8uLXy
2zNRk4Gae2GO6PfGrxqE/9s/+sg/2APXerh6QM1b72p8QNLZd4Lvy9efQj0Vlf5HwEQZnnG0AHSs
y/t5L3UX/Fe1QXvWuC3+KuPgjxjno6iF9lhXP6i2Fq0XhKAvAvgDqcCthdZezVdMBcDReTfJOSZW
X4jIT0kZA0vLSMQUaX2rl0QCnzv8dA+qBFENr5xM9SyJfZe1HaKIzi8saREP36HOxR9BwTgsi4pU
rih/87S7VvsdMtMAmVHBoP/Oklse1qU6FrvSsl/9hdD4GbleyBT1Hhu3lJiEDzFIR5J6PFpuzVWz
dachYhu7MdvVBZd1v9S00lEuVy5Gw1Ztv+yJ7nY+Q2ms2fOSUq0RWGxvWN4APZvbWLX2gC6NIWNQ
mocNs0UzIQFuoH2e3LdlnlUTtkiffuTjkzk1sg9EJ1edtPHsV3GwkM6238fNQY0cUwbKIXpt2WF8
2rmVhnCWkqZNf1I6fCXrxzZY1ObKs+egSA5uqIWTs0tUl8X40DlAQqNJSEjiiDwvINXZsZxjCDMD
qgKpvvnXrpC1Xd6Zu/XN+XDbMxhn2p4VoMxfzvoRAUJVdgWd1l0HhKbEDCuwATyiJSNBZOrgfS+H
U2+k38+7Jk7Af4LfDmr/gGZnRW4buY4tKYKUEne73bIbVhc0nnAgQe69HQc6ayUJZEjahD4axyCK
aZ9z1QSvxvFqMqYDAyUbQ2xAtcT9klZ5PRzH7Uk5jG+f3a8UTn+ckJwK3y75upgkyMVnrpL78npr
zyAO5aJ8ccU5aApe/VGxzKv0Obs/2S0rAdcHwPxu3IUlHpMmcfeRzdmvU2ZXcxRvuz0Okb9/f5L7
PcwEZsVaNGS+1+YUl5a+42qoyuDRpsq59fHlSWL0s6CMM50vtuqm07sxbLIG5NV4DIiA5EuVoPpL
md2Unj+AArS6OpqysxKREt71UBwyQbt+rbmwUM043ZIJGy8r6aJCFl1aQEKxGARjRvL9AiQ5lZnw
Ho+dBMDkUZgsxXywAc1mZTttJdA/8SKUsBA65JtTNgRpr7kSW+fDIVHF1BYrmL47P/xHQEfcUWn9
g7f1sZPkg8YLWiLZzpdPmENrqWvRdp1FVpgOwxkToGJa5pNiQyKk+QcnpNpg6daMk9zMnoaad1UC
0iKOCFFBtbJFzBnudMSq1cItwpYDuR/dTQaKduo8MG87INNFzgbKR24wB0PwVirJ73NGIy8FmNk0
4DS75ohW036T77fT+vcOtlq5WUQDnnSg/8dsduJlvJBOhtwvlNQUT0fIoHNfdNsetJM9S+2DHJfK
7tWEriFvkW6F8s7BoEml+jANqzh0Sw7CYcbE4vnsgBG6T17z9tbhlDID2ZJ1vqnMGBmvCQjYPVVy
VvU2VGGbpB3DuxMb4iyjnTlrUWKi7o1knCV1ablysETiEHumTIDw8XmCOBDLr4bTjrn2HmocZf20
aqy7EsXwY2TRDnjkO66JjDNbk0cR7z5YWDsGvela04KZEjEkS4turrMRoGHrVU6YcbSz4JRVL0Ws
T/7L26AgBHijuJnjO8c4cSylE9f2eYvHfCkea5QEcjgy8eFzze4bnr40jiF2ih6lfLdMKP5MXqud
Ie+k5rseft/66FC7OJrOC+6SB4u00Hgf1gxQe+k7+neRNSVh+8sIL2IPt6P2W1t3mqwvkA30UyHj
aIWycxY3JSyIeHgIJKcni2YelfDsEa1q2oDmANYy4YzfXxIyNw1qoQy6ZfGm5Gaf8JMs37g5ZH9h
MBpVAjR8Rx+0Nm5DvPXHAEBb+abW7yhPQ3EpxrI9GuwiHOjTQEB8KnWCLyTBvhWR/ZQsudxKchDc
k8bSECUE1sEvbsvh0qMFIPcS8eglWynKV/WUnkWdB3oATUntPHk8UrBT+K/lmjhvHZaGQtzmjh/s
0k/zAPWNxPMdF19DrJJyU9shp2BNcr4LoTewRwHS5r5Th4s2BcZQzipfswdG84WRD7+nQ1vNGHkX
eqLwEoydHJGc0GaLnLawm5hi1dKk2hGXAhQ9MpE8iNg9DSARXlRg3phFH0Ozprgv552iIWPLTZFj
u7MQAWP2DfvhR613GuZC1Lq7x3qUpU+RaoZQk9jgOQvMd8ZVTQxGUqkCRlBOCv90IBgPE2jkEHV7
1Q8CptTT/g4jbF21i5eZ15Djb/s0ZEwkQ8wc1NOj1Qb+0Aa/ehs3O/hVyvjy9uI0q3jOOhiOIJ2r
bTsRxlUu5C3tsEfctXkcqET2OT1Mv43yHZX+FQFEAraxkrT9Py7Pq6gX8JJeue5ebLveoNO9szS4
cn3B6k/M54Bm6+Mi9W9ZMVairOmEHhrmbX/ZgeRXGZ1Idb8bzOtbYSRiERPs3Uqm3P9fuq/ICtew
WI0wagt7PY7INLGNN0LXrNREM/e50DwSwHE8N3z+LViATg7TJCiurXPWqviCtNI/43Rb0l2Wktg1
Iwk6Vtx8XGkWs2qYNMwvNy3P357+gXcwjTz3hQi6davhQcYUGaFPL48SathzLRj3o/dGFwezN1N9
y2S7pHFgJBrAT1IA2uT5NZgkpB8JGfP+uazXU86bcS57gQUfmVRnuv1/DjnWu6SY7tLbFY5n38Pk
AmRLzInxnnvXCWEcFjg9uwXx1+wv8kMIuKeBrCJN5RuHc6OtGhFqFOPZFqbkbkZERwSP8XlYamzy
Dumv5BjX3JL0k+1WnHSQpRm6KwLJhJGlWUYJ+PUOvKWmMMNtHou5mi2uHXPTEkfvtysWwj8pi0ih
b30F/cHirSVlBQQlG8YF0Nt0kVrse3u5GD/o1yUgibLw9sLgDXyT3rMYD6j0vfm7X3dkKq4cNO6w
VdptCk8wEroz3HVDe4CmXi0bXyG4umZ+8T6aCo/T1UGjcfG/SHOoTJctMNMJZIgicfRq48sstRQp
aBEsquDIVclZLCOmSydSY7eMNkuVyt0V7mDOXyxR7GJidFkn78IAAaDPOtkDh33OfJffd9olAE/C
KseRPNnq8KpTYiDwsOPdRg0vx6iTclS5pBmDYnDi9KjGvZ61Sv1J6nOQWqr3TYlO5xnnjKt++fgj
GLuNVcT3Z4VhE4IGCpQzVut7knrg0ho00RvMYS3NBCNxcftifiR+tXmv0D4LuaiwW0/QGaJ0uF7Z
C0ELx98yNsU/x4/wu50tJRzXewjbPhL36JxtZEZGM29pg9f1tMzXr8KUB7t7YjuOEkiBHPke705L
L6f0UmO/u0ZPetaeAv0caqD3MkvVAHhWEMaQkrLCc7DBWVSv2mom7fMHqhZIJTnWsOC46bVXPXRX
gzobsMBUmYdVig/zrN8j4qtYoNZag9g6CI9DssLlE+EeAy3f+hs786jJOHKKyLDG6SH+RVVlIr7C
/MUGFtML0TVtdKIe87oW/hSG2+PghwXqA8L1rDKx+dfwY/yS5HyWUc9ruAbnqL9Yh2Cbe8WA5GlK
ca0FFCTVByIVvE0JAZo5DnplYwA8q9ybpnMGgduErm/QI6/EY/BZS28ng2UIx0o2hrQsKk+1y6qW
BpTtq5c0qgi1zRfETfXhm1zgZHsErFjyiEC8nBu5nod6+7hCMrT3k2rRvP+c7vaspwlRQ45EsFlQ
TXsjd6UA3sM4b6z9YLeJTkm1CEmkpEKoMtIYMNcBRelL4o6kud8Ti3LDg3zqvyPykWllA7mdDu45
XXQtbf5Vmyj8TX9JYWUNswbNKlUCj2UDDzhsPGzGc5geIH8eXEVRWchEZANxEfoqcvPPTH/3MfQz
rpbwMLY9po6mQGjkUDXzAGEzsYV5rxLQAIuYIyYYL2J94JK3g5fEnphnq/gwVDGTS25UYUtl/Riw
OaR+Tf0fjAZFK9WkTQkMo3MuqJz0FAVa9PZIx1IFoddKwIqAQIh/Cw/rOdXNJZEgMfy/DmlSqxjp
Te5hMFCaR7awq6VhjOatpjUysT2kR/iEQolz6bBFLC8Pih+SSW/ZHFxKh+TurA7CAf80Aue3DzRZ
8mId18DUFzwctPWE0XKlM87+79P34qccMLNQkQlxlu7SEvubnSc01FsrewLV5N7WO1kFlg8CtW+n
9aO8Rhpxtz83iRQW7JaU/bs+29aADBdnCTyCAiCK6yLFqHWs/q8WvZOvfBu/Uakzh+lO9jnQIiKW
RDVqbhMthgJyHMSH9FX35+lX6gyln2e3WF8tDt2FJVwlepxQ+ZBi/AQQovhPkJfisL7BlUD/BhM9
e+nvJPVuCcgjgHbsYyCO43ZAjqk+HCqojrTInTt1CY3bFzdKUIyQ6w16ygFanax9FrWDknYvDCRY
+7KECVFz2mAiFAfFTDw56yfW7fFyhcyc3YlRC9VQYKpyYy3bQBbMYL+09SsTcHi2WOjJJo0SF4g1
F28houoc2giwTM/EEwyV/MHDmkfLh5mVyyxdl67mWxOXJiDkyIKuAB0jC2Vt9yIIqrKSyXaOnjwm
eKg1v4lTwcWQehUJI7azOHEsyjgIvfq0EgpYHmC1udyOhBIToLIlWAYe2slYmBsubwrX2cdkHmJJ
8wxKYAj1wuu1n+4pTTwtg2Yplz9YVAjcx2d28BOUP32MP4xivPOLXQzs27Y3dLZTysv0FVNt1rAb
xQXivtFlbl47trMaJ4QEpgng44XC1dhZfl3TRdvo4v9mGZUSuwAh2+Xc4k3l4rKBZDq7ntBu3633
wQg4VZB7XV2fxcdOEAA+Nu14bjQUV9MQe0Ln6klRFksu4gzH35DHp/OyYvIVu3pJ6Y4sDDN8EQs5
ASAnPd0R8BVp+BnFzSmSIp4aOwfinqcH4dWwkVVwEJsT7sP2ccGGBwmh24hldXhKDUluZbeQ5vaH
TwrC9K3vxVmmptdYjbR7QzU5N1x76uz1HZK4x8cwnFFl3F69/GLJoEfDtkAWUy5DT3E53UaUyAZA
vlPC07QpeuAsgMbE4KfCprVhh4gAQdf0l3Lwzi85HqQR0etKJN78x6/AsRFALC+EonZVQK5Ej86d
u3RqdKcEyJePmzhSK5/5ZweWL0J5CEbNMDopu7bEKDbAX2NYTorV3GuU7z7DkUZxd6Hu4+h75JnI
Zp9NNKVy5TOgOSYQqE7K3Tc4E9y5UDdHSySeZjqThq4hgBtlmC8Zpk4AgXUZwLDZ/kz7/kI1ZSYI
kpJvCrhqocWdBdgoYrLdL/l4BIlXfPRLPCfJAurJR7EtsVf7sD3wiLPxdlMRMzPUwjLmO1KI7Lkv
q126gX0IF8Hys0sB8xRF8pRYSGiF3oIK9v4tTUtej9TrQA78Pb6I4XY0JU21pbqjSxUOwZgy/zp8
BoW+AkEi/6wfDn96ylF4gFQASfypJ/WkJrF+tsSaYbulMRdF5z43mVBOiKFJUwwxYeal13uSfD43
1Q16XNSI9mcqMA0AHgA85HSYDOKsz1gIMce1/270XCuvodHm5yQkXgYTL/3qU40yWImn+hjT6kHx
vxGoOqBTfb7ykwbNGYQ30GmX3YTSdRnMAIOxZ/3yeQJ4sCB8YZuH+1Z/Dv9Ej/ZLxYdpewxvKjUO
RA62JuCCW4O5YYZs0A1kUsNh+nQJ6bLj3ODJUAKxc0Ry2r1JqqPj7sSzW1IeEPzetY9cgWh9n3xa
SMTaq+DXuWXKDkDysHsJP1H9sEYUq6HXmpqPEOy4fIJACXTI3cSnlGA0UilFMVXZ7wC8HFgNwHcK
VLcAMH+YIDDhQUttNZNswzpRDnHDAr22+p6hRme4zDFW6k8xOrVv8gBLIEAq7QuQb/zzsOOnSnn3
kYhRrQmvZkME3gvIr91KSJ/pJKrliGBSOzzOOkdshkLS8j89AI288xboggrO3td5F3r1SDGZC4Oo
Q6lHv7fEseVgXnUj99A1/I0EmEDVy9P/DFN36a7h7zYUdZ51NtCsptqH0xLDOlfQS3F8wyR0/hBf
qNNqi0sr+87aZN6enY6AGLxKMqrDPo/zUT1ORYwxG5ugi5XTdhMuGNyYbQIgnJDAdSWw/4rG+nmb
uM3njGzHMjFUcMpUaS+YvzQe2uCMAOXpQKfyrX9UcLj+I250ayisV2jqNF7eNe0UFD60t8BtGS42
eX3gIjQ9NUP3Ii6t+o7DjRbznM5kQhSn+QVhHy0Ca2vgrISgKiyow25dGPxtOy/gL+iJmoCdCjEe
l9N0YsXbqDfvHiySMCds4amFocKbrJDxk3kP3oQcognnDE7lG6AS4nwRX7ZxTnTddFXrAFejLBgH
ayQejfGd1Hf/35saMm5kBlrX/a3NQWPTtPqsoRkquaPg2R21k91JVbxurnoQEQTDrZcRl0Ce+ZPc
l9ZFTOgLMU0nmoal6AaDE4+xuHxI4hUYctGtHWBawSUaIxHVMgCw0Rxze8pHX5fLhXCj1E5ctGjk
VoyeUjTDC8iLuzeO5XEHibcxmGYHU0dZduSa9YWHL45gNeAYYpy6HOVzrUr+3M/19CwyxeeV7xVv
C2eNWDlJ5LY7Fg4Z2OjCGderOVRQ0FI38fEpMFcdk4rxPFa6bD03ejkJTxw1bCwRxE2WLt7+lG/Q
xL06ppHMxoTXanlSMO8MsH+l8Gd5LdAjuNOXR7paV1Qv7r/b1aCQ0Rj8WmULtcHE/maHBC4KxB42
FTUYgHrAV92ZaLxuuOGGxBZZSPm/JIBmF97/7jhr3e9DUjuIPZyjPqZNzfuqzmxORi+sZy3ojH+S
//y1XlsDM4xy3fl06BNvMpdb8oOfUbKIcqBnPfEVaASxytqsfJxnf53FVlWzcykkPnZTJvfF0ccs
C5SN1eBfd5PKhzikxblHfn8uH9eaThXt6cFPaAvFpH1VMLZoFgufKS8+nT5Ntec03qEp+gFJqLE6
kl+DXSHCZaBZF2F6mKJgINtXSxbIx/9GUxQkTzuDrwOevFfDjN/sWkYh/B3QmVISVe8r27i/Osil
rYbCj49u/gLh5dkm8WNDFseLQenkyAjbDXsSlq5b1YtoI02rfE1/o50YBVvMn9RiS55f06syXU/+
tg5xZkT9lrWTwql1eJZu87KiV3sYe/0i/AJ7pqsOmVQ8uLxB+wZbhWpFqg1bcxGTQZLGj/ORzZdH
FyMII3nkzRi84Irkm6cK1iI+t/jJ8o/cVNAdLZujNRetMEE+vYw4/Z9ILXrcf46bJ6EFR20/NdK9
H60/3X5BI2Pv6elTeZiWgn/0Ob7N+KDzTdFKvwrNP8AptVB5nMKe37I9nASmFhAC3oe/IGnl5svP
5gjla3Wj6g14v0UfuMA8/0STdPbG3D9cUI1B0/6RtxD3ftG6l46hei9a1WoGUesdDnR7nxOXBnXC
oK0BtI9RJrPD1pNatuhv7GGmYu/OKoLvnjT3soZgaq78NYgu7mxlIBeVAzozgYE4WT1yUWLEDWjU
w4rvwCXxg3tNXCotx/SMRAhvDLbsmSinl/5CfddpMpNbwZEkM9af66eCsc1ClTbH7K7Xp6RralFU
2IcVdX0VPNFtIea9tqRjlzCN2z5QnVr5xZI8DCbZcgDGV2dpf5pxvXdZTrjhjghanH7v/awZzVWk
4wal8WbUeeZDM7lHBr4XPoiObEIG763zKkIHpEHqjHAkmStI7tsyCn4XjphNiXrEPw+qEpc12qw9
N5uG9mnOR9/h+yEuiHmaiFFE/cQCpUotTDnqvF28kqhVIrrUH3mrtbUoC0V4sCbm/ioRGFAhQKNy
00KEh7WH1nBM2mJ8CM49S201FdJsTdKHD52z+btUfVYrXrYAS3O42Jii/Gw46RfX5m8l5GRvRQKI
Yzchfsp457GNBS6fwsG+TgLor5YZXN1boWpnIC9Vfn69zhr6ACgt3NjecEGRl1tgLzyH8PpIxC9q
WSA6LUyzMXTjKi0Et7hVH1zkHABDIiY3OQwAbPHNjSG9LKWCAlsN5OsyxWvfhQJ5J9b7MbsBFpH3
/Jbzam3t4STcnD7F6zH8FZklPe9iJxZzd0gSKui+gpn1Sr1h8MlNBpLbbahcyrsThU6fOax0JdwU
+bZIEGe/Ht0BTM+gfBFkSSdc9mbQjFRsEcIlWNffIoQTW4mT4/t/szJtudzDoPM3GzQpBJ8mcx6g
ZWf1esdJCpG3Fbm6po3vDTjdzJL+W08zV3oKKkVbaDe1Is+bKOOX5hVhwarl2Rp1ckxs7FWjZOS7
uQ6HI5sdLdEe4wMlZ7sRql42xB7oeSe4rMF5akSTqs81tHOIFMBvbaMWODdvNJbKzFuYngyhfOAp
mZ9N29shytz59hI37lQ5BEyEife7tzBsOTyp829HXg/yjcqglqP1YjkbFfHkt7cbGr7aRBGeSY+Z
U7+mXeb4MvJpjfYBDBl9sGMa7+3gbw54aknxfyBkrP+mNDXQEO7ughLlnbE1/C+9X4P3lQnNDrKv
vfS0ricU/fw6myPeFbq4hLTGf+doFvfYnaGYVe8tUwpI+tnNUJQPdfmcx7C0tModV7rs3NCB6e4t
nluXYvsPAc7UkOxC5j4k0JTeyDwUOSZ8ZCIy8R+QpnZN5rYcpCNh26/Xm1PZLK9GBn7tho9GAU27
8eO+szLW9o97bEce8nnIIpJqlZCXMguCX79E6KAM+QhYeF2r5qlSFsT7dNw4n22xf/FtYWrzeUDU
fqnkR1h1fJ+bt4PlCYzEuzKbTu6ZwEZ62yKjOpsPQ5cTT2xuKnhDdz9vEvL684WV6UcZygieUBMZ
kot9qBSRKwxOrq/WQSIOkER8roTvpmWYYWAG9PLdt/yDEjsPIH7a71n0M4rtbSN889AyGqU4h1qF
ayNznx70CmggynbGHt4SAKLRneSUvs62k6ZDoiE7tU/Sqi6m+hb4BYwByFuyXw7X3kh4hL9KLBOX
WVv2yk1o3zRVrsiL1FzNvQIIrYDtisBxkIXzjajWDmUYsZpzCeIqRRzbTBxk3+t3ItOpkGDFJaBy
+2BBnXrgkGftKPQ8u68p8cwADk4hCPPX9S8eyV+VVyom0Du1VWr9+MOdkjmc5R3SMbpGi5AhpTgS
4zj5APuACkJXQce9yRDsG0vnfw53Jxq3YvjJofL7y/UjoTPM74scL+J9znDGorEKV5UpN3X7Acju
GdWo7oSSDJlgwQCMqvWQ2pBfLclhK7vHxtb981uActYogq75LGU3CNQbK+9wJEWIEi2EXmlePHgI
dIb+yPtGCOfBrBF2W595Txte5IYkiHurxEH32DX4ivIKFJbj1mcYejZrIyTZMeSEk7XQsQMPGu48
EGRKrpnLgPRa1oBSSn1/pRnumYgwUZpVb8B3fqfJgPFcMlkoMb7YL/5iQyvBaS3QIoFxhqYFGw5M
Fim/9Wp/3cJ9MDY9yN75/3anSx+0eINX4UzWnzgo5JvxqiRhYMdSQJrxff2wN6jLk/5lU+N7e0vU
DjlJ9GCQB7uBQjRIemLj9dxVge41WNhejBHS+C2Ok1MiviD9eqiGYyiB+QirLsFgek62tLgklrhP
lgJLr1tMq6zFRWyXH5lMq2mDfMGvZjnuyn+AJjc2ZYeY/U+Hu62YuItVbg+32HJXERnUMoajGxpH
h+Lb7eAeaMCiktXaj8/Ya83vdahP5kivAY07BJjgYPCJmXf29MqpKdsb9gkBV2Xz4oY6WJj4fFJi
2kguTuW8AYgon6RyRFiNTP+uEyquEFPm0sTaT/ryerEpSb5/32eJdj6vXfBNfF1x/+jwlo2l3s9x
sgn6KiShLrvfgVRyteLMII51SDiTDVycriWupxeXAF8EOW9ATWtQan0MgJ3thPYj04kZIc5SroBg
T++9Svfsnh/vk/BUTkikOEy4L2Mvr6fC7K2NHXVCd0CXUS68WGW8Ah5OC9V1Tf0k+EYLMPLG1T44
t+ZYO99W6dregJBY0Qm+xlBVBJi8Yo1DTrOM9qIM4Fg1GAX7W2Zwawjgs9Og6p9rQFz1RVnMeoDu
bO+es0PcXEHYdDMVvX/HJtz8NzL4VwZeCdPydpkeO6GZNww/gHDuLRJO6PL529GF06c5vz0yKhAA
OYG3JJed9+bxrygAplZDCLY8C/5RpiC8jDnVx6nNcahNabgUd3fnIPHvXzdId3sdZjqIAvDo/z2q
oPBpPTCGjkD+Jjxs3vDdgcIkIWI2Kwaom0y/eifCm1iX36HUgD1yuKNSZ2nd8fS/9MBXPCoZFjyJ
6KAxMHmFspXhtvTDH7xaPCi8zL+NlXXUO1tzMitllaBXF17DPrBLtnp/wKXgIprHlgkhOjJRfzXp
D8ImALIbQ9jcWkGm8zLHK6WlMBT3vNgZb86uE18katcI4otAAcIEtpaRCg6S5Ky7TkjW4831fUIw
YBuearpJMMgB/iMIY2u6y2CZUvX6TP50OGj80wtHl2GDYqM2Ax4XHsNZsmZkSAdWBjEGSTMnNqGr
1ZGSeNX2v/0Nv5UvR4OEJgCZjfwYIKOejZ8aTVtktLAbC0F6LHMS220UG2uWbxu5IyRQeuUflYo2
FvdjMpiYIodKNQF2R5UyF1St2nfk5eK7B+qn7YKqBSzX//bcVtQL23gJhN9I7kpM8n65tCzdyN9S
9TAgjnjbXIqR2GX2Kfkch+oNWvfxxSyuZSJqNC6co2atSv587skhFpKDBm2I1ej43R91O7H6aoro
uBaKevdNS7vYy7sXj6t13piltxpDer69c29E8CM9J8eYS5mxftjxqRGD28AOiV67ZQt7XlG6jC2Y
UteVMy7VDZ+CAA3GxJ9BF5zXtoXYqdAudxoIpOiMCDZXaLBq8ytE9bkYGH1YBu5i6glrgTVsiW58
bt777898tz3CYZl2E3lPmyuztAEFWLzBp1pDc1NUYEo/KID18m3FnN1+9WX9IrbZi8iZ4fp4lM/q
xOkjZNvnt13LJaGk23nawxokAOBe/tu6BonS3m2hE4fKuy1ZzOSj00pcSHWj1iJZ6jz6TsZ4RQ75
30+MOSnBS27B7cfkOaKI4QzLIQoGscGdwq0ZqUZd8NEvxhUBiQeXYhrgYUnl0VQG3boseCKwMJoN
Ox7fNxu2Kh9a9E+AudA0vaGD41/g7YfLE1bujEIND10yuqVwv8ErK6/Cs3Gv4mCL3Y8aSjzOKXoL
6BQNymqWy4Dvlgp2pAhVSbGg65uC29AVWRAZ5+FsNRg8pZVE//JGgfyEBGcXxVrXCfmaYde5bTp8
NblItcrPFfaoTZguN6NI4F3TxOP8qkZXQ1hgT0w3uWgVI3KV1251jZL0XsboFVz5O7oRWzoqtvv/
9VBqbVHbNJvofSZB7VSHkjQXJ8DoEQMAVzTvPbBY1LRv23xsrG0o3xdAzA80LsqJZwEblG4DdjQL
mvqR04No4WVngAvtL2x/m945ErUAe9p+oWfloDa/x3KYvlQIQIvPpbXVTgq4ZMRZmHrZ2YEvkJzk
o7WeiULFSGNZadoO/lgg36Rw02pYJDPieVIK5ki3RQKvl++UnQk3B8pkj/On26hSCYt1kjY8K96c
noSRJjRVkHwEZ7j5OtqmvNz+9H8qH0OKJlRMH6VnPm7U0lp+cI9mePOwNM9DzCzowAyDV7ccFdHZ
eg6EaI+at32UexG4qe05KgRY7r8F4E2uHySShjm8IT5b4KpCHd6gmr/3GCERPHeHRwPggj1alD4b
HVXkfw/9xt/UHximdAFDMXx2F8rvEZE5aCn2YCLL/oUqOOQ/gaZIp/3EDAKVhhivTowfXMZac8TS
a9woueQDBJeyabPWUgOOGxMkgWlCpMEGzbaBdxtjxf2y89YW/8mpGRDJp5bAM/UlaSoFBWYndYBz
5D0aE4PLReJ0B9msb3w8cJmwRwwKHW/JISHxR8MP0FRjizBcxfYJcg/txLV1526BrPTKK0JfhH2P
P9Do328z4eDf8q1eKGAwdRJkt8Y0jWPoolvsQEmgypao7HXZwL3xIwbngZfIW+KTOatXH1orfekr
QxvxNFRfwNiRgdxtJYD1cvWvCCXGBocDlF54O6dEZi2WFoL2FVXsgjb7fJ8ZojDNkIjBdDtbFfro
eA+CaMhDFCWDl8YwAbZKwjvn6EeToVvQlBxNawEeH7gr77J+J3DjwaR4l2ksummPKR2LByn6DEND
eFRo9O+MbfOUUtnKJ0Rp9tNionAEaPCkYzRT15CFSbL0iZJ4HEQ14L+BSSjel7CUcmJzONFfpo9Z
cYdD3TzBW8327vQ8Mu1etf0xYS2G+mkp0EK9oUz0Zgz2YuMIHUJ0RR19QRfFA7WXJAVnPEP09lSm
BSGf8oLfUzX2wsZj33dzWmUlFZ1xh0Us6z3te0YS2+XHK9ICsoKR+zndHzFFk0257Ov9bCQJURZ0
Az7It3HChgJbf2pqy2EPunOy1JcLhv65zRQy+HB42Ny1UppEjW/RE8N3Z1zOeaxzaWPsLTA6AMBP
YyXVD0ROEFicHZgrHB9RHC3DQZn5qgV7Q+sejcXuHbUjp/Ta1h6aa3JaquWifbcg+aG9IbGBr340
omJABorN3fy3Rf5zwkPyBGw8vUHajgY29/luga0wG4Y3fql6Eid0AhZTjFlRh15twDSkrTgxDttK
WGs/r4jIQn5DN25fp03RKcPvBvkGPOZXcOK6fONDG7aHcrkhw4XEzswU9w8WVpkWLNXJLdRhhsj/
3qA9qsSwXaY42eqomSn4iieW9POsXomwdw05ozIjBixfqTpfEeTnmMgop4fcyOJ4XU0CacsOqPok
FFKqgiyD6zfyrRyBUVu7AHeoe4R0Zek0s4bPjZjIX9y3ehkkEFsJA7NTUPJNprQqf1SfKObTgIBO
9Vi3Wb+Bo23dufFUc5qO3H8mD5T+1eWGvAcS3sV3Y1HvNYVrSolw8kRUmxybj/N8AtY7VFWPEDjj
LG8qRKTgMA6m8UpMS6vDDB4eES7mBZSerm+rMlPZzDOZc2z5R3vjUREY+NzavhJlGFzWREKd7MNI
EHYpr9Fitz3IMkmFFfmZMfbSkvfPpVGLuFV0OXpQ5/TczjUfwTW4VY3a9m2oSENx6cAYUgQwtNlE
r4gOJSwwXC7YrEMywJTgTrHn7abdmoDU4GTDygZOVXvq4a/HHZa5S6iNp+XMWMjZT4Vc5lMoBOv/
T5taNFFejK887oxm78NuSqd4Iv2zwK2ZXTuhHVOsKMPjht7elQIf0tJVSyI/nsR+75oop4wqXmxL
hcDDhY9NUvvWEcP6nerc1B7HB3JPQYkGjigVVd+vtGshs/gZPu7+wE/oVNnSH4Q5H6VkI3/mq2Qm
lLnmMCtWUPlxFMhhjbJkSd+RFtz8G8Endc8sjfcetkZG4kjqDgbAnXRTY6MjmyX+KcbAtZDe5D1D
eTg8lSrAuc7WqAecCkHHhD5oFkwVxrF+Y9/uBUU5REP/R72vA/BPb7KoYuYn/nkXjhPskRy4J77r
+we2VZKsDqPwBxAX2xildktmdW+LXDa8h+NPI7UMelKnIc444p6+1wYBhpHR7T6iVSjKeEMbr39L
OfYjex/0SWQMcc/5sH0rMWHr6CpDxVR36RQPOI4bj6ND7vTeDU4lTtMeheMJVBGfgzoUUb2DqGv+
SGN5MXPRM8LCdX+ivph+Dp3TWGlNhWngg0Ycl3gZi5M2bpqLzUpWNqeOr5RAF0DA7B6jsVrqglxk
pU57jjnxKmahjXKdYk+k8goUQ6k/inl0rDrdf5ReiflWJ69WZxBgq1uJ2wPJQTP0WuEcd4FRyjmD
Iwy3Rq9hUZ4SnfVIvmkFU6kyhONBeVUCEkkaF44UoioTIv6IMrXLnoEW2eHS72mTW7vrHfuEmbx+
RuM9sHOOTuUkksx4KhdaLZud9IZyIIIerAih3u53jdZ+g0BUBm/ts5EH7GI439WTXNamqsuvVKM8
m/B66QLA2sAnavedGnGutvxzTVU4XgqrV8Y9drB4zDG+mnH10gE2Tpw6PORdTfe1B2cv0WXabe06
QLYFl9nK7ToMjl7l1YdDzWaJVj5SCGnj71kX/Fa4cJSxajWuqrAZ2tDEkyrjmiNYHqoJMdMht75J
JUN9RIiIndQdiJtl1FnK0AIOvg5SHyDqsLH+KMMOICzrbILYr7pJY7Cczq5weqsbWJ6eek4Oh6Mi
bP2F+IAWpdd5JyInPlY3LSieaEnWZ3RsCAbvXGl3Vk+u9Z0DWtEghhlOr4G2J5PsLB2UlVOz7AEF
VpU2XiocwoGJ++gFKevJmUyYVRF6GNjeLGTGb/AjR2KUaW1OFAdZ0b8f4DZO6Bw7kXeE/Lk6eHzZ
upK+zlStAiji8hu0ZxWxYw0rLM3Us1yDeueEyAplhjLaOYV0PNRd6sQrVtAEZLP+Ws/gGMwSrgCv
qo3N3yK8OJYPNKLgiqAY2ns0eIQyHJYqEWUuORCYYyHa//U+vlOp0Rapk/3ckLvUKK8kSxhi3HAV
LOVtFXxqjy8YlN/TqcVyTHeTRHfe0LY+XmgG9dk+LyuOiMHZ6K7lrDuyEBVS/MHMR4MXmEUgFxIv
iVOuMZStOENYYfY8iS36yby4TpHRkgLsAb97csxI5m1xKg5w9tXOD2CCyMpaioXX4Z7OkmR2dadX
oFudnlHsHNPgZiGskXPFdhSG7CNOAk0kdOtnxQmUltNk3kP3ZVj3X7dubWM6BBuqiqg40tEJFQeH
mJG1ritXEu5gz5cbepXTq48Sl2nWRGkxVBFF7UqZ9syt3PgT7V1zF3wppJ6pTC5v7/xCKfK04QGV
purVB+sw+2cdIyPMEeXYhuPtTBUDi8tjoRmR/egGmY/eIClGi4xpZDm9zpfWMeuR4+61PD202KUg
ALNH2NqiA0g9QRoC/HUnGNP5UPr00WqSkrJraa+6Z2DrFtCHvk0h9HYe0v8ZOdzQ5yzO1/qxm5Rw
rwZnphOtSywMtiW0PTOwnD9nfzObQC8Eq/390woqCxVZoyxjob6ACvJ0Nqg2HpoC5eIQdLJ1ol01
b9UO5dnM9h/d48uUTsI5smjkZykMW5FRrggK66Vhf1HXNDAGW0/xy/0enV0RB+qCQADNZDmMMhNo
lZ41mAkdbZsuWhI2Gijm3BZQYL+xHwOIWdSVDCdHuTGkawf10tp5+rlTdg80nTJa8VrpZyL/aEr2
+6/qWTNmrTR87FkqIAbMBijwtdcP89Qs8Bwnuj6BkBJX85hkeNXHz8qklS3PwRNP0dspcKod1B1V
pUVNgWi+iy9uPzKs79dKpfWdA81P9MqBQaoCiKZDUrOTCUoCY3XoKpxfo/va02SzTIvNxhmiCf3s
kkmFzZvgDHbFwvSaVC7JrZrxcXPyqyk+AcQvcexPLYmc4vX2aZuK/E3JUS7IOWl15gwbNqSlybR6
7fSJxcHqT7IlgZwZRheeMROHU53pbMu5HIS3xUNerwp1zxn6Ll/SCTghyp7M2gd3NScDY8b7RHzH
56VRCI1JoxiJjj03RRa/6l7WY4rb4bOABrdo3dje7tRILjdFacee2fnQL0mhnoySL5a35ZF7jU4S
3srzgrUVQGjh/bNtrsqrS4HLH9SEQkVm2EQiJmsQXd0R6jIXGAr42ugEtxN5evLVdsFzMTrXZHI+
+zYln0xMzx9Z/ngCiwagDCf0WeakmbZfWMiJaDIApLdWcOi/QNzW054lGZoJ+ENvIqOiIo85r4my
jWFlAfmkYq2BTnk5AAa0Ly6SPlPI9J4tUrJui6AGwiOKvc0kiXpzycOaM7Vo8B45awqR6JGYG6Xq
2PojP2Jiru48yhwsR8LNLBfACpa3p5dyLA2olI684VgzkDxJ8K5n95keWlOyVNqM2ChKfqoxZlG+
fC0tuCL4l/gt+oZ4vUr8R2zOsR3mxm9V4gZAjJMN6NgDjfbwGDwcrGW7RWMNthyXRLQz0NuZ7kl2
hteIQrF4sZ2naDWknAHtjJzDfo3xE+jE0K2kf5Nz8SftR79xAAS8RADWYNAKHq+0JgC4IYL7+lHp
74XXUx1Uv1uPV7M1CGf3TlNvoi5naCk/1nn1g1mxoy9+TIqu20tY4lUk5groDO6O34tAwYC16Hsq
Iin55oQJqLShHivkRGBYpK2ubtU7TPnGrkwvtZ6aVYFnAQY8BQ5BiYHnxs/uBzg/NrsGo7JFEc7p
jZcaS69FmN+wEVBPJzf6753XLDfFYmQnGv4E6BG/x7sx0XmXtoFeQ6+WSGg7VOvU54HrMxCi3mKX
8USNPzj2A9Fl0DsB9eFrPzML0hqP2ycD27+Y/Ebyfo4KyC2qiQMZOdlhwu67VwApI9339CrY1A1g
bEl0KvIiDuUuFPlM5+Bk4IAI9Xa/lfSrX6feqaoclW++EE6FC2rYhMbupDKQVOqEPbiuANaKFaXY
mEIwDNFpkngoWCIKECJYFu9LZFKs9eQblTvcB7AnTL4+k0n4aCHpYUankcl7Tg69eyen4f5ZIoes
Z0Jph7IVMn11O+tUGGSRVWH/dcJRY/UwiWSMWgsXEDYxS1bsncfKRKz4TiqSPMeUXB89dH7gYkgJ
jGlNolmk1UGQgdafzi27sUAnj6mDl0Q2vtA2Py/23I1bDjUcK7l/vIPS9gZvGkCjeG9ig5HFuQm9
eRXM7kbdWO+yLntSNNDGHVAc8Lw/Etgbv819oSg6GfpYsvE+fSW0jG4r7LHqZac1OVxKnF6FTy4k
I5Yh/+G2FuIJjrHJbSx4SiUsUp6i+dS9G5cz+cuKKxILKx/OLT1Iv0bo0Biz0rVebm+z6lDzXN8m
K5haS1Cmwz1twAREwijZA8dnkmpYuMKt3ip6AGBKbblEQ8nquj2dbly11QHV2zYo0CVuafjWkfdC
eJ846vwGakBDRyBHOTNHnv07jY8ThpwymKrbZkUJCv421MoHvnbKiknQz8cjEzIU3x//L4I/FUI2
2MXjrT11F3+BrFpWArxl8G1sm0ERiDVd7jcoP6QoXCBn7jZzWISQMzt/vnnYAShg/aM7Yo2/3keF
XVVGwoQieUn9nQ+i8gjnWsqKVUM8RgIn2TluZhjxmAraWrd40Mg52WLkujWqHOXDCiVbQWyOpiAi
858N3aS4T6vm3X51tTSag3CFviTaBPOs60rnmQITHeXh/c8/n6qdsUUE5IOCrFy85lRs+Unlcwql
ZGTe0QcTWvE1p0aVLls0KjfxPc9DZS2cI8MtyCI3g2UQQ2Nvz/yZOMIGV0tInOFK9b/q6uWLmQOB
xT006JWnoqiv9JivXlc8nnwCTPiUIdWhhZUwDgCcuI4DbPkY7XL/hXzp0Vphr61BfPP2htflJin/
/MYE2OgU8XdrG6wq70t9VgxavSHfvRsqGraPWX6x3xm/QeLWRl9DazEQGhdjPkleOA3n4tu7CN9m
dZ8pJFL26QE8va4rBOuLjPEuirYIi7U+OzF/Sa0qOj08XMhBccbglSPPod8fCcCp6UcrB+I959y5
SHjz5VlyNJrnItYfic8vlSRBXUah0PdgdBZJlf73XxWScV0+Y7uOV5VZZZmrVWylmUSxrKL3ihZ0
jMQYmllolZvl6N6YzlOcuXTP490fswF3niEQfTRpPcckdZJ6ydZpCg6Ts5AxUp74KRDPXQE+J7C0
m9mzGoVeOB878LJPd1R4V+1/RzPVm7tMun/eEqPHI/Jq5X0Pix2YYlJO1DVcMHKMNAfP6T6ZGzhT
asQz/mshJ/bPl1H4MwJ2mO9/Uy6FbgX/umFFR+xmdZcLWVkS+pNVgLHTtwL63G8I7bnTipziRFy9
qKO3bmpoM5SaUftYZ1B63rMAsbtiCLSdUIjOHQPjB3ovqjEu6Fy1j+vWvmpVp7mtKbWLURiWRIBq
JRPur5JD0LNBFnPtnuPO0C6t7uN2YB0XbHBMCfNydA8LN188gW2vi++bqxrCkiQVe+gQ//fPFLM3
13xlRGHTq1HQmkhTaHL3hBOVBXDmuotp1oIu8q5h8zg5lj4AN6PIECbvZOkkm8hYpyVm6Wxs+UpV
D7vBUq9h+O8lARpGSCAkRZQIN5S+tcwHx3LDrqBoONMmAmEo7GeG1ZAiy2e8KEbBCCYYjSXQ+NyZ
KpQLbVdGikZ6C9Ddb9ZISg+yDiw/1OF7VnlZlFZxOOQJDhW1slp+0qFNYBL3YkJzQLgr25Y4Vg3m
RRLeQpEdVafXFUqOSwujZXh22hvLFjTBiQece9v0dbcjb8sjAzk5sVvVCHic1CW35/ZtE1SeaUv9
s9/zgvpHfgZzupqy98j5Jb4UqkkozSePYW6bPqF85aHp78yX2qmA8oJiFfCTT1Bnrn6iP3WqRFjA
HRsUSbS9cZw3gtt+KbEpIGl9zfRFCkMrUZvX/WE/R2BQrzXi2ZDmah9mCtgeqz5SJKCIk+BmaOhE
sSv/Vw1tnSEgcRJEsqkGJ/UXHOvXMCzTl90Z+COIe2uHBPVpAaWOMDW9l/eBX9xn3U8trXZ/8LIp
GXz7FwlSrFjnhHuAA0AwW/wcqUOKEe6888LR9KFDh7Ha0DMLTY49qQhAe45iNlqutvyAWfNghB9d
+7A9arLwOOE6XLa/Z61Kp5cWaBHztIsnxkATk/S985H1EXxBR7vUOMhWXa1gCfr8Z1Q4GnXXZ0cR
RAGI8/8OlD/2ECoNOcgSdb5R+Iyq8hm/ECHDn/ocj13AxDYdg1l+bUYUgRcz/VPWhJmYXYM9woVs
+SFqjfcvhp5gk9m+HCAnGnkCTsvY0GGMPjOd/rYjGlD5xYvglghx5Vf/N2kgusBkHtlpzoD4Uv3D
mh2Mt+dXCV3pp1t9QUMJySZPsXurXw2jxIPvivvJ6M0+82zDxdvx+EE8eM/BwED4B+EmeX/cLEOJ
1+MdPuWnA1bS8BIGgyZjRHcLb+p0EbA5iwZzO3M8e5Nk8xesgocwbGcbFQYc9jnqxqo6ieibGRS9
A+5f7uLOoQPLRk8jROQg4tgQezsDiR6QsCJyW3Z038UThfeFQHysjvwqY5tbl8dbiYxG2s0Y6ZM0
UZKDYj100pIdMQ+S18C8n+P2ewpF6dWvcQhqkH3iqEM+Q4jtJgHqPdQXNaWi/1+8okXO/5Lw9RYJ
JCoBqpyzt/s9AmOAMNFCngcYsAuiZulF4VTwbzLJdL68+UxwpdcgGbBza8WAbE929k7C8crPuJgz
ax5iOxuA6KvSqZG2RCdU2XT61W5VfLP3Ej5NEnaEXNCmyHj8ToAc2QygWmXz/nye58NucaklPTDx
oM2E6NykxXxvlLfls5PQsk5V1dGiIosVahcMSJNdbT0G9gIZlBigIUmzCaHXNPe6QvYaD6SOFIfD
6Hu3kLborfJVNL5y+OYnsFQvI3qY+88Ko6g7Qi7pRLXm9ljtEkf6sD5Qu30tydCO7XxBD2VJncy/
Wtsx4HpSL8tQTXAku3Jr/DJ9ulnEIS2qarF4DWJ81OmQaYyG9wZu9pmMNEqx9nzBK5WrSEGUDnl2
eW3UAvJ3UBuFP8NClsx0vG4YafCyVajI/BDoe8DSc2Tc8UCA20zWrKys4FYchoTAjPMy3HyrslR0
fh+PKQGUoq2uBSGaDGi/Xh5dM+t9fx3IjY+oH6t+jmydKskWEs+lMdnyU6QAOsLfof5tEYZu7h/z
+LbpTM3n0EmbDz+Tc845yFrH6r2rAhRhYIZ9+bHKYq2zhJmjqDGNbkpLsHQFPBQvvEvHCej5Klbp
JbDDzBP3DUya/BJ46bbe9X+VSOQMz0jXaDlds1+DLmeG0/Ud/KnX6pYIfWXeV1OTxnpAP6P6QOOP
kX8fOtbD7nPnMJxBC7NLCj3vMqI9ZpaNgVYs74qY2HCcAOjf5gw2/k0+9GOx6ln4Ko7SGsc6Av2G
lC2vWr8R3itC4Pcl2Fq+ZnFBKvH+ug8SABvGYlawSxHyVc698+LGKCHTSy0pjMnnHP43VW/6upzX
VnaiIKFk9VT7R/LHrxq7AMt05E+njgJWcbeN517WZY4X+U78R4veDbhlhkWp9kpaqrNVIFE9BItB
+3NnbQjqqkzgIEATJHaQEcEnP8H4RDNE5qmbhcZY5DdJAyzqGBbEUwJxaIT6szgiUu1PpQ4m22IZ
IA2yEZLLzlF8/Pb1tBD6Yfp4jkZRVMwOZG9aMz2CRijQA1+yDnQ96Yygi3hU/j75LWPBBtTHtseZ
3Ykt1JInJuDArBTeCKksyWqUb5yolz00BoYkp0WksSz11I3jEHjRpnJO1x/TE10jQ8F8+20XTY4y
w4S3tEZYm7TCuIABJsaZOXDoWYVIDdUUN5O7A3B0PgoQuctUr0E/4HxDH4kIpxirAtu7s/3u0oAD
GxC7+WEfotH8qiHXsoRN19dFIeru6paICqcMBfEVq0c8HkxhFtfe/j87OEXpqt8ONcotT/RBQC79
fEenacdzJ4w5OBZKwi6L+N7QrLoUzNbjLZri5LyqKNceMt7QoL+2ogkDuzqLHCsCTTmcxucpxAxB
TXBSemFePLychbFJ92CrUt9SNP5KWIE+s3lCYFQ2CFFCoREOPytMeOdn2ubQIMMt2SnqqZmYTzGe
fsDv8G0CK1AEhYuEgp9w7cPwi68Z6Sj7WJPIbzPfWZ4HIomnPfNvl96IJxVnXG+LzD+Z1lIKnrxZ
AzwmU0aIbRGsnCKYASyXaCKIUbR1Jbe+1poSPSVi2p7vvT1GvOh+cQdCdtnXbK8pc89Et0hZy6AT
OWNUBStu5IPEskT4e+CKaok1ouS9j8HHFIAjDsOuO1zSJZDeJ7HUm8/+fuJ22AvSPuGmHVbeOhgN
qsC3q5SSmLn8aYh3eeeMmyFWwwEGIHZ5FLGBmD6Uf5BrRTurjghi8lHHTLPmb8vXbH6qR8DhyiEq
Px+Yto/cJ5fKAmybWbPz1jdf+lZctspki9pEK7IYyCQJFv+5nTEZjwgZfC24hJdvXtOLxjUGLnwz
pRR9/49V81aTdgLXKJy2GfqaODiaB06XTZSyzJ0BRSd4T9Iiwnqp3diYu3VnklhQQxzYxPROEEDk
Hj1aQ8WYb2Xl/mX19K1cj1iWU4IAnGTY3rhoDJRD7nrKiNtWlnceij0O9814QbxV/PTZokI5zt4I
6pNVy/+Q8uGwV8XyabyYACN+iGz7URt4/wKa8o/ZrfmfeQ6TVYnjG9jpFN1SGmpQ+CoNjXHMU+FS
/lmKd3CWbDH3Gs7G/9TH5n9tG4UWtSWKd9w6izU2VJuXTdYd8tVWTLA/+Mao1zYwZMMsC3RFimz1
zX8DkKPp/t7WnOL6KA0pJDRwPnRUFs6AsJJBPS235eg/DqlYQXb/9m95+fjlMf7AFT3UkQIMgYow
w/TsYv12uG86d8a2x99mDNhGzSv2IM+PhrKT9dIS8Ro3mvq3Hs2eN2+oA2ULg/FemWQR+4WoMm7V
8YlD0px/u+U/Mwz09bid2X3nwfnfa0fYA9vZlQGvLBvmdtgUb9o0by+dWmEidqhHTo8WhpKq9o0f
/YaXQrfs/x51xK4tY8F7I1UCG0O4ar0NgHkMCR4BJPvLpexc3oJq6wGClhj3exCmPLf+mYkRD2gs
DTVqa91ye+lex4QBmc3PrjWf+oBURJ40m5AiMm48dED2hhaSea2kBO6QCYaSDTz3HVDcItXpB0JA
RuboFimjyQd0aicFyM6od4YrAQ0t130uhJlMEw3d9GY9dbi3LS73o7c8C4jIp5RVer/4WAtTqZLF
Z+6D1zeEdhytrIBwVLHx3goyRISRIqYg9hoLVv36gY9otbDRylMNObNL3S4bekRux7FHD0H5mIda
FRzgpg2Z7vKteCEBO4x9Jo9A17FsfO6NtVXKeHQZramHddmsHTglv9jhSyBAc0EozP2wpRRdRhRD
/pkLQc5GuYyUFlq+Ztmh4RXEAKrt9iuCJLsakh3ifiZu849n8yk3sTsnkUXSxfIZrGQN4xaOVatd
lOUPbEFe6KHVBhcDaFHKATHHZ1f4/KwEWgkWyTuX5hDBm8U4FrhFUnFxNgGcSQkpvGhAnF6oiRet
iFYW0rjEgl3j4iAIS9qg0B4fhCfvVQ8++j9ScvKKir5iUZ0GahL+/lkLG3T1rjB/P2/Z5TCYyabH
SPC1CLO0XyaS2zUJYD/9FozpBd9iLSmgxKM5+LSC/b9KO0/87voR5fI7pEZyT8wjc19tC32mAyYX
7wzFOZaF0AMQRLy0wAgjO51gmrdoEQhM6wBnSqxFfoUZfjuCoW8mlr/qGfFkNXK64oULMO/2EFAK
jU1NKcs/0FN4prCJkpgO+jeLYm0Aou7L8ZbddtNROPUuserVeVaeqgyiWEFwxWRWKQNlOtlHRKr3
RzNCFwHNqgy+/czMCN6Hzfvo2TTIhogfxOAtQNa2YfXuzUfnj0h0iYPXXflRtTkaRKvaxl9RPcta
kKeIXhc930Hub/Qh1XhwIWr2mETbrrZLT43RaCDwJyY3WRQbYw7Zc62vdYogz8KhZEyxny19IAXb
xPiG2//oNbrz6Jthgq4IIbPpO+JKYQGE2wV4Ur7dLyhtHRdxLSMCEmn2/ic8xZuwr1r9pHZbzw+x
X3ddR60m2uyfsyzNNGCj3aYAMr2l+AVpBioucukajCLfTLM6KF5EC/CUfGKNpqiT8MY54CR9SCAf
1rd1jliuAR4npJwdx34lJBYmhf9P6dFA/ei6ENXaqRwAF7Lw4IjGMwqZ9OE82fbkl/KeHgwLmCm1
DTvcSWdZol/4Poak8hTNspzFZEPrWG0zefQSiw2taExAbunBZnYjpf3lsh/htpErL2dmigkmTAl8
wgw26VOnmq6hYv4Stjx56gvH4YGkEg1CBWjXT0F6knajlbM7mETUd8OALgoYBxMFFpvifeUxY4oc
3ACJSxJxaETo/l4bcA/0KZ3sGPRbHE4XCR2ZqVayc6drG9hRVYlwHszzKqQPZbIKX9DNMhtp9sre
JypiAM4Gt8JfwVk7Y9CxSN1DLAWiFQopfYa4IIZqwS3zR4doZXYkauRS0bVOMpoT6aSu1mtpVRGG
a3OiRSz0pvJjO7lv09SNBYWhgvKNfzgoYmx1VXdd1Z82HX+N4mDAcYBZn43twSJWAhwL3xl1q0eB
RxANgX6UEJIe7y4r+GN5BpHld+T8e5M7/erRLGaHLI3Jb175Bqp6RyLj/Qmr4f8mRGpJ9DOvlUeb
txi2ylWos7KVbv3dEceZbo5Tpn8j6Psv72mmt52/1SPA7KKjKGY40s2eiw2hYGPs/Z3NaOCq1OCe
f10NaJ07qM7+CTiRUq3DHa1KXxehcjaXZ+TY41Q/Xqy08PmHlAzSbI8tZddJAuKc/t7MYxqV4SC5
f7P21gqC73uXAFgAx2s63qZsjbIFDrBe0pJwg1r4ueufTWdonDwL65iBQpS/+LSgX8FLvyCDEdcK
8ZbY+uCyH4WKgmDsBNQoM9zK30ZiECOBfdSN5qnv8LAv+twgbrfEstTG34mVUqm8bsDY0C+RSR28
fRo7XBpzUV1ZCBZbfLcYNaUUrzzPBGM5bzY/upIwx+IexTL1Uu4zsjtjAPP/j4UqPTolgws8+xRE
Q6M11M8qa4xEJF4Yt196RFU9sIycxOcAO/kOuC+VD9IwNdDctxhN8aE59Q8mYNUQsh0xJgSeEttz
B0Lyr+52gsC9yfVKQPGZtIdLe4sdEV+IZxJ3pCRK+Zh3Ct6yZ1XybDgejuOCzAi+cAA/+l7AXTCE
GHozHKrIs5wepmqXXWSS87GW5PZR+8oqRYmSYhXzCiFco1tc2yzjtMFdn426Ps3zzwW2mtbxGET8
SuWRh+PvbiMNBzyG40qnWDu6khUGSZcH5WRkLjE8iNyXakeXB2F/4sly++Y9j+VjrtMqB18Sf9L4
1FRxZ10j5yzh5uTzqBM9fOLsZ0E7LPoH7lxzKWbmDsy4HYqW5/rkmmYXM95fgjv4b2Jl2/samgY3
+UdzKUScYXJSJUO0il/s4HqnwoA57q+8t0Zz+3U/VDILmflKQ3slZswNP3LYHKtAKBi0Az1OFBTD
WQCJxY9oFJ4uGtRLuXq0IWabLDLO+ZRc1j7JZbKIySMa4MSnNHWHB6VOYwKAkLsZpHLTg5nqrrrX
L0AQPs6gkjE27+JgEgx4iIxr0mPCJBlhujip0fzYF08bs0DwOWpHn/zB3bUse/RLIC9iYLka/GSM
KwthBIeR+XZx6M+5yrgzfRLwauamSC239u6j+VXbg95h4X5KV84q/IV2SsEuevCKQl9pg3K+UH6L
VzsJajsCbjVVnxeLASi9Z3zq1Qspv9HIp63QSa96jV+6Jf0BOECSuqoE6fyTHstSgirwyV4utD1f
8pVA1FTp/G12eu7Vr+Va+lR6JRsvBJoWK0gIt+apKo1ii7F1Bl5RCXGjgde57+c5KkaToYIIoacE
0DDy6m4IJfbIZyQn757ZtpSrDI/tWchkhi62muRLEvWVcKI8TZMxvfMxP7cm4osvYoIJ7S/nvf5g
zH61dCs8yexwkwbaokbH68O8eY3VC1yjSseUy+wn04snONpNw6IOgkJdUTM+NhFwPlb4IPpbMt94
4ZYGXW8vFRl6xGfbO6gfgwJVs+Qs5m1vo/AcZpMy1KT9D/ugRx5rc+oF7vGlhhYcBsxFjtxbQEu5
OjCWE3L8ivWNN/AunsUGKTD0aw5snqQ27O3xNLbRK25sdnbnMDLs89bVT4scLN8G12rjhC6eVbve
flxmmjdRgQTlrLxvoWhuECmIEKiNsp7ww5egcnb/cijITeJCjMaCuuqXFAmXCDi+q8lNqeZcqOmK
uXie2isbdui2bT7Gn4fp+rwlLnkMpBgKqvxCR4KYIZsOrEJajLu7omaitvl7HVNy0NdOVWvtb6/M
oIj2K/k6TNAaqIz9b+++uHmAEaSnQMfSawpsCZybP+lGgRO0CxN8Apl2lNXZXl2n3DHZO1c7PKRU
dKZi1iNIJ8rJdrcfQPAYcMmLxxcRqLO5uEFhp4r91vH8y5r4PSd0Kbyr2NKw9X890MnPg87dEjko
cuvKFQV5DOT4cCLeDFStX2eFjMCGgQap8u8lgT56nq3biSZENnWBU5uNSo7mfR+oBz3SIt9gwxAC
PxO7n/CIxdwFnKRpOX65Vw6gH8oo1T5XOB4vdJO0Rzoc5DuQjANNzEHWJXJPf3319f6rsQy9sdYo
2hjosfkKnRo38x7PdePggs9GV+w6BiJ7x7EE/fhDVL/J5IXgsRs/QDNmxSsteVUJWcSChdhZEi+1
y4AeuomNvUlj/0I4226qFryQEWHoiv4Ko3WleO5MXV4dFhZSf0s2Zze/k05r1D23DLwH9o8cT4Xf
gs+asMsMYKJ2rbcBQL6RmMdmIglIX7Ekv+uPa4GnF3vi4n9qbcMRsCaGwZHeg/141j+yx29xU7fg
2Kprt9d4FCANWMKrcvb64a64ZGSmtSodRUcng3z3bOQ6yAG7a7SXpIn58ho3KADGjgEw8F95jcvk
22Mnv9/Z20QKkJghcXRkzzuXozejK1aFlpCUxh1S6iBM7jjtkL7B+uYCh9cyzZL2d9W9dn2q06Hd
WegnioVgg/HiPFAkBxQQuQZ2VTjYZwDUm03p8uDWFheB9NJ5Z9dntwKuEbvAJH5+b4mr8z+nQpIr
azxNDlPpLKmTo6J7vXWpjbfXETMLjPTGg7H+2VC01V9XX5uFDZAJxlRFQHZNxuDxKuokDWLtv/al
hg9Y1BP5/KqEEZEC+fJAtq6V+EZh8ld0iRVJtGcQTmQ3JfyzWXaw+TdS+dw4uwMk1I0CSaZSxHAx
N9tSFkKE4La5TcUfwWamWuukCfFBNqVgIzEjl4r2xhQaI5DHegzOS794+18/GwVDLrMCXFZE6f6f
ZyCYFffn5PGQl1KGLdfqab/VLSPmoK2VAKvVTyR+tY8bbGx6ThpbQDYT+zaXzIyUPuFXXvj5mDwR
fTU8WwSJdg8jrmTtWLjZojIZ/QyYIE5cvihCCe2gZ0SoeMJdBeCfW+p/QGaQ2xyMe9qBgBNV1jqU
84tnEjc/DiD8ZkdYVUsktzJAOrAeZkhocOAWdOv/3rXyluCFG3VzW9Gxi3Isz11mLtaoePdkqNeV
LUdEmIQJle9R2HPzNyc490Bkw+wcacnjLSW1cr724TAWsi4/OyyZmEWIiV+3WD8xoT6C7y6kVBMy
L1fo1Kdb4+/soCVrGwGdODALtI4Y3H6I0KKEW1ZmxxPqGfG1eXgA0o7B0CJP7pYq5BRHZ+sFiExc
Z+eIuvzUHK2fFXr87Am//66lJt9RTO5BnDWYfhu886t0tC6FndZlaqzc8dL/bOtwuPmOrP+VLVUj
rmhgHF9YiNVbxVWVLjVTvvgoRVpramWopI3suJ/7Zx8WFFmnXewvppTwzZtcdn98ZBNfKt5Jvioa
Jy4XHIezf6MKKl2aJAN4t2MxEHQ4kuDt2XZVfH/6rftuLfQp44jnZO6/N5Y5vlSWC0LDzm3cO12o
7ZGHuKrWULo/BnbFVilw0sYKsb1gpa5+3Su7Nv0UZ1Zx2yIKIfEaXT1LNCJitJGYKtKJDZcA85cs
LxsdZDyRG2Wao2MQnYSo1Dg2Q893qho5aKK/HkQEf5TcyGRHeY1I4H/h2ug6Ou1wv6U1RLgISeGU
V7jFHih+S+MweH45Fik9u21Uoog8+kLVJewdoNhuu5QDvfMvcEjgR7yAvFXozL27XDg0lZE3WXYG
X78omXPaCKvEHIMe1IgyGUPNnMqmbh7hEArM0ekanxlqnB1B00Py0OsX6OOdWn1EOX2Z8KLoyNPz
HRItPXpM01KeXOp2wqrgRX4I0CpY79TAMnu2Wfps2YvS3aHk1xlpOK5ZmRAZ1IyCb1G+O5k0ABrA
REnbEZFNxkO7g5TysLcOxmk9e2ua42i66GJAUgXUSF/QfImmR1u/jocyWxYYVHgoMBQxPCYqcdIF
iuUEHln8Tlkmq0zp+R50p6ptAFz4CX93AJeUwgleQNYvadV5crvi54Jokk1gdU2Ro3/eXkBuYr1x
iFkrH34sAOddlM7Goo+NYSQI5DveXjxk3mn2vhVQyj9rD3sto2B7ecV3Q653SzJOpCWddF/GhgPi
SLDljdVR0aFT066/pbboPOfLPseTxvvPRwQn7SxnjF5pgJnVI01FNReBSk0xyp7Afdvu2sn8KqpV
WB+EF2tRE+XdIxTcGkoVtpVJvKI8U/wwuFRgVuT1l2pCjT27frN3FxuP2mq7JzxGMkrA8/vwzNqg
BGNBpg0CocvTGlNjdMZn3gbV960NjA6w+yV6ZeWVOTeRpVIhaUcBPRTA8BaKh4X9Blo1tInnZemp
yuzCeYUMRKKcTzSgjS5+jbiovaBxYTeN9dgh851LK2QmF50nz1A2RNLVnmiZarulCt0VwJWGynA3
vNS7El99tSK26+RSao0RUvo5nLmCLy7KF2yBTPRV+yxA2KzNbKitQOSGh+Xg5QENPUjgsiHw78k5
rlIdKqvDDct+AZGMH9tLwaV3AkgZsCYl5/GUPBY11inMjgPrU5A2c35cTXeCrZmRQrU3SI28ojOU
H3gAIF6PZJV54isd19Y0Bra7XLGJ3MR6lc3V8BbjmuynDTfsPFdOiPppSSEY7/jhua3LaG8RcrVs
8Ro3mDdUavyVC7b+x/uLh/LNU9uRKYjgvGVY/24sqwIJi6BYdYyD5gmNGe+yInmjPwaq5Y0onaPd
wKqBBhb0H1ABiPaiww1HBeCmdtShh6snjrGDr5FURrGATS/nlFn/smNS200pQUcPiUw4xGM1pUH3
eAKWt5grWNcKWqIlcso6YhuPMKLrG7Bi7MUSfVR1A9V29lN1LQZvGx/Ds1YJOjyLcw9N2qcHIu6j
dhEsLPn8iZSnrR8IkxdW3w1xijt8TSEzd7Boevu0RsZwl2YGPvAkn/4XzI/501KIUc44XCQ1SZDj
tlLEigp3C2ea5yjfEYLj+a/tUrry7pNy9XBIks2XUlpqDG/4TvN/Kzb7R9Zs01vf/0jfquoIxOws
LR5hzyyKcNfPYUEQbzVUaVWWViuMPjgsj2ZSHFBNi2JUnyCu2MuEZqRJ/p74mesbhuCqzisW8kF/
SAkn9ioMkUWi2mW0CbbNa9pjPBSwQJnpQGgBLF34s5sxhH9/COZbQHL01lURkICXGhJoxQ//J85d
KwsSGHItQLiqN2+eFo2xM1+kAK2cgyv7B15OxSiZSHF5fK5ktLOv8Gmc7LAoqNIz2zuE6wbxoTAo
wFIiuiGBScO2Q1q1oPWK811lMcrIOQpDDea0lYKwe1BJ4m9EgTNeAq0NW9JZMqj9OO6cYsArkwIo
eagjoJ+pninwK9qgX9+brRrDuJUfVDLZoCh1bQHdPex8Muv0xLx+of1SkvOfoTqc5tbTdRO6Xsbl
gH6GE8rH0bkUZpB1b/eC6Psa2KVxq+l3oOZYXQAuXtjPHYZdbFuK7uDnWNkiglXogfFyAIFH9zLw
ileIakjj/74a8rWRgGre+y6zc61AtgDFCziuEgxd+2ABPOVqiBZyGG0nupvS2Bt/I2SZGGggW4Ku
hjxQ+YDwDCLLmieWMkHoGertTJYKleZt6PjZVkVVeo5ITxgHhQaZKcBx92j3I8RdKQOtT8No+jUP
/hPvgk1irk1zoI34Z7NfcTufqGL+frvOhYQCVa2B1s9vHV0FTZzRI0Osao0HGXxU+/RjTCjduJo9
QxvLdAqE+jQkeC8qBQeNj0mI5C8Gbv/W+aAtS+87YQQ8vXrcCHycJC4BIVnPR6Qd4qy0oRFhIwE3
i8f8MKHjtiPxqc3T47RWv704e4IEdiSXUZ0ZsKB4npQPn+ias1s1Zp0FdN723//+EZ2T3+SYpcTC
rH9h952k5h3f1CS67b5SlT93OwglFVPkXv/eEEUKhbovDS6JFBGy00uzs9br8+Vs534K4Xcg3lmk
n1PZ8ODWcWarleuBWUHwcqjEKHKQOSLj0V1wGGxCV4pGRqgIeaVBl+Ir5llcVjQ/FZiAexIWMjhj
Ce7/qGW772j6ZotgSiY5kxvhW3qX7b1aXKymH7H4zA+qLCnOAhW0fNMoLGj6dpMOTnCLi/ap3uBV
i5AgZtL9r7nCDOoRWKmJTcJJKekU8I6IY15wTeaXL/NGTyxCno5IHtw4K5rlecnPfRxy2RRBs58J
PtU9hnYFO0SOhSIpEKYk9sazp97OkJlKIkD6JYBUaUhK04HIvVfCsJgnuL7WsUkGDo331sUrMAZR
IMbWRMND/5I2nxOC2nSsQLp87rnXK4MrRNWo11F52oV1tjlRZBrFdC6ex24gBGpOv8vdgB17tO3+
gvH4Som4aVWVepGHsO4mPTe48AXLr+e78LoW1DTRM0IVPaWbNKQH4rn+dYClFRpj4yb9332eqmIW
PrTP21ZcJs0wBiio6CwAI3DSzXlFq2HCVEkngX8XxS33Uz0tCo6k4NaLZEcujJyAFMWHTrmzHI2z
o32EGbtv77hr5szc8J6coxvYAgtBTHwLFvJApSHclFru6NivgE2z8XIcq1TJ5QNz9+pmBCPVyuPJ
J+1aHaWlsV2X8TgsGdvXlSWO8iAK+nLI0UaMlyjAC1l7D2LbqQPSXM6lTPTsiKG94LkbvZErJWgA
LYsuML9CJXC0UTMSckQsBeuV9VveIBV3HoT7TwsyxR43H4SjlHAv4wo/QHVksSjqn0k2uG9Ne6K+
fN0ysOwgh0h3H+QSH/yZhZC97SI7kICTw3aTSAAAjCbp4ebtRy3buzy+iAi47YauwQYqIX2LieI7
Ot6sGGPqeaNWVSDnFsLKxxVZkFHtw+Y2vEr2/JrmMV8UOSej5qmRu0Zu7rMs1C0RETZqGSn5WrcG
NkgJExG7YAxHb9UUFPfiSJkPSCwhCKN4eYOTz7LAEnaOqgRNSqNc6R3Zwn6llZ1ufXAS7Qn/Oh36
SsrF+t7VlwCtjsJ1m1hZmvvk/3T+N+ZceMm5utA8aKGh6kcyr4BoglUmuKVgwgoumxQprYL1tMv4
psWYDK8AO/asR9si5nOCF4PKcEf+2HEhM0m6bk3SL+MXlL39icGik9MTq6HVEd2x2F+xgZlQJy+r
6QHWext1DyE9VqAG1zOnnZBWGbmdkdptYCE0yIPnR8QLGS8awuDATQlcbWVZvSZIy0BnkPIvUi+9
fQo/gtK+zmbfjTItD4jvbAYH30gLZ39DJng96YwA3s+1lS4kIhU1tPg+rcK0/7J8HjwNr1huB/HV
R+AHgHuWsYzEjdv7Kmo/9QqHENXOcrjzHLzPM94SxPPvldJawy5g+ggsgWvHBckRcQ6iZzPbu2y8
xMr9n9KN63NjBo3BPluQp0ZlgrAoll3XP25Y5848/zvy6v6KqAUE9NRjRYsjX0y6pMB69Wxa8e4J
UMf0d7sO9EMES3nq+XuIzhaPjObuYi4bFWyYO0yGRtCwZWjb9hPPk7gT+3IOlZACFUchxDPyfnh+
gNkAk5XJ4F3XxOu+m8B6SWOyuMR0w2lpu9wH3qBKRsZjyemUnzaBtCY75vIg+6bTXv/cvvukPP8P
NVsylEomPzY/J0Lvcb/oJPpRmbGyyoaRqkj7w/RTox6zCsbFfIW37zEDE5nbOTeZKpBaJKdgPjFd
Oe7Y22q50803AD2WrIapmFitweHaRA516yHrdLuQG4uIm0pG1LzF6Tzl8O6Ch5181imxQzTc1k8h
9J7yhf1y2UIYiRoZ78Q4lTvk+W5H9kIrSloyudTBZ/0nW4AMQsaXgp2hq3VKJxfhbxZsB4ml5xJ0
8Prm3FYdswEh/Fd5K+1TsKBEVTvCWRbI3qhXIny2xP2X0grQazfSEqcfpEZc+XVmr1EOAdErA8r5
YAUyBUD5Y/mw2SaDNdFrLdE+pgvyYNDZH09hP2tnwUXdyJMEBus4Snif7vNNFor3UcQBa4Udju4F
19yx82jY77G7+3buYqEGD03qs4XWANFcwUBxrdYSO7vrdWGp9inIjUImfwkKi6Z18lN/jFwHXV+4
Cwhziccc9TW0GRdgVvZSCW+QhITzZ2Nm7U+AaXC3AHcPRlw50Civ6IXQJr+UPXanrV4p6p+cXcYd
oll2xPCMFcsoEbIqt9ZoMxq6Y1oVX/sHntMBec3/LcA8IpD8h1rAuZUjGWRpE9bOksAb4v6xe9KM
1waCASi6lhVKb0/JoofOoSHlGlC5xeQAljrU5XpQ4meUBpM7ZHmUDx9Sasq4tOvMO/m2GcGDt3NM
fluGnUNaePQ4LrJI/oWJBgk2zEn5vR0gcsly+e6FjXx4bCrKENGg9/fCfqogxn1PpdpbnGKzd2eX
244+m/cjp+fLyAVOUT73WJk+h/MnZ9hWexf9vSs3YuQ8BRKtsFn2+p0tdAQ4XYnbhQj/+XVy5Rlq
cuFBCk+jM7gEwxbZmmw+tnOSYPD9Ka1gYkjIA3461V4otK7tAUtH+J9FWOKKlFFFd4Sho8gKPVXo
MF5pwHlKnh22xtEPE9BfCz1lOh+iOoDyiQPLFtzorAtfHNnSen2p7BwckcbjGfkkwDS6QzyXzDoe
kPeQ4eW7B1zWDbymSQ4osQE37BQGwlAPM3hd+wxu5iqHmSFH8/bEVDunWnuru5p1ePDIiF/KZfjR
YXLZBB1aDOZWCFPr3F2I2Sc2ZdC76YZD69KHTrL3rd925kI4vifZ5PfTJ43UAp3SX+vFVE8ptd6C
W4blSDKGzdeuWYX1+IygnfvDxh/CHaoST464ovE8NaD3nJ5XdugzJmmi/0CX6KYzoyK7csjzyiRf
7mrz3lBY+NjKzr3w67nH2L6bhrEw439AiSXh4/QEDhl1EzsLP8UB2maAAxLfpnSTyalfhxRJp5O/
CJhi8VjibjPsi3yjwYOSpPOR3ahLzxZPRynZX6vHQdWTz0e6+Z/ZZ8hbaukddzOm+zWX9jiH/P4g
1BSlC7HbY7MxvTnOl38mQehkr0DWhp+Z0e/iN7kS7d84qojB+KngbJioxgCr9rtPznt8CpIJyOQB
tjbQ80yhkrD+jMj1WuyexLdHV1OioLngwp3W2LVz0Gvrff2HnJy3tclOlWiRFi4SZkr7lNOqrSbd
thobqnrANhessItjfDSkfhtgvnh6yumUd5UHHpO4g7nIbmp5SSUwG+GSVAchYE6LbnYdxGGskOla
i0NJQwzYw7YHYH9J+5XupJjF+VAVEiiiT011SYA13FSiT/D8RHD1zKV06m2MYph+Y75itkGNvehN
jyjZoKXzDdZyD1t7OLSXahiXLf+fDwmLEffrj6FtjrwMYwu+s9JsjW2588TrhCYlntFJmUOX5f+N
7d6MHZ4cg6eeBkexZd1aftQ+mV+/2uKEknP0mxVXCL3VKqHB/c/b1V9Rzu11E2mNywNPb6yid8+O
v6/rDu5rrdX/ZsdlXsh53kSGABWGyf9prKu08lQe8Ek4PgPjXLCs/t9nYLFoDeuDMdEMUh7ytiZE
dZMBOJn5i+2mIyea6IGj7vMR7xL0Jpe0oJyCpiD90THRpmG0eUO8cZNsn5BvEd9P0AdLU43bIwNH
X3WO40Mcsi1KoB9NoSvZUTx72QsTrwR3yCupQPwxhzNXcfhMWRFR3Eg/Qm5Ew4rEZhFs3lZ9G+SL
GkU+68/T+LR4hvqgZoINvKurlq9mBXSvrb8qOhLjyFw3/PLfEsGJKDg3TvYwK5GPqPdO3xNzaopl
eCKthEwC7n2DMiiRmEr2aOZnMHRCp5APDsB67HaFTs1FTVK9BDSa0Zv0F7bc1kMqTtO2fkAdWCjN
zAVYS0IVPtAq0EOMB7ejfmuDRI5bLHTwfzCYWEMmW9WqKgNHf1/2Vfiuhw5ow23SIlHxBmZa2nJ+
bG2vq6tEU8bo9U50rAZWRaYw2osup0cLBcjWwdPe3fsVU3I1K7I34sS2fDshn+IFFd2CE0rK46Yo
jubIqLow4RU2GxQxCB9lJPV8ZlCeNCF5OT4WVIJSGQ2myft7OLO1+BPyMuAM0CCBTx5T1dVs/M1/
L22IEAR8ABTY2IiT9YgfltBTBnCXjRYaQ5XeDghFet4xgJXjIRj8sn/QhQB4SM/Y0w2C7HMmq9Gg
/NE+wgdnTNvFG9qu6ARTdoRo+4TQf3k3+jLKKzzI8M3+vLweAbKjjRvqrjv1Ug2+pO1QHaQhqCyU
zlz4NIxA92kHjPI7NSzFMnibrjYmlcpXFbW71b/ec7l5TXUQd8WeFXgeUUfOTQBGJn40lW5Al8oh
s9CMzpwYpJpBfa6tWrUkNJsTDKUuwO1t43gfVRHUnUJfAZGsX0v49P0apYT7G9Isd2SV5IxSPfMu
R0IaSHHSf8WkbI0DiQdpcrBjckwN8mEMqR/Xnxa4940PmOpRiOXFQHTWGK4f3c1NSGvscm0WVN7+
O9IjIM61+ZXMYUemm4UmRL4/UGG/oCIvQMV5jLk2zBSiT2rODobciroSMl1kScPleEm5FsEcQx/8
PuKmNMDR9qKh9IKnM9sVu1rymvR1X12c185l3esJg2FpS2iAVNlqLaqu5r+X8ACCrwy0BS9zYRnI
nFONP7R/v+jlCx2rb1TRkfQgICXQL5CyXTlrbyI6ae7NGlFBj+hlYZIC0G5Ar3Ie3Qw6B4T/DyFj
HPQbb7DJHIeeqkvkrfUdGCo/1qBi8rht3R8kCpH0raTEwuV8qwUK87t6NfFwQ6w28h5G+LWBp59k
VS7R+64l8keV0xgsDCVAZwNi9b618TJqmTmFzJyXE8l/MQWUXOboEIGKdMBsUqgnp5y+54WkzZyj
l+xnsg3YT5LiVtXi8uubYPNuv8u08iA0wriYDzNaZZPoYrOPdyEz4FG/DyD8wSI6Iywnt+uzmbtU
fDDY8VRizDTFxlFNo4ICoNVjGeol44IL2VG+sKUFaP1YnPZDaI0CM3T4jPDl+j5mzZXaezNGFdc0
ZifnjcIDuqgAwq/uUNccgoEGmdi/yLMjOLJQky+xdmVc5jBeatj5mmsG2+8+mDQhZA6yK7Y/Nce3
O/cE3cP/8kyP6Fe1bD3NbJUQHHk087ywKaUHc7ok+u4pdG8W6rNr9OHTtIj5zsqznCgKqJgApYCE
xlllnUnpLIydtwPoc4MiLi7dw4dy7ew8C14GKn3NKFJKj9UGLV45OCXuQxROipd6OsmzuuXYYsGO
0W6VJPAjhYOs44bfruknyuGaGHErW/55FMBuL4EeZRlYPq+4xmOvZemneXghtLg+JFLlLtbEvIR1
tyb54QvpSXSGtyOjFXXvNT/Y8JkFgauoWqb35xdDvNGFIYWBHHG/hygpz+qLMru3/GjZDf8dNOTQ
7MzNG+LU/Pl9LH+Xfl64lQbAYxAT+hHzuPod1JVcRswdVsW7cCeh5z3L6L3H7d6fca6S1DwUr28+
+aAxO+s8DibEwtB3j2neBdszsukaJgYoaqD7QfoJURJDu40OQZHSillZSbTnaanQQKFFbXgGDWkf
AW7Q1+EIxR1A9BPJX8D1wbmL48HfJROmmW3QGR3PuzCMEn99pbs4eB83+n8nMiZcfqVUL3LVyJe0
qy/LDPc0/fqLT0SC+sDZVenvWSePArt/LMt0vGmF3rildKkBSEGMuBkYAdZ4XHiacu9aT8PDVUf0
pvXevFsfCQbXZcNaFHY5mq6y23a6/JRyg9MiUdTcmzw2GYh/aZMopauwpKmnx1dRBtmBAoO40QNU
vEuYk+1ihDiNvppUH9ZLKH/qC4lbf0PlvMcSrhLdtyc7H5VWLuD8KY3+k1PYLc2+aanYmTEI3Twf
iLlASw3YqeP1KLNOs9wAC/MgrVcRL4Wq8cHtHGxM7DBOoWL7MIMMENjMW+nBUSAXcC/UG+BoHD6S
jA6GlncsDzUBcUC/UFrE3wDVr1Z6RdLbUXytTXakHwo+Sl8oDl9ZbSSwESy+idkX0Za9gMBLStRJ
1jenAJPRPulEuwjFKiRQ3yD+RQSHEQnZ8e1Schpdy2iz35NsYqBOm5KKbMazGu0CNRHI3XGMqUv+
NTAlmbCSsq/RkSfUUrHKevX44fQKsf6V/q17vkCfqqRETTfTtnnFt+7SB8NF1FCGqISkTAszplIe
tpPVxUnWQP8XUf69z1GOdf/OwyB2oHZS3+t10Nu5uf+im0BHQisczjriXosaGTy67BamsLZj3PYV
ndgFzSoGhQECRyVMtGHS6bIDUdBCNzfLF8QfCrWg1e5LvdHnKkH9Qc+5ym0uaSH5QTO44TI8NYvz
Adei+/QcSAQ2owe+z7jpey/urZ7CFGkFGEvAJlJusD+ZHw3iDWpQ9TEPrjfWm7sqCwYEYQwCK+1f
HmMbRRiD3b01MxT74Sk69xeShtkUeRxtlQW2Z8Xg1pPtiPjq6T3UC3y4jzqvkZYgK3TMZWjxpvOP
vgQHv0egqfgDWZV/XOxNydbmg1earkHtdHEz0kpsSDjSlz9adNyxkOzYQdoIMDTY1lpaWLQwKR/6
ukLF6oAnZehHv84kdG+fo31eJ2fnyOrYa38IIMUmCAgi8CCSZqNtErZjgV/DEFwzLwyY9HsfnUpe
4wuI81G2D2uAY3JH1QiCHVnKP0Z9SD5/BxkxP4daryX2yz/QDLQduauRvJ17+Qf1d89LRYwnTMvN
GewI8pZYDclS0iWhw8YJYRJJ9KqFYTGrNi/t3SGgFGz8t18COeG0tIs5vvN8FC/XH9ke9ho11NfE
h2F+9P66f+Slj3vEb44Y5KXfPFM0LWy3IJR5qyV0JkBLWiLDufFSAH2Rh0+zdNMSlxAq3u8khdZq
eCS14s4LmBBRd8AJjtrFkLuybPyVO4enZXuUpafsApCHd4wvTfElITPmEPTXQ0rXmObhgy+YfesM
+LHlHI4Kv10AvegZxmLotlHkySmsYuad1UKvPnga79BKwng8Z7gv1F559vNnxUiRqLtMw2cHgjnJ
5c5bThnWj81DnR2b/sajsEgo8gJyNo4Q8PAqLR5BbvBue1ByhnlU98KXN9OBE4QT4e7Esha4WUnm
hCJ9zF9W9qr80D6ZGN3WJg2bUyaT5ZRMHpSCWbPyi3v/COPHu810BUMplgAz24DjeAfeqaPk1RjS
VXoJH7CWi9wriKOuCFMWPBuE8IkpjrOIH8WlLV8Pz1lmVtGDflccWdCdVAkc8yeyt4c5NCXCGxh1
BZK9K+C8PVEzDF+ab5dciQFjK0pOJI392JHMdYgdApGhOPA1HlkeU5wRS7eRgiPmD5zAYo2AlXIs
2O241n27+HGvHOoFRoAdsOyR7BcWyQgZFSyJs93ngH4yRDjoLg1jzeIb5/XAHkssMV/hUh9r95KB
iCYpC+uNl4GWXbbjmrDxdeBGZNKlk28kEppJ1fIhwFl/ZyynATakinwtUjUWyZPGTOP/ncRD4MXR
B1kg2qNzEulgMKVRRlYGzsc274szbHumCj25HralGHQ5FAK4B5srxqG/SHoGaDsZhdNfBozvm+np
u6DuU8D6F8rhQgUD13/GCnui1XV3qrGWgB16Mg5Oom0n2OaQHvGH1ZswXbZ8Q4IkK5soAkYQw+6q
Ra4J+7++0AQWfdA9cqQtmBLt2E1w4cFpLuEBKqasvmx9aR+Vcum0CQLTuyBdzrXxZ5hsEmkKcf8n
s3BGx77U0aEV1it1AIp7GVIJSHC5giLUqXNmbRJWveQ8T4KCKmtIO6JzkQVNgL8yc2JGY4EDe0SX
3IK8/s8nBcU7JfKtZFycXtlf0w/TTd1tvNYw53eWACg7veE/KCnHbCbbumDQulp9T23RTH42ztb4
IAJ1Dp8352eIrF5KFEHSCKSdP8rJcJMZ0XlGvB243KW4EfADqeQSe6aqZWupQ8MZjg1omzKUhGtU
7xAFvQXJRP/WxnK+8Un1+W3AaT7ewYQtJHbqBRJmrYDcos1k66yEiVuHWeHRo3iPi0k6eWx/i2Bd
T0SINjvKWHxZ3e2X9Ga3QasZBpFlzDeuw6UpnJrqFztWvzra2NS3eZKKvQAOusyvHHXxKbSGX8GF
t4XtsYtq5/zItRXIrADzHreetQVPYYc3hx4HQDZ/b0zXjX5nrmz1AtQESV8EWxG12ez4sly2qvOR
gExXBlet3MHLKoORuO6/69eoCoVYP5dV6Q2xO9JxIxLw+dWooKdY7bmWOWU6URbFlT8ONMRu3fPm
vPChyf7Mymz0rxdLboGToGapvNKBNoit1BwV0GQD70RjTr1wUeBbbIXhZ/dkkYUfUiQWDE/kKl1b
Rr/5akIgwaRdJR/TK5rJIOL3wJt20AJGE4b1wJHO4ZznLtUgT2eRSDd/Wzft3SCGkWgEKYicpumS
CzjMRbEAJRglS8v1Y7SZ0jEuOcdicQe4HtEynDOzMR70/hlKytNeHn9tIsSuaZDZa/mHMc9Xt3eh
vq9CQPPbvq0ktmcJfbbwtRCiUKBxvoFgdjW/9a26onAX5pfuMbyzgrOxWz3mi9keRcNIzURJW0c/
S+FNrwA6l5P860D7VR8bsYjBVMHrQY7YQI0w0L4CAi5m3BSe5/9GUV685glKsJ9y8UuYr6tvq9+t
83mS5flCx0MJfHHUsgWdIP71yHyj7bFwRk1wIki3cmcaWm/0KIPy/MPjqE5kuag6HakODfGiAENI
s1WvXFI5z6oPs7WPXCFX3EOcLhh1BdeDVrK/tv011ExzcfvjqeMl0wCzeteljFkeEXrz/LCFDN0l
GJgPFC30HNJjnM/wGEdv5qXvjd82ZcX4lKLzUrN/UuFAtRCnquMuslDmiCgywn12VatcH1cJS8oD
i+cYPlB75/N6JTkX36L3h1hHzdj0dcIhRggN5lJ0XVAhr7mx7t/unTHJc09LShi8VtIp8GjIy6We
bT8wgGFZMtmGyvmZJBgieKMyx8BkSaml/HUjcwZ9U65DMUg7PurxxbVgKFeTippxD5CUp3q7FeOz
vRbht3+3yGS9HDya4UqNPFbHJI9R5DQ3wANdzN74xFPFr2iQBQ0MuWKUDqC468Y6KBdSPC6cynu6
zCeV0rrThtJ1LKgxy+BaXzCG8bPZWO9sxhFHOaa1HZ2YXFgX1DZNoGZ3FONA3oM2cY23sqab3k/1
IiW53000wTmO5NLLRNDJ8Q7VRs0DyE18m6KZsRVp1ewmr9yShC4ksapI/z0gldb4Os6ccmkoSiVp
LxBerDbNMlp6pAWQEb2955gNCJQAQFJdr14HUTi75hAVYgX+5yi0+j89WBZpVrqZF8Q9MSu9bGsq
vRpyhIj6EE/Ww/QnKrSm7QBKcCSuPhuQpVZlugUEj18LvVIi/qt7ojxELON7uDaUsxHe7iwbnqdY
tz5IcHjJnD1xag4gZPgYH/WLVb8E/rCU+o2/iRhHiq8lwXSwUFabj2qsB3rdN063R1AkeWaku56m
lrzUoL6VbOiZdfqvgP2rqqFLED1lPpAQOTT0oSZkcHGFM7Pd+I6AnlLRTaEYmNSjAOCL/f8FMwez
8Qz+kESxfVROHpoN8uBNJcg81oYbHExdI1zyEL06nLusyyzpKWxea7P2FsL+lV7jgrsrUqbRFTTC
9XDzNOrbPsSlFA5K775IEhiasa+wv2H6iN8KAYtV2tJCrCDT5cPxa/lymh1a4xpHEKYRK5nf9iYR
xBZQq7erDVzIjX1XfBzxbob2vKk2cm/cUJtZApTKN4kU0N4CQwTWqWASHaP/C5jDwv6pf2m8r6Zo
y79+Zx/5+VZ4AMU7IOLsgtJj0buip9A1k69iCXkgrPLyYxqNoMMidkMimaLOrCCRZqAYpYak7PqY
59I/fCseu+bBYz1uZ88f0sgiWvAXuVQOjtYk50ZUa+ry+nR+Ex3IZyaSu5k8MLaO0xEvOYNybNTA
3gr1C/076nmRXdzhjwqoh5Kt5P6CRR1CjfbuZR5PoR9rzr9h/N1/tn9VWaMZd6S28t1/x245aBZf
goRJ1TaI8UW3lih87hmRNk6LQ4j7oLyhl+bbr/cUVo/oZkvFOw/umO4P8b1rR8NrGaiM/00lsnrK
zuYZn9frf18ZP51hPp+pZ/T+dQdPekmvx/4md8phjB6s/6eZPaxliAMkWmu3uqnCC9Y/cvwPcJn3
vmKnXHMX3lNPLxrXCXMVuFzikscNhHgUU3A582wRyU9OVZou8v5eq80NYE/bU90u7jzxC5QVo0x3
5nFryHzl7F7mkgXrJyh6/0TEUFXvxtjboOrlNCx8SlYz2z2i5Tvp3nyuU2qtTZ3aFRIoGdjJiERN
r4HGW3Wjww9Ct2YFjmKI4+qpcGP5xiL55lfeX5ItXBke0OzqobU/606hdXs5yCSedGVLcjMz9vop
ccFuutjKgoa+RF6hIVK3e36QmBeWlwqsHDcVTua6WfPe2Pqd86BCfS6QAGH2Xa/LfToQCak8Bj23
BbnAhR+rs3cDSQfqToMDTjgHaxIyke7SiSWTYe5Z/Kl/lifgj0WrEshlv8nyXtL3/vgcsrS2NULr
YtZH6yL3x38gywVHsi3wzHU0/N8Nz6jdRaeY/lyKJAaTFWmk6Ijk+/PH/86JBfekNLEXjmP8mhTH
PuWoKbhLd7/LGDVbwtQbQ2a0BpWFMP0RElEzPINvTy617Y/zgh3jc9Pn0lhHeXPNYKUuxEY/M/x9
2vj1gM/tVq7PeciDw4XLF2ToaCg2Nme90nAgvSeWR01k6ptIs3KZgSBBaofisdPt8uGjBPO+TRT6
PAWSLK4L6G7/gs89wqTW3YRTt0wG6nl/BbWp4Vp6dMCnl53Hj6tCVoirLzZ8MSo63g/U9tgF7YYk
okU8yhrF0I7+ub0dSdGpXTGqhF0rfOzHwMS0tFTTDBEjxkuAGYArLpG6IX8iU/ORvMD/11XM/s+5
XDQWucOnHpv5bdS0EgKuLqH3WmuRJrL97RgDV/hJe/GplJVgzrpYUZz680nFsyJPS//EV+Smy7Ke
toFIPqT5wjfQMDn5lc9qV6VXYW6OjhXAXIFTZcB14TTSiXbyDUdoUcYXtOqSA7BE3UMjt8TafD6Y
U0V4GbePYu0rmcmGHhcwWafGkddVrbxtbryU5+XtdL7snTStwVrxGjMLysAyfQ647uPW1r4hgQKA
L2ZxfNHrYx1AMNWw4y6zojdHc7leDKMv8vk14VAmWU/p++/hTlmJseZpphanxvJplOOnTMmztRHT
5a1B7Pcu/x/BhOsVckJIIMYDlYRViM8p20hdDY9eHZ99sFffZ6Nt5O2JVyAZg7tyAkvO23DWNSsI
hIAN+ZTKfdCiH0NUUf3wELn/iLluMI1YegIMGrzWh8t8jBvPT7wBeDbiHrJ0oKPEYomms9fvHRTs
E2H7UaRevaiLlUJ+NkL8gKLbrdHOSyXQCUyt3ga23tVAMWoWz8wbOoMkAaftW50vo/ECOG03e9A2
jw4iFC7gA6BhA6Cj/ZuKqnvTWgF7/bkHVzKrDMgE0iYXk2NC/dRjwoLitF6dE25xtJNx+USiMvb1
dh0+PTbmEvs3qdc9D0kJbhxr6956ZnuQiNRwoobc+yTaZhpyQPpcZTbY6EqPmc6CinQaEP+cQTmq
LIqK+Vqp7qVhMp1fgpN4QXEbFXydUseQpA5kgkGii/eY+Z00BteFkMyh0ruIsFzHQNAgKCoulB+a
z089N9wso1VtAy6uUc8QgFzVtnPB1b58flgPy0OqtLmlr23WF9gdT9FErBjhtSRv3sBux/NbaTSf
vMwYlWl0jP/l/74Xqbmr0VHD/ECVs+9vEDgZn95AUStiwpIV+jSTSps4tXo1UJ+NIzjgVzsRXP7X
qaRAOviyoRCkrSR0IpaefvVjhhPYx1Ry/eJL3eFvDzBeFf8fVzSCXYtc0F+lfl7h0DejO30J7+nT
aBu0uymT76NjCIIpLeV3EU63zXHPz1BbFyN/DpGFy6f17ho/zUniKV/IjDRlXQTAbXNwBd5JOOq6
GOjuWL0B5xynn8/U04EnjUL5r3a0NeGzqIYjXJIyOX/H5fQ3RdaGe5KXBGMjlYrLABOwru8Q7E32
Q9tXmCSJ06rEx4pCCZA1mK0iNE7kFJyHc04eE9v1MyimHIVaB0BjYvrrcgjz5+pYutWP2zOlCyUW
41CSeCE8wUSTDBELh8UEE4cJncWTveruJr26kFmvorHH6JX42kN2ZXsEFtNvL3+gMzQ3HkdTQsBH
MViJbKunYF+s9TCbjVW9WsnQnl/4W5QRORqF3n2TlY3Ep39jmooi3mruIFS/jWY9tIiUfL8USPJZ
55LA8NOYGwDrK0raVBRhZBlW/PtXzliiiy95EWHa8/k9ulfUL6OJtLyqAZD6K48MRfMS2GhzzpNz
Jv05FM6kJSNZfiRfpAJDCmq/VpWSZ3kt9bs4I1tZrrj2BVTP5+Pz4FKMy5iIk6ej3BioX4hESZZU
LdDzYHPYqAp1axvWbUqKSuAkuSQhUIfQrK4yCqzgYXo6kPG1THKZd4FqTlC/H2UeiFD8ODJtT+9J
4SNMLUYY5In2QoD2V2MobsXXh+/lsoVkYEUBn3DWwd5TrrbNwHMyddcA/2rRVtGMRutlhL1bV3aS
fl2mKqvbTIaSpHN4NccRtUzahtBEQS1MzOXAMst5BCNhN30yR4RELkpa7W2BLwbFzbljPVhXhXRo
d4oeRvwT5zUyiExaP/gPN6u+Ic/x33xjyr/Yq5FUqg2HqeAUTYA/esfPFqiRSqn6Zpfj/xS2X7uF
moPeEhHqoiFBsNXBUJbY6Qx4TJAIl95l7EXv3eZv6+tUNyqnLl8f8PEhHOdqL2Hatj0BFmoN5UsI
TFNf19+eLpNmn27XMTEOdxhD+AIy2tx7CveTua4OsQvmFWRjSG6Xpzg+OmmxAhYFusxSnbnpwp+R
T/VO/PEdxuQtW12a8SngWK8g44U+n8dtK3nciDubwi+/Gs6vE22/Jo8ILPC21vkY6s/MFnvbqU6C
KqHGfCodn79mlOv8i+/NNbrJM9S58l6rRmlEOI4jZQNBR92sIUkeUL1JygIkV+9QdzwKtmK9wC0d
mizV9CNMnn7O619httCNBPxQ2SIePMikTYBmm1o8VFjm25RmJ6ihY6MVswTzLtZG40ezB/cljx3B
K+Tc41r9GwKOqds44MJCM8oQfrzR5WyxFNkyP5Esp260F9kBD1LJAY5ZEaqVOwCXDnmtX2+x+TWo
UgMxioaV9RT33HCJv6JaitCbPvyrHsvqUjC7ZPGPNNts1cVZbBXcm6RKolexeXhixbfJxxMPd8J2
QF4ch6YXsQQuzPEMtx1HjHOkSIDB6KlKDipgd/oAvgr5MZQTsde4+2Y5lQ5GZMDl7AyzfcAnE10s
1a0RFKnMKf90kaWOQOIjipDHIXltjb6Pxk0Z3oiEE84txHIVxzzmaqY7udGf3ulzIsP+AkRyEeul
A355oXlVoFONVvNKWVm7zJOW3K51bHWJiXhPx//dPpOqihuBsAj9St8sHC11Wltwgt3om0MJOehq
qmm1a/D0cXDaiwyyMLX8bG9zQqvUMW80wGzi0OWUpDvziC7JGx/wjzTGeOV8P0swN1zpkmsF2TWc
U/Lx7gqss5OgGG2fbQSgLEHA1fH6bV3cIhGRUZxw3KXUPIbcS4HFmQzYrv7fPr5gl3BpweKiPQGJ
30xizShGMFlf1xq5jCN2wl+jiQhl9+lk0otG2+2ugaRStNEc/W5Wqh+5GubLiROusOu5MU4gfc45
+/wI8W0SPW494NlMlgQWYtUTHVpy3lD0qgHpwDPTbBCeHxN+QUBOOrj6K0Jp33Ihq/vaaQ2/4kB0
to+vBzoAhpnr/MHAp2UatV+9laIWRR0263sBgkjAlPXw7S2mnvA3YP3RGdGyoRYxao6T082+3mcd
xLlkrtJY+LU8Kr9pV5uJ8VGrPHN60DCu6349jwE14thTLxK8zGZrrMCr5Vk4PhFJVWKaClnvv7IS
xRu/qxUM/zkjCGP5v6nz+zeZlLbkR7ehiH1wuYGJa/WF9QIMdOjB/zymuOZ4eN+lS4f3BsPsG3hk
6RqETGCeEOmveFkHKddg9xnz4iR7h7JTWvS3+1BV1VXqH2gzKMWVFiXWLH+pormKbp6QopEAtWlb
fbD1+ftLO965jnI7Gb9lx5fbhhfCHyGJlxjwfifVIN/fi8bCO6AImbZE9SOMzIzPQzFiQ6SeO/GM
PL1Zvggheb2QFAPLtp6GFUNtA6ksD5Mw9XhhlWpw1dQhDrjmld8nPDzy5uQarsJwTz6KweAuWOn2
0SeTGPJGf+rNWP3Fr3GEXA3Z1AL6nb9sf1cc9ou3lNHphwkRrH9SJU+BPfKVnGU9DH28hDF+K5KY
eg6FJFkyDAWdoHVg8b3fayGKwV3IBE/InNVCBGKigQaJYPkIwFVeY30FCWcLZMw8XS4LwGavQDf+
lCY/bnOhF5+jLh8PGfMij4AHNvgFxfcAw1pH7VdQRgMelVCX+2UoiLd3eVGFbVRNiSHPtvbYfzPC
IkmPOXzWZjLugmXsJVQzpIAV1L5jsfKd2He8mfmNiRTsCaFPKWY4Mn3ZFgfLfmq9RMcLmXJfTL7q
QkZf9kgJ6V2ygOYQj+uuI+eYOF1a47+YOKKkazmeshpFXMXP7RDgySLcLVBgOpySq7oi9IwThp+a
sbjMmfwjdwSRxVEDrMOh6pwCp5sFniQU4S0CsOlCeZyyNl92jEK85tvtPvcen0OtJ23GJNgELXCM
yWk+cAblkjxuQIybQRq8K0hkftB8gp/vDRn8TmHH+HBQuvd6HGokZO40F6/Tb3wO0IEOHWo5tXbi
NcQr2YzcO4BnzfxrMOJs2D27zkjAXV/T5JxccE6U2IfLBCXUDpBpWAQQEyqSuNTwkLqLlTtqIj17
A6RRnFfRwRY8Ms+N+86lyipbukCU0wpzjGIm4q1PGx7QqvIvVoxIqkXnn3Qxx1bXWDTVz10RWz10
+WyoHmeb99JMwKWbgjHdAcBuWS+1YGeoevX4RXYOwbT0rkP0Mn3Rr4sskJiTkH2CvB2PLXIpbxUj
tFC+NORqv3PTabEHxWQ2XcykbNDdgfV3gvIG3op6WIyh2oEf/PxOjvAiYTKeh847s4A8UBeMZMjI
CRqnp5DcTT4HVB5q7k36/HhKdbkGreU9CqBiCKkUnXPC0D1w33jBt4qH8SX0sSvFDIQjdDt7yB7g
cmWf2CUzIUn2kVKEkbWMurZRcq1JzNa3BgvXPxDEx2ygvYxVcVTIAWvER2xl8fr0lJFQgyhb3xOY
UYS6wTXGEzAOms50/CppsN+9N1WdQ+zJdwXeEW+vYO9Ub1IFGzyob4KxuC4uls2MY4cisua/Q1x4
OeutxFU7p0rFmYAm7IacbE43MQ9SGq/iOZc3oo7pW48TnlbWbQeHdkdE0NqJO8GGf73md/egW5WY
sOtUJO64WH3sn7H3otPM9UhX4RO4Os+eCq1rkJagHvBE/ihbK7bGt1QEiYZs68MxBeRVwjwbs/XI
E59xtZJBoCnTP6DLvKAfErZbxXYW6UAw2q9aJ6JVOXwSKVrGzMP+4xBbAGrqTu8p2szBcyBQIUoz
DIBkFMRSrJjD/Z24i4aIhwDtyUO0SF5kI04Fy/+GxfDjnAyWikK8Wud3O4atEqx1yRjpSVKMMCYd
JytWeJc0fJ7xIhqQdoGE+Y76WrfLku+h0VM9LxyIZwTGY4Wtk9iPHSXeA3gLFsajA7MLNB+oTG8+
xAd/VmQhyyl8jkQXmRxPh7lN7yOIDhXA+6HiSTPgFhibaiIT17vnOGjD+dOtH7rCQlvaWcvWtlik
XpIKJzrpAh6VeQrgYHa51Rel6AXgkzc5x0opGW9MzCupegcE+PEV/enafDNhzjXw83dQw+4chg9c
fB3lG/ZKKCgJezAESLiFmeKnw0IKA7h/zZsUNMyVKqK8RfNlXb3K4v1NvkWednSl8+ujhfEeVhgt
pAfE4e/zhPJDCGzxRsJcCgVLP+iwkVDYQ+a1ZgxKoKxIQD9XUz1s7+7So62LSx4YIbQIi1BbmgsW
jTE84R2kjP33XAsy3XciqlwVn6400F+qE00N/z5x6fcFDOl/jqOBn71dW/FM/VxNJGFPpMIEsPEC
yLwJY5JUkeegUjDMPEjVSzKuPP24mk0bYfLTJDHbe/fWd9kQRtSYmNjfRuKtZmC2zzYAJCeRDAH9
LMrggrGrTerwP/wbL9TxyF8seg3rvfjwg4pNdZdpuTrBO2i/nUk0hgp/3SCAflueVs9Adv3SbBrj
+ZRfADMz4QYkzBUkmNXf0nJGN5XNoYusTDIYRVW1Zje+241HdkAO9iGjaZogNozNrSZhMr4gPUJt
dcgaNYMf98H4Lh9FlF9vNnPOuEF0gBQC9MUjDXC60Pk8kxuSr1o2akH0V/xr/mwhhSwLe7aZBAin
zxxVYenxH20zND9mFunRkTbWZ3/ULizZnugx68MR+sn4nSwfAkXzW0WbiJcByrOEviVrMp3lUBUQ
ZxZMtNVJupbJTqTK79ZQ3GtDP4ZGl8DgZ1NqmLL+2Ua4GU3ADP1qD76s1mqdtKYPr0H5DJGlqaUo
/RYcnaB2KvMeInH3+frFi6Qj+f2MYgTIfr8dwmd3epAak7HEZTggoYuCEFsCf/BY8517v9M/JLky
E6Q9VDcKdcCZ+w9/enE8t/mk5pCDjV+p4x/2vbyFp+UFW//Vs2nNlSz2iXaiC2NjYzkZRi1LG1bn
XnJsZZyFWHS8vclVwdswiGCEqGi4prSmQd+CUE8fKh1Xh5pu1Pqa915hRzzxmUw8kE2GA0Bgdj6+
KozL9IcvB/WF5+GzeA0WENl1tkRClhu81Z1WEFtbVPUpzFCXQiZN9uQpP6b69kE0DQUkbeTiAofV
LQqjgG6KwWNG32OqcblCTQz4ojDuKJIXyoHozlN5vU5mOiQgSkRjJIeklv8ILbqCHgduLnv6jChW
eCyBAvS0W3UBLkdgtxi9JgnB/ekLTUWmzeVjnB7ML+ZvG5MCY9ZigNr0oc4zV6Ka1HotbILFqUUU
0ZtItYutn6qqQBdTgmYWWSSzh4yqDRft6PDWQZ4OP/9OnEk1eao+Nl2aLlJoqkCQVOsnF445I2m6
N4zrkfE2/7/m0//ldCInMB3f0f1qUyVthkfs8pL4lDJllrjv7ts/z8Ek9lOaGD6KDXUYc9BfjWSs
RH54OC8maKaz5vLv/1wjoewN9mjEvgzwhRd9YTTmnotaxNK6sKHay9bNwHQp4cFjgHfqeWakOZ72
dyJhjkfyuP4+0jlpOx31HXgtkq/H2qU3LvEDyD2eBSAuJ928svaq94osqpXI9tnU/+30bMSaawnQ
7imvesRGWSsY059EHjExU+Ey5Uw/urP6ppM0f9Pj5RXJP8Tw6BX0uPtKst7w7o+AnQ0WrYSJa/XJ
h5o1puKhcBh+R+lmjnGPnV5nYwRYQMpfRW6Y69Z3RqM99t0kgfb7DFaMfvsBG3A1AfymZN4XIf1K
/iwzS05lWIw7ipP6RwYSr/v//M5GNcfQY92U8etnAsAsnoA+Jnptr+38tg/JHXY2AdWh6LGmaO5u
Ztv8b37cNwtvKtsVf6aXA3T7TLoYN9A2757PneP9pvq/co6PYr/1QAc5PA/x8Mkqbi/IBNayG1mI
vwn60pdpEwR2Fuc0m4PBZ9Vskilq9fMBfv9bUdo+EPNjFw7+r2Xu6LyZgrMUUBEoGnyx4cJPNVqH
tDVRVcXcu1+kKYiWlpRXVhz3kI6vQ4NqQof96iNpWDZ8TlUUSCGtW2K2Mpj2puQojPsSBOPBluOQ
DzJcOJU2ZusQZ6lIFaX0UklsxQyJ2+BKwBDSNhQMJOpH832vDZGEjFtLvM/6N5rDYB0gsIQLNzks
PYFxhFxhGUJznZmAf/K4xwuLuaAuV/vjPFjDFvnnjoC0Uigd3jBetNf1WL+nEQAAGTnQDDv4RID2
6hZZBfiXtinkjhGLJwdJw2XmzDy3EbotGcKkG+Q+CkPRhwUttD02wj30DQNK0tf+haJj66o3wWEr
6xacrKnqCq4AjR0B8F+UUe/OYZe5YCPk/5nnUXaMVgIhhm9zJ6S54Ctazqt1HooMSogZF6jfNod9
CbBmL7x4TYtVksHpdUVvpAE5yHDwGGE2ux0Jq3CduuKgHE4t3xeUNSEchOEPsLidDBvvAQRrFkIF
yNVzfQYjxSNcg8cSJCxD7unlM37qC/NGO0jIUQ3ItiTdFZADLntu2urYTW7nHqKfHdQQeOU/b/fK
Fy8nqWg1QSbAR5Ka1EJodN8WbY86QHI7FTn30I1yEbi6ODs16Tyac60PUUJ3v9T3WVQXL1WHPh+4
tXRSqulX70qD7EUDdsURJORiQGa7mOx+OVpjocyxVR6/0zTHUzk9M9i6RDUpTBH2LBSx3ERd4qvW
+6EVwy12okOQgLHbZbvEB4aA14FJ2/lpo2QqpzOxZzi0sETSbsufYiaJpDyMA2FyfSI+5FAH2MvR
6pbQTWRQS/lxq+Lhpb0714S8OoIpCtbwKyCGqse+HNH0hk79TgD38VvHlfvWW4+sqKo7npAsQeYS
QleFn5MT99Ay7y9qH9zQDadenwpVcc9WaSnuOuWvYZ/7UxxxVJL2th9/Cz4k5fwRuLUlXvNXj3nR
um6Z3bApR+R8E66xzWAND7J5KNFIXFsCYDuuZT1XZoC9tT70xcCQYscVRkmtj+Wb4h8A0Z1Y3FZY
rl45a24BSse47D+fkCKzrKRilCc7ZlkmQ68qAt//VaZShvI2M1veQHbZHIYlTxX0h+Or68QEIbBq
jlKusd4K7mlevgm5A+ppfbf2Zd/TdY/fOPSFl0rbaqvsfT+2zBjolilnTddnUDvkniXY7y2huXw4
TdcMXMfBtGzoNWV6vxvy9YFmp7FNypybX9epgw2QBPCK70zvuAWWwpNGR+PwtNnkIDYIiERy/MOD
iiQXkAcc6uq9i3K7yZWBUg9oPX4wolfTIZf52OfdYG2B1awu+sw9ogBpqz9tdgkc/bTZ6KwjKH5R
ZhUbOEMhjbQ7zdwaeKK8UNCS2Jb/pqEh5drezNFzgVMkQ3Gun6qMi775CCzjBgNs+QkhcCwyHFhI
IyweR3WQdnJ+PHMIlwyjCn/fX8ZrWRkAmwDX1q5ZGMfue/Pj3FTr3DIINIwiLoWzUDPyPhuCUwXc
qWPX95cFliLlbxJqJj/6zNf321/ZrqqEKBxxilSS4rsrEdDYrOCdY5n8QMW0EO1SdJ+MRtqoDfR9
k6ODN60QE8xabeJ3pcRur/1cGDIMtnMtLyubF3iRYzs47Ah8OBqo1jhU2B74hF7SlcmYBze3itZU
fht/qV7iyIqdmMbZOOxQGJQoYGKaSiOSyj/BAwwv7eu/vGfDsU+86VkgQYyQZznI8e07gSW4RSjI
F2hJ3nxB/bMDHqlPTB0PzPxDrBiLWCerhsO/9V5d05mPfZK0/6T9YizpNxqDRrdd4WjpR1FhPhRv
8CErrzYPFoJvUTIIDXW+qIGfxLjW9WP7o9B4WCrMpoXlRo4YxU85TgAEnpo3wR7FrxKhZAfnN4/5
QF0Sm2CsIpB+Jc4ylfzXNAD6XODXL2V8MBqbIHdT5hR+rfznoDQJ3fA8OPmnqXubbThaCziQC8Xy
A9wUFfHNDJAyrefa2+XL62VhuyDAIsmBfED94CDQ5yvzPf1PF9uk308oYRe1pxznbT39pBXXu0S4
2BBnAFXvwI0SsQylwgACGMGFC4KdwDNuUPrirW7n8ZJ10nGaL45DmwXw4ThzjqfcK820sViD/CBa
SRySrN2ryTpB1/fJZwAKh/G0VL/Vv+eEOAXIcyWLsroUXvYKzV5KYKnGs4FZ20bzhLNeNez0xvDI
+kOWVab/OfKufA72NsKdyjbqzbMHb09MI15zK6zGhVLRq8qWP6pv5OdQA9IOYb4y7bD9X5FbLSLN
JuzLiWoa/IELX9qeMW0jqJQFYw1N2+Z8pF/xhVNDRnofBWdPUsEFOY2Eiq5egoJn5+wGfiwKoH9U
T9Q5pKJwVTRwj6lnDvqXyEa89bbQYfIhujgtF7LM/gSfAPtTQckhnwAXalGBy5Wp87iIdZYuDjev
Hxot8KYnXhIoPU4XTf4cweMwUSUs5lT+jN1E6Jn7xROtw+TAdtMx92NBWpkc9NPcxTS2XePwwmpi
/zWUD2oI3vo710bVFhWmGzxg6QejAaxuFzooPAkhH55UJfTEQcsc9PbCFg3z09y/NTem1j4I9v7y
aGxNvzQo2Tnp6E3Y7Lqj1BP0iuOIACX8MPX9goTDeRDja5aBguhmp2uN2Tx7h+SaMWd7896o3gj/
Vwy222VDjPzeLOcveMhSzlOgQecqZMV8semekPv9XHMHlc4an/yg/efKbv3uYWFlvvyr8mxIEO0b
O8k8XDiA44x0Tj/8s7TKLf5RXGsGJ3tqKMYQLT0+o3QweZCFqZLE7kYQ1ZdHaB1MbCnRsl2IUMr1
wWZGkhvEcoegDw/g5X7nFiUAMCuOPFJeGER845ltLBQznKP0axFp3ffdxQQ3fW294hWzq+Is53Y3
GsTV8xlvIZ4VulCVoQrHN6WtmzoK8/NlQ2glvpzwxpf8Z/+zpJ8ipXMa4F0aspX6qJyrgAe40MFh
pa13xShLfcOkovGCfISi/Nens3i+vu8DE2fulIC7LrJm2j9hei5Xv2/2WWeu1hl/Jm2A8u14bpDg
THcaIYcjDv1KgAhFr24M+73u4CN4v1A3DVyFL0/vVnRV58SAEfyTf6zI/Vht45HQgldPtKnEKi6o
5DTjryT/GAl0A8HqJPZ8BujIVl7FkqMQPdDYkw/OrZIma/qbxK010Qce5JTj9kAeWSbh5j8v6B33
tQJQUaMGOuAPavNfXCvx1LxAUce9b/OW77p25B078HkI92M5j7uxEhLsbbwatGLyGiOczSwmoY0l
yfO/EPOsgFb1gxrgsKwkINBveKIslKd3DYwj//Pf2REbZtwI4apyQB1TQBYpYkgr8QZjdw8FHBVp
HjUN9+QPMpyAtP3Vd09VkNr/6/bMYA39AhjA9skwBsQxSg6DUN1FEKKwctH1DIh2/gyqpzvcrFkE
gn/xdRt/4Crwxm5a9iCzk14VTzujqmx0u89FE36rd4TrEYxFR+gjbRQ0QfnsQRbBRIpus5zeLtbZ
BRZpfHBYLi7ElveJkolzwYWzj/yb70l54WR6SkRVF3g5DhJGtvli/rpYlY7zCYLWrYckwaySXyhf
1chOJ51tf2azAiy5V934PyklMPZWXFYhdt0bm0LE9l/D/lCujm2XlzAiNuVwcqN3v9F09Wl1oVUX
m7pgYh2MJEYC6arbO10zJTXVT32clhJbtdSyXMC3AyM0qe7BcUNBNVYx0zjl7AMDyEmDg2Eb1KvA
1MUgIDH4VS4ymf3N3GkoOm+EAMt8js00bYdbfcKsQC6rVxxztjl9cCHe3ujXio2O1JiHh07XIPKf
B3GpPuUEljuyWcMpj6eVszYMKKNs5HpiEKDyhrhLG2uX6VEWTRtvmS6cXW1T6jr3NGXA20Q9QKO5
c6ImwBaJXt2EnF1mQXOC6ZirNjpceLiZBj8h4jJDP7MNBrFBJggU2Tzq6aGSwVRRqwEo4WfkNl0M
HUDxqbJ4+mdFGW73pQYYY7llfG0T9x7TionLN6ZM/QkAjSeo5EWIHSTtXqVMSkRDC9mFYn/wvAaI
l2Ojbfo0cupPtPB0jx8k5vVSCt58Q6c/9ZX6WsR/95rYyuNxPk80SQyVROmmk+JJPfy+76be9CdF
7V0YS4Mv+jjaDWwhtVKZg3BYXdv0P8aP4NoZiZz8u/qtuS1t2wZSyEjgbBtetzetvxQw4oHaWtNJ
O7rg28jrXdR8f/MoBdpYi19TPebwJXCAImXIrKWvC5bJbiv9bgxl4RrNtE7pUcNOJ6YcgTxhNhXR
AmOx/7VMIPUc4pAPvc1iN+my3qFnfBmtuAZuseHr1PRAhWIZRZL35LCetdccd5fnbSgHbMiMoznH
xw0FkxQAj1OjgvdUQQLsX3A1WhJwTM2QuqeTyMZUMgcGNOsgxEu/9OFfYZF1h82sPmz/7ON0tmfb
PktN6iQWwVE/gmPgOh4tKY+vZWxaJqPvCbHcqnhLG805lOp+hWoP+7ETs9WFvdb3qxr+QyRDKyMB
+XnaUpAebn8hDExFqEwEBUtBmixk83DOsncA7xyvAZq80EflEZAAUL5XKBgW3sg63oofw0uERfNL
NaaW4K6pI83iLHruTpZFY0AGM3km+83c8jc9svxYCagx9bn+s1y9uFSX5fB64iuTZWGeZ9EYvkJq
bZsTNQgaecJoVh8lp7S8VKY3XVQMbcowvWJT06FrG5RaR0sWP2xuyD+vmg7vgPdTNr8b3rZml+FU
VZl/wu32Ycbk0HjRZIx9T6uZkp7C/wmgmA/i4yKJ5uEgj5v3Q59PUOEKCEZSp9RxJwYQKDUHzOG6
pyNRw8w3LGeG2PwtynolCgqLZsNzQHYYXruX+WN/HNXk9EUY4+PkfKMkONEHpjXov37EUd4fxoel
ZFG1z1fI/QgkNpL5MqMY2wqFgnnJYAle/gsPunF4ClzwzXZw6+Z/4svfJWjSslh/W9n/yYqRz344
2/E6v+e10TyNCvQtGi22aWC0s9gm0/XAh371FaRm6bQ0HoIQ5HzS14A522g3Vkif1YNXYmbgVkfs
a2l+s3lArpkpQsU8ayPHGwxdzNn5pLwRHqxbUxPITmNhsLTAQugcAo1OCrPTyuKG6YO84UNuWv5R
pvxyU5f0gOaT3MAMT/Lwx6n+5ZvdiDS7UEvMWjCUA1FPLFf0DCqXC1ZYjlp7W0asa22yQNHTkctx
TIOtqAPVEKbQbT2pOMcdjVjjDdsF0nkqUGkYp3iECLl4m1eStV2nwcY8cH6CnHDJAMF47z38UIYr
bD864V4iLTfGFc45ZM6EIaqZgb7WYanC5BLW4K0oy0MmqwBPQXL7g2qmCTqxI+Z3J9s3mMbwESz9
PaWJSWo1X/NJNDLlMyGR/0GZW4ftFbssewrnA4OV/CuIyz5eQPlyNdFfAQkDxqA/IuQzVeYUR2Wz
MJHRmyiw955K/P+DNePCHjP7ClbjZMkFVAKRU4fXT9bC7S8CvACx+Y2adAv+4ub9dZBVWvMa/2vs
rlZY1gie45ADCh6fh1yT6SAXa7UNrvlIq2HwSyF8AXgeZUg8fn6QCcsyTwYSAUOyWhW8UCF23lMP
3C+UT/rzmkW6iylEMnuHeU+WbsZaz81zQ48z2K2o5mUj/34rxgTZxVzBWtHpjAwz03Bnfaun0P8R
OAQApIssd6l1MZ0L3+C+axDYSVzNQ7aIaVCb0lHEVEijnTRaPpskP95OIzw8SGx8ZBYD2oaTTLsd
WnyXtsO/E/RK/3G+txK7du7gP8GzbTVH0nlC2bT4+2XVLHu8wWRgTB9l/+keXiJuMV8/5WvS+gn7
K6VLLsN5eNSaGJ354uiO9J4wgtSoKNKT6Z0iIkJGgvdr+iRbrA7dFOXy2cGGcmyIscUmVTE4aaN2
RT1O9SZ8cQ5J8+xJp8XSETVJD8uh00nzH4SJDxblr0gFgeoM7V9IwLWw49kLD2xyBkOM504we3cM
/pfSQByY9lUHyi5NbRoVn58Lr0KP5dPazTXwP3J5fPdB6CshfULxBqCZ1BQ+Gel5S+ldgoIztbr/
WCKd0BZnXPBE4wkgct7SFPy+5s+vHwtf+h+YdNE7t+1k7fzDAZ6ouDArwsxP6oc28oOgE2KiMcTE
b0zcnxehUg2YyHn2ecJmTEbZJoLcyex9cDKYUr2GXXoH8Kza7WdL5Ic7KS4nqw88Zshl6FXnSdwx
TyUixu0zRIeciT12/s65j6cyrxVaNmXOvzAPuSs+V5TvGgp/3yF0aC9B/KSAaAr77Qw+gW/azDOt
jTLqP2m5Y4oadmyxoTfWpOmBqRUwh/WV60DFt0RRScyRjKKX9QyFhUgIprncNXAqTU5UB1tClBK0
gJerrRU5zkijXZ9AhDxzWu+tjdPM+nCBP+e5hZXzACyNVJ6zKskujlE/ulLqZMINYPyGoliGauW1
q9gSPcvBHXoACpug0YWxzFAy9F/Wh+oPYy7PUwp+pIxg3QkzPQCJCyYP3MPDtE4HY5ISzzY7lSNF
4112VHPbZd7zRebUlfuFb4Kq8/r3OMOpUbRmU2rAIcC1gRtVV3EWVGMsJ1NfKMbyll0yMcgJJjT9
DQL7ucRZj8OhVtBYAMBJAC1YDQPRb9Olwugm2vqMNLsJ7xCu8Ge17UHxP55dHw847ViJKZUmhqrx
z6Rmio5IxuBPvflAzYbVuSNI6TlOILF5JMb8fH6UTotWUvxfWMx3/S6PNJ3kK5WgaPPxWOleFGMt
HwrY5y+9C4f3gkFurgeXWWbeSv/AunXrEK4j+iU9vOI3bkuphOBQmmeVHm9N2ItUeq+uwpo3L095
BpQqJ3FEJNF+eDSjGi6zODlKHEgT2rLCB0j9EMxjNXhXxc5LU+hCiYIKwHiWWfQeHZ1lB4EYIgzA
lZdA/IVqlKquHwRyHEBQBKOzIXWNBOLn94wFC2gYxXxsNPQ32IrGXKV15sOEu4TcLJeCi8XOtlfb
W80aNDzHfJTI+lbI2hyN6VLBwEaHL4qXs0rKNFLls8bk/nujq7Qzrn47xC/Y2lcpU4QUufEfDfu7
N9g829uT5SLTNUcxEFbgTg05Xl9kFmPXGU2PJdxokqdw/BDhd98wrN9OC6ntLiB8jD5RgC5+0/S0
FpkTGXu/xbhm/1As2sqXoy0NbATPZ9mqy+UNkChtBBC+8tti1QWsaMWvQhz9jG5Z1iJOfcEb2jDb
aXy0vLArwN3BaDsmicCL/yjhwJ4GfaZ3AuvzBwVPm//bBYmc1sxvJowgxghqLvx84OVhKFyA1OSg
qYWZqFK3xII4Nk/sY9ZB2o3ByU4fGZZTC4AMjRMGJY0IaZ9tjVhwUKPiLdu/Xfa5yp+XFwvGr1/9
icQvRul+9rfvDq8fTrKu0oxljKTLIgx62VQHpm8YhRUp4DNb2ffeWRnMOaMykdCtbC57q5FlRLCO
/wNV/gGaGHKpiMWT/1ci2Io59jgCVgOLrlK4WCx2Nad2u2dLhzL9c/CCRu0Ebtp2UpfmTCB4Ph68
uME18B5sAvLgkoJr1JoYrc6sKzzbDPmXkRPpUAcUKzvMh8lDFFQU8G3LC9XA71k7LhEdHjApyzXR
jcOkRy3utpbCBcrlH0LObxfQe2kaSweYfu3BIlHOl/qOiULt4Wi4++fEJULO51qIU1PeoWq/GmTY
lSrg27rgRHgbXAmpOqMm3DoCGV31xmkYUD1HJjjwMuDqXYhYwbFXfeU9Nfez6gO0kvbrfa6BToPJ
WHQtHM1mbJ445Y4C0VxJYXzlNdq6WlcmsxiiPvrw7Z0+QtnYjL6FzO4x0MibfBiG+9UKkBVjfyYi
DKIEZOqX8C/l/S3B/F4H9iMAA80XFvLEl44qGkLPhyxzO3J/ANE5ovUAIrFBFcEJAITnmWNv9clK
VgGsUH/ynxefXrDv7udLULAyAbkYgFbw2aDKwb+jrVg+EJwa8cWKaBNoYSOHbIJAqX7cgpt3CXt7
oH7YezriHzN63QzstdhURQDflMaqbWDJaYdI9fSpAsQi7Fv7klUt5DbzC99L5zKZCrcQoSgKRprC
GftK5ELMSHukh923/9r+q2JfHEbPQBkD/PKUGb64bySU6XMcO7CgfRc4FFgJTXBSkyYAkxJS1+s1
mApkdV2YdP2SEKxYqYDoWBvwbe2ZD9kq6XFCsOg9Dk5iKIyXQgswqYGohonJDhDujv5QEWDoSFWX
Pkw4foO1CbZSFfKPkHuZ1S4B0d8a3hBBrC0n7kxas0wRfla0WIxaup4SCsyqGmgGxQlItYD3EGlY
+cR5vrixSB72+PsDM1LnsY0GrBy71PcrFWwoyM/63wVa4kCSvhUf8/UBXcvh8wIS4VQA7IfS70Ho
b8zWB3RrQGuM7gWCTyEcoobTw9Ii0JYBQayJDHLuhFh41U+CbncjZuUt/y4dGovry9HZUdQZ9VQQ
pPRJ7bSw2L5thkBixRXIANRTMkPLYJ4U0sTncgmmPxOnN17IQLfz50aMU9K7+ib95bmEtC4T3p71
MFdTyYP7a1mrBdK03uH5HTVwhs+6DCkt3junkdXGGLvqmXuweSIN3OvA23QLMN0xFjmvNt6bmp7m
uiaqrhLGFfvutXmNUGR+B5H5v+pfH1nwBpFsczSYtG0KbWF/FnSCFprXqomTUAFWueYuBv/LElmY
HiQ2ByisRD3Z1i2hsiKOemHADfN1cAKtJ8SnWggJFyc/Ws8gUbyzVdV1UzHAP1q5YdJQw6YxH0xK
bqPslzVvK6MRGSEXnL5dLZUfTjH5c2+Numl0Lx3VYey8TA8FnSeNoNwXScLAvqOIofUuum/9n++q
Dav3wxHvadfKPb/n13NZUNGu5jNF0AVHDui4W2caARQYb0q5rEcQXIb3OHllae6UEtFnUmGLWm5u
N5TXPckBesFipn7Uz1TJiyjoGZ+P01JDvcZjn68JddNKya4Zk0YUdFGbQdZsUxStEVGCb7cYQkH6
y3GqoIW3Zwgw90l3AR6O7vVLT0LltwE7Kx83erdmTvuHQinUjG9/Kxj+wzVJbmRN5WYXBoIpdCpy
TlJEtdRlN41UX4qxj2R9vcsCnfu9Yvpuuqodtc2C7Qb9gCRjFaDitg8NtGyGRBdAlceVNiqf4LgU
Lmw5UkNCQX6x+q6KmmEGPGnIScZzJOKSTfBmr5WJNQFpU+n1bH93vnfv4qT5XPGpC/4AyKWHT86s
W/NUvR3bhD4d/BUdRPMADG1fzeLB7LzHAPGN+EGNbgyQIfIZegu/9KYqtBAYKZHJsP0He4Cmyabk
YXS+7pIjxWpk0MbILVTxJyEdmaAmJO15ndp6SjP0uKU3gaEnchEZJa3d7NaPuz5PtuZ13CeiOGDv
uZZo4c9TQ/ZTvYKz3FHrtf/e/1YjP6poOch3JeXrObd8C+ZM0fK1Nr0YsN6Vp88rNECwjEDCuC5o
OEyrpyRN3RGOyYs8QyjrgLWEczsf8h+BaNGnvXDcJr74EsS2gYWsNKCEn43pkzXDBOOsih2u4Im9
6vCsbWVCyGV3Wnl4CdoAOJ6P6mOQIEcMzmH+6ZKjNUWKRK0XvwcGx+R/YVH5vDkxQP8YFnAWq6Ie
pTJsAZUUfKMG//MTsN5uEETALGOAbS4FwEpk5INszZ+XEdoup0TOPi+RH2vbR2MWL3NanEtSsD4v
erIPKnbe17WFqFUQIxIxH9soALQTEDiwlYT3fEzyBAjTS6x1IfgPgTuVq0UN+p+DBbe2E74rrFtu
adc7Cx6PF4c6FPyucEvLz7xyTjKjaHWXbklPVxc50RigMgQ7IauNXYJdl+EH1l6Zur+09B2j+KNU
9GL/XApXpvp4nbi+ydebqgDl+W48pV1XAIgY1GR7YQ8pemfYicG/nqZj+ZBlUbOSfJp73yHPOeJM
/S1PeoF5KqWrrN+WyD3QsmpbVYKJNBdlZy28O//rXmucYgsXipW+iOQkKcXdfvLqbbO4gkjyOn7I
l4nfdnNB3z/NuqoLSxcSjwKq6fZFrCyN1JZXgPL1Rw7d6o/ykuoQLjNBAKRc03EIRlN9Z98BaJ47
XnnXeolvpPkxB/Hn9WibZ16fY65NchUzmtlYLQd+OgnrL26h9AeOPfbZ8hsbigTAr5tQAvYweCaP
V/ukd+kb34XUaL8rvXIM4pz4+MlqR2ZRMSams+0FbtqoX85RnUj8EaGo1Fa/k5Yo9BYi0e5oaxdd
AhG1287QNfxjye7b6o9GQDDvwZIgyJHulUPGBEjRUgP++Seak62mdHzAo4OtzM5RUN4eTJC5zCMl
JpDmD3htCexmtIkYvo55weR0f34RmOzRRrNgxKmcAa80SiugpXJ3ZDlqQ+9FT3UrkNe+a/jR6NaA
2EODhMPrvxXqufxUB8QJiw56t/Iw/a63igr+olXuw20d+eGNi+0qBNUDJ3Wt7DurylpjVKFkbSKs
ufoNJP37H7+dcZGAf74sumSn/46e64+NHSpN6IchWFy+qlvMUMqEZMGe5enkXILA9xWhp8r0bOSX
kFyT6YS/JYev5iIufplhGniQMnKDpJ7pgtb0Lxo95U9ASe6aInIP0ESEXd+aQsvL6uHQpmIapxyw
2XypYVTvJMxfW12YKDHpmj3DurWeXs/1U3FsLYrP0W6/NUS4KkhTLloH5NP7UFu0Yx15ovX4rMcg
BlKkN0FsAXlj5tVr+5HIfHx2VnSHE/cJiaCM4fGX7RFtnTxA+bFm8RHNcMLGge3C4wLidZy8ZC91
kbRod0ZEHRfFZG6hydWUX6AlSAOoSZzbxjtwisCyivhApJ0E68bcRBcKOf7QIcwoPTE9HuX0aFtb
8E2XoEVbrCX53XNgpnc6Y5/RXo1x2lSp0/EoyYL3JdkodrMnQ2mWKQUu9sEYaVqTK8zrlOWH2QBE
DqzCaExFgyPaF5PIoCSOJMaYkycPOZ4GIRn77yUX9KrYD00hq0BSB1V7OKw9rT3i7QuFyz/MmTcF
swIFoqYtWBAMPxhueYGaxJYlpdLdb4oaoXkRHBdWZhWyPmD4duInBVvh0hUa43QHsLpayJSV8rEB
vX4bI3uRd8Iv5FTkouxZeIbBq2gRWL5a4kgDfhE0B4eZRLBq8muVFAqJ7LJvVsCYcZztdPRmxyU6
O10Ncublbkh0CVk8Cw9OFosTgmAAlvo+EMcgADM3oHRbwug056l5QV2WvHMTziD+1DVKcENthpIW
kizNK5cVhzCOef5HjeXQdjTvNrcPtteHjf2e4Micn2VVg9Y86FCogrJtGeT+kZ1/t9oVNQzgkadC
HMpzd+kuwhg6V/aJ9g5wOVcJ9i36K/suwDkMRg0hrukVox0gVcQcEOHa7d1+Y08wKJud6kDXTVyr
xfZDGBKcfIzvUAXdtvPrfH5MYClLSJKmCXuV1NZPKntWGe+ybO63XfW9rGohOaKj/Di3hCGZvR6N
T1SpMM2amlk5ajqwjdUzAD0k8ZiA/zPCxOiUQdI2wzVmpptmKNo+pEiDvqG/6xtg3lkVt2TqtQ6z
2vT7W2Kj10LnD/bcYEksTRLnZ/9vdOLc251twUzov3AycohpRk8H5MYo9zmqTdCDUTmdDwzqjYjJ
CiJsevZpy7F7IkEK+z1zr5KDvtys3EGHnmzFu63UiHVrwU9lhya3LqXkylqZBEYnwQD4CiV5fTke
JNo95JGDEr0eD7xCEDPkWCmG5BI0jzZ0Y6Sc8r3KbK6OYEmikSb+l/mLyYUEgXFWQ4lytULu4wjA
0UPXJQHCQ3QhowrHHRojXRddetqKdWsmS1nN45b//qfQMCtnUe2IXEuTSS3okYE6ZQxRVvBvJl6o
k0rgr6a7rdMVMDF3KB9DbtYvuH5eBvZIFlZdcTRRYfmAnoJxS1lVtxztr4EDTrVE23prGCFOCUM6
hcvfwzRQ+IViSQDUnjr6XZBr/AXJ934sAjYnWlEvKEx0F3OI/+UeDv3Q7BfqLShYUjp6F/WIPokh
W1XgCbwd6dIE0cNc9o0aJNIUx1wPEFi7bPk1phKyfDmXxfS6HS/72JVfS7aa4TlErh9X1zRa0R4N
QHTs8/Bsqx3XlxOSUn1CpDgX2BgxqzUOgXrkm+DVxUQktI9PE2TSG+QmCz30auXg/RjVtZAmrua4
5LB6yjX8hWfEpsFXlwETjrlg3VFPFQ005fLQVubm6aYqtXEx6ddj+X9fC2y+XEVBp/YuKrXNwH0Y
73AIbaDcq9zZG2KfZoT4bSuWWWsS2PJ1PI//MXYk7qMhiGgvwGzYScziniJ6DjvwRBYRko68KcN6
VkujGoJqBQNkO1Fuigbi0ib9DIWL8Uwfdk3juVqUmRo8ImR8iFmXBkM0Bt03bj89KPcTxmPCPO6s
qVxUhMuTxZA0oDNrMgNe617XbEHKGZ7WEYu9vxef0nW3cWigWr65NBeHXN6RbjHrVMhwVOn3io/6
Y3b0Z6TuzbXkeaIH/LcEjuc/SJIXDf1Xxs3VR784qgmp2jPXpj9kL6KtQiIfKLZoaWmqONauR2N1
OsBeTMhiKRO1n71vpJ86DzKQujse8KiSgbahStcneT0QcWCn9O+9AtxkqusWSUOBQX/mL10U3GrJ
A4Jm0xl6O5m/ujrvzOZ1yb0vj6Hd4lt7EgmPP2mVqAixfh02/oHwUtFaEPaL14CJ4OXxZIHpIVvx
uUC9ySHn30bqHb+oSocaWFVkSBay+u6UgDAvLl9RaP31kZRwPNtHM+GXSquGlAfbVtNK3T4xN/Qz
B3X33WMHaakin+ZqUuRwpMpIiaM4SDwvZCTDoDXJcDLG+81HqtqyQZbZjMcDFG4dL2PqDCZd9fKI
ohgZ/XU3JqTvWYsbINF0WUQ5YKFDGhs07abIVO4uGEVLdgtnj+MNWY2X9kgEBBxDPNsqCLgHYZNR
fxNkkS1wUCDgtUln8K2rbTIv2tCQTdv53dcGy9odTPe8rzVT/ypaeQXucrjQhAK8yBnsTetcSLaO
sUrZfArS73qYNOq6keI/vL5Ggkh0x1R5SN6JMFD8qePyoW19XMX/rZ4V6gytoNb4SziQ7y8Bb5QU
KRYfpUSZlQUxTcMpHx7jAJV1CYfnpg7e+5WA54Np+9ukKSyUdqH2KFC4SoNDnhjRqeYnLLatCS/u
OMehSunNYd9khS00AGINrUuWQFO/Eq+msKx4oIyqHCsiBDUjjD+uns3Yk4mT2M8ymxHMcuqYZStQ
XMeXnDAYjZN8+h4LQEzEAx+QyRweHTKlBFQDb/g4HjjkL2uOC6iY9Mw8ln/H1fWjiJY/i8skpxjP
Ib7sPBNYy/eIeyUEnZcluPIqg5MW25O91lQ85lguDGHeAenO0RdFpWVRejB9ONsDhRN51PO+MqGk
Ab7iIR3kxwhyRFIV6ixAWYTj7ijMBXzfNvpVCKq5PxKlRNoTrtEo4gpFq2UNxvUQAIISVFpdkjZe
Hpy0r7IPO8JLddfYaokfmbXaZbEEX2jYWR3qPSshVg2K41EQ4r0cjkyRYBQ08x58+Nud/9LACyPW
NOpIhYyHPvCshShfJRMN9iMAxykg5WczPnBDHVtmPi2pY9VjPtDlMmS4ZbB4SglsekO5E16LA9fa
Dg66zBTRVK9V1ztYZD9NiS+/7xBYaAQh0BQDq54PYha3+X1aSCF3k4L5wXnBSqfqWcTyms/m6ND4
C/Aj4wTHIuyIJLm4MyGmiMM4t6HcXwMyAQw0CGrmQ82acHqw0awn8o3ZydrijeJBumLYrwCbq5KQ
34TELVYmcDc3V5hqmcJTOKH5v6444DG/oXkzadVgdMtickC1trGIwwrei6AFKO2XviaJexcslRzO
1jmPoV1/rHLxUhZMaV5ZfkP9X3BunazujbnpE9qiQtU3xhaBS3r8ha6U4S4MgFWInKUDpogLrPPR
McvRRGiixhZiCHUrk7zsNcrsnuxAwR7LsxTVLh+xnWHQS5/vBgpcaOc0VcOsbocYHBAd3lhYcikL
3yzpTa8fwX7eIX5ITW7kpU1U2vRLh6BXtNApEDg8wDzWbjyyZ7MYClKySAzmWdM6tYVGFwIYEoCZ
f/BbFRPOPdtOKJVsMu8tqP4ZiEv31nmM+8vbA6lSRU13+jRKAWNtvqD/g8wWwG3VdNb8GTmzLprT
LOGFKq5qbUO3Jbox01IJ3pswe3ClHQHmmjcNSUrVje8/kEs4h2pdZuXcUzKFMMkgz8er7yx22tNV
GWl6/2X2s7QI/+sqRCZRGLvY92Qqe/NW6z69wmi1rl5ORoTzj2i+AwN9wcGXzKUcNFtHlR4bpXaG
45uORhdicNweFHWyLfcwTJ1pKdTxU0dH1LXglpmwFZDVCgy/CszY0rctcuDNcHYpExyM6B+UL4eM
VE5PtVXy+2q7pKm/AZpCYFpTYkdBgfVVnYyiiq4yGzUp0fPh0gu8m2GJNLVFIALqhRgkPSEzwEpE
xSngtO3UsiiWPQVrSRf6ePoB5jDmeXp6iii5JT7087A0c+HT8AdJwc/Lf1LFXO5B7JY0y9+IlNa7
TLUShaRo0BGUvTcIiZbPU3XoITHLFH/8IZU+4Gpm7oxEwBNoqf+mfCHtchvPWMGeSNNbJSvHce6q
xce1rpoWZ2xdX0iAXz9oc3Nrbr1Suiw3DfmfLx0k0WWZAqJw/3g+8yx9dVoLhk5fEQscMGVbqtvI
13EjU1B3mM5m02woI8xLpA/u1/UqZW9t143CYTpEA/r8nzDcqHyuk0SJB+c5rBaOSQTdr3/BsLnN
vDd8pEkXfJGTnWoIBVZZ6R1XDMpmB+4EkMa+DQbZ/qTOxS8RGOFoDImInLJ3pOPZsrJhTnZpNJ5N
RtTvaMH/wfoNED7xMG+GrkSrCBVBZsMBAJT8k9hIh/zdEQac7PL/HpO7bi18v28Y1ekDSgnKkGe1
O0wRJbxUm7BXNIkp57jysD13rElaKFJJKows0Y6eRxcKLrKar34wyUe5Y5hSUTzjQqET27OglSZo
BXPsbKDZXwQS3Q5biFssl7mPdhix+lT5doyLNauSF/W9JaFst8CO10hINQZj9bj0MHFj9u8K2QfG
8AmFm0jRKj0vrPfQGWb3s+6Tae70YLwPZnT/gnjE5T7K+tTBEYHxZ6juT1E8GYNcTfodtRFFbzk6
9wS/xY/UmO5n/SwJYdP0/2Xogg8/o0kLQfTl+fLrTPvsBXGaYQgyums+YzgW0Mjsjz47u0zcC1bg
8nc/a+5LkkgLkSRuEuschjUA3CDyoPqzHtOfdIX53L7eAwDyiTBM93RYehkCfdDc4RlrSTaL1Qgb
RPk0uUBmm8R/OPoC2Cykx+dXfXznyPYZ1iG/GOxrH2kFqUBqmRh4PWpRwd3Jd7t7ohAkqljU0uBx
RAsZWOTUoQcK0UkY4uh7qEAxmU+tCCAGawYIvnzQHn30BtHUkct43yPJEgQyYqN0TFmnQ5UjSt48
3wAJLtrkUgDVaODRXSv8tJVTHT9v6oRtAwIbzlSWT0CYEmDu5JLxs8yasd+RdD4hTwPtGKQ0ygGo
GuX7RST20aio4YZGl0kUptQa9UXQ6fOWH9b8hzG6JeVh46GvppJWh2DweHOPQ/s5h71BhUtZ7tTc
zAWj3dVT6TldiA0hDQFeiSCq6+aj18toLo2XHeefJGSj3lLvgqGnCKKhLddSToOYn1fz6UcYxBkq
oYTeRlSHMpFnUfvdgB4Gy/PuEVI6/OHummj9Hp2pPiHYzun95jSnK2oiXTrOgm5xiKhuN+EPkRmU
mhFd0ljEeincsILhitoUfpotKRGs5d2w29UhzSn/GFyjFApSCQSCh3GfeeWiNVZT5hLT7ylSQZsl
xCAlfN0DAKra/l1oLWfjnFV51MgpJo4KhrjrYcDIRmcnCStb6RVW5M7tLOel9omipwM4JsBGJd0e
jYt++pTPJeJPuOcEIJFCus2RLWc0sPdAOVT3Jb5cKHuulmjKU+Qc8PmdYDvCz1uvN7HnDFi3l+B6
fnkwU0g4+LMO3ybPwxLv0KXTBLH8OwX87rwEq7WWrCli/tmVuf5ogsinvSs+6aRLJOUgHMKvEVRk
wmdZWd5QC03INnhNUfM1VIm6lvEhVjpg7iGU8PG1cm2xBeUbJf9rXJM2f7vgq/ePWleDZLG/AI6D
F/i92afAU0hOxXZ8UvYOlwroSR4gPKM139MZa1ZeXQuodYt0JSsTmp55G9LTYKW92UvRFMdDTTzu
MgYCG+7UpSDYK5aFYvfDG2PMThifkbDdGc5jFPGb28tlco4OJxJJ5jT9cxtXAaCwkmQXGJmlt4DI
bRiwDfcslMiMH+DZDGdGLOGsLgwlv9AeW0UYRL0CVRlKvR9uQlJOvKWS4KCIFp2/R+oBXI3ZIWdq
bR9I7WnCDeUmg+KaMjyXghqHXEU3Yfo9eI6NtfgJqFHfS2Br7eHn42ufIDX0IvdSKHyQEJ/kODgs
veqdprqNn4i2pBKELw0IrRN8gi39jP4Hm41SERC6V8+zztGoRY5AW62JWE7xNlcl5w3UeoMb5V7Q
rNhCrm6U4l8kOODxmKT5CKw0YyRZnDJ5Z3u2sYeV6J4Z40xKdKxGNsKmaCwrns84EwnBiQe39P2u
9VnHKhnNC/bzB8ySdOerGERy26gRNQt1SSmgidyuxrWDkZlaeHPeQtfqBRn/rbyDwQDjPOiqmxUa
bmKWO7aedlE//gx0cQiGKSQdtUfOl483tpsjWk5pTRes3mk8tgOr5TOfjDLA6SMgN1MnTgJd/oQT
ewIky0K2EtoBC7JPmUG5R7SVJNeevaggfr5fGyOviW3qVWXBrkcc2chNw9RVd1ezLov0tt0J/Sz0
p0HXt2/fDUdwz/xK4TpK/yba0TwUWjUmZmP8VopLUvVqIuLDh/vBg483gvxUP05WloMPi2jkgkOI
0Zq6FTfXVg7dH58ffqgbN6EUOee+8JBDrYbzE3+F8HiAG9jCG5O24m4VRbd1wZwQm79/YX0VCej4
r3tYKoBcI9kqizrmL7C87v3gjpgArgu1crC9DI2rHHbwZn+1IfT4x63OPul2/lxL/4mAVAS6i78A
KIQa6DwfQ1OWdoqZuf5j8twjCbyQmiDlt8GDOJERuXPBWAeeVsiBU1abQ7ZrxgnLVl5opGDWmkP7
ILJRoNggOC5fWnIX0sNlQZK0W9iTS52kjRdiArgYpvr/pKyp8ryGnwtScnPSR9JSBwAAIzVX/Y9u
Kn5tGRrUPpHcDpRKIcusA/t7uyae91hKIIdDSze+TDxAhtP8UA5DkyCyL4DPzdDNfakxz8sqqX6s
Dn8bot9P6M3I3lBVXbcp67b/q933EgpOR9FiRjHNGtj4MymLuM/JAfPBRy9vApL2EdXVWktIJkiH
BNrk3MOHH6Bla/Ix1nF+Am/P9soq0Koo2tHMdq7AY3lPqhz8JC0hf1Q6evCIN5ih9X9cUgJVCdQE
BCVnD4t4e4+/Bwi/XdH7I2h9sukTXbldIXKKMdJs9t1UrnAlrxktiklvFbLhdCdufQgl17Mz59sz
CQ0eF8k6ZNA9u5HdS51tmOOCefW22UXDxLtfWvz4N9eiUUwVkGdmZbO0Hq0mzvOBQ1Yz8o9Z+n0s
nOIwLeXU6a4VQ2qiDmdRtOwTFlC/W+6aSVwk6Byx4sTnz+XmTvwhCef3W6xSxbFL+oYZ8mbRfSJ6
l80ccaLDcOUXFTMocRnPe8z0rmnOi4Oj8S0/n3MBV43ISaCob/d6Am1RR5CiKNVPvZaYgpgH0CKj
obuAbBNL6m2fQ9CzJ4Ej9UKSuxn0AFkIqJxu82531q9oLvVcp4dnMRaHv0WAgcNPDOfghXLXl10w
5ivr/7uP933JYFZjEwdvH3NC4+GIT7Z4DdM6+zNBd7SdsweuMB+NcDcnYJ2qToLI6pHSUWGFuvAf
RwMk4AATnZK2t6PN92pU/y/C2BZYySFfqRki85LvloqRMmF22lIbQULJxSLdHat+uq90gr0d50dv
QnWArE+hjQvmQwEbzA61nhNuhWrNGaL3a098iSkGc5nGd8tEkyiWaJl6LLPsjEPBFD/QvwBXg4dh
hPHgt0w3bCZy5nDMK/tMCfZHYjocrToopIRuJuaYY7W8a/lDVk4tMMtFk924pd7HI2+A7bcMEFaR
u6yoaJuPBbKPxnp8cV5GpOphpciGVgZ9XbTpRMk0soTKpe4f7CcZT1pil+LCyzclNxypGiDyIIjM
m2nDs0FWYTloNdaVcHzHaInj7aLlciW338yM913uQAgPfS1zst+tYoA/HhvFuF5OPKe7Ez7dBQas
FCxbtcIfTT0OjwFJXHNByVh25sC1w6BEc8uIzrVtKO5mo1qB4rh2wfa+un1DhsgHeqefO/DUzS9A
AAdJEP1kebCZgbfhWBB6h7yuunfgkcLu1p5/jVzUoOxwTm7Mr11klMSMb0KwQllklbatKjhVzQwu
3IIg6xrDPiaNuwL/CyiJNkgXAM0Gl7FITcdtlPaHs2lBCmFi/gotcgjwbNx4gxminsjTeDIIAB0c
xO5Ye7ubwjwg0Ec6rIRJUG+O/qY0SXiLJEpdUWBOwFU4GVs1qnGKHLVefhPO/JTC5IpxiyNch4Lh
nl+xs4a8vV3k4JsAbD8j+FiJBkc5UXmcGv8a1t7Slub25ug8tm1w7Cg8Hsbxvq+D4cIZSHjIR2KF
WmOESiF/TXHpKA6tYZb066CQDx7WGhBgiGGhv+yrQoce/DlnckkhRhiB5oOnQbhgqlUI/kaoChvU
G7ZloOSyfCkyvseSRcz2xUW+2bUW9jPN/b2kAVuX8j3ylYBaEUMLrwK2Nmf5TFHuWpkb/ikpAoVx
31gvcAPK6EDPQ0lP/wqansuDnQPcs36fZwE6zKEhf3JujWtJMhGFLFlGKDJ8gRp9n+HybAWmcJoH
FCtbsZ0M2UnykwdVIvrV4XZ8z+4x4wNgor8/aHbNVUflhLAoe0jbH9UucdlSP95WzYtV/rY0nVCd
vmmv5xwPCxFc2ugnr/yh7b608zH1nFeyX1YqKhbaHLksTcvHYFJfVsrHHus5oSOxiTnTiHdxoxZV
SnhyIJUZpcMOhmLMZ1b7ckYrWCTWWthHJEenK1lCH+tIq9+LutZ2JzoxNNTmixx6pIJytT9Z6Lcn
4FsIWhXiBfEbbr8SIwHnVpcBt2RlT0lu9HlRf2S+2rba0Rulh4im7nnGHOQ82aCA335Cu3MIFQ7n
F6cEZCIZx5nXMgIBZf1JwfJQATRIgsTDIFyAcCVDQqp+W/2WyFZ97Mqtt++KYSz2oiH/2uBfJVc6
f0HBWA6HmC+rDPzuEbC4VC3cgq+QR3liMeQJbnMCzfkj/DsR9QWW1zx1QIcpjNpkha8u9VJJyP4e
r2xuXQFdHkzjqJ+ef0oLOvUq3dW3Ark5WKoDO4KaZj1TCVA2A0smiruZf+NalSfLxrAmJdoSgSq8
7mWgYuzBq/T/dpvVsXXQZLZGZXMR4y4MNWLn1iosihXH9XjNmvVm2wKBoDRjpMfCAHgjmFuhjY7c
BYFHFpNM5Dr7coYrXI+40Zz4RCVJiqYuzwOe9XvMIxbeWcEmljDyDu0PQSpE9yhjYnc5KiAjPa/K
sR18HQE+7s5OzhWWIpmWFaN96BW+Mec6E+RyYtqjE0RqvFgRX2JOedVs/NXTp2PBwavBfeXlJn3b
Lf7uCS8qBtnZPlZeFLj5AUCvrhpHukuqasIGMthU8iWmMBTJAzftPtnMoj/g16sQJDr82ScLeO2p
681z7PUEEJT22c65FUG6m4eKTG5lnVupShon6xwZLNb52kBDNRiX/HZ/xVINkxqGlYZd+3QD1Iuw
KmV2fV8SHKfA+BqQuxKFJSXjSJeyq2L2+kxfE4uV8W+qUIgfYRS5ylsNULlF7q3gHi/Dsw9+SiuH
vJurgyQ/ADZanmZ/0v+txN1ZVbR6FIM2zBCC98nbyNZVMkH0SAlb0BRoefeD1cjSDlDFrVwa+McB
wMynvh5RmQYjj+2n+Xu84iNQbzfgp652MKekXv2E+EUzI35ADJzf3Q1PDz1CBrxWt0Y9f/mH39Gx
KWjdTWF5qGmWl4RWyTNbPkfM/ZBveFjhqJov1DeKtaMhSd6HAmGDiXgZnmbAC9h4vbNvh0J2ze5u
P1Y+nC4EptvdGBJ9ly9H3vLWhyAZrNAvpm4e/DrkGOMWUQ+tMdAAuUqUdStQm+yWnh3f5xwlhgrA
ruM/9JU9+jzBEivFL5fEgRjREB1Z5lI1Y8u2ZdyKWIdp1HAp/zERu+A8rh5RK9Ji5MOAGQSMMIJb
A0PBhLwME5YwcZmmxwqZW1BX3yK3Y8ube0puNYqUj5AUYlwaDzXkEOCse3WphqcQoiHVRU7ncx64
H4s7D+Rk6/4TXHAE/fGlRcPRbdGLeRDuaBKIvGMIP7pfPP4CfJSh7t+G4hXIxNCmTBCkJa13DcRm
Dm1kuizp82WagZNCTjlfLoT/gXt6Ir/YUT862Tu4yAuNEcLQgC6djy0EL5DSndLhIRjqGXO5RIM6
SsNuFSzwOvhGxF+1K+W4Dj1IoTIMXHvE1keHErYYmJZXD3jmT4AFzJCtYCtsNnNbNmdMAXBNdgqM
S6ENMGbx5P7apSEx2+F/TZRTX51suQe12kkuOE1VarFSDDmCqv/ta/G5WHtxAnhRTXjRt1EjVC/l
WnODsONx78xz+DfuuibzejsmxKn4UvqKVgqffSxgTSdu4tIzZ87Zd0iVte4DKZc8M3t5PT9itSvm
OuQgdieR9z67KhFthptRvbb/Whf7qHUUO131kEC6t65n28t5noKgBbwkc+KKSLI0Kjl99eyVj3rX
E+lyWWGHJiCkATdP7IlahZliHO8DDszKs1nnrszRYxPuXSYsIruebl6JwXMLaBQPDHFAvyibPTaj
y+gI+A+iz83tNy2Xp2jEFhElSbWwWiFLuLbay81FugJtfs4WtsxUQW6w71UjeVzXgP3iJQANGCAQ
Mmv5QQ5VmdEf33T51phbTwH7sFesuCrtvoEaM9y2GHfXjzFqAA3ROE1iqJNCmPVzEZhFzqfGE2wS
2vE4iv1qCBuKByJMqqnOn9skLKhK01EkY4J8LKx4SJWcAKAyZumSfkLpKykLjBYpcyklJ/gggSzE
LpkrIN8o/4S3TL0fbcWtQPunfID42SwPn/WYGrd/zfn+CAj3+QV5+yHD2+fuqgEPPEO15gN+k1Ky
8mcZPSV884RtPfgv8J7OKKxC4jpNrdTbv9aannys2Mgp0HHCfZlVO2Wh7a4CQ9Ug0Hb9se+yOrTa
Io1FE0AL9ZJhQeWfRCt7WMKcOUCAQaCuIij2km1xpKrv6hxIM2VchSqTVnfXlX5fi7l70ZpPocw/
JdOEJmIAuA7Xarw1pasM1lgqiluawPlyT4Al5kh/iy5eXyx808SB10DMWX633fToS0quipSw90Xh
GVMJnR7e9iPBdM9zlRBXZunY+eyenFbp/DdyMCXQ+RtapsejXXWtdFsQwZLs3X0HB7FJ/SIGBJ0V
CYnlCWpimx/XqaobB9R4Xla+ELKsoditgiAQkP4oMUGYaGMdR1rfeAYtLEFuIKS/H51jtWbxDtou
3BLKCdDUAmdRyNCsE9Bj5EnYiQziGKIMtYUmXfCPUwLJpzF3jKRGFQf6ub16VsEoppE81X/Dgpgh
YUjcV6ny9YC36yiyWt6ItEX4/FmAk9C7ea1xG7xG7rQetEgpFyPGROo67Mznpf3UoPu6d6GMT0DJ
AW8U6HLVHALQz17wzyrAMkCcu7dU0R5LmH2RdxnNIrHBzQjsiTRcC+LChGDOmAiLsyMr9hgYObhU
RBZCNdwXycue81cUf7k+GCPVI80ek6RcDnvlJ+s1jow7HkabmdjS8Md2+PKC2e/ePNYFE47y4dGZ
s3D+lebolFWUQTCsFoRRmokKvnNFzoRuI8yiMOJCDicm2UAF0n9HxN4GMcNQsjgDgyjT3xmamvie
L7XhZS7u3sUsHzRh4Xg44tqznaJ5j6gEaMCFFvGMn9ccA0fodlLudaugrBVqE4XOvcUwx4KSHvv8
x/866Lyb31ErcQG7vG/maomekuXk9fnB8/ceqy4gVxRHa776hljhAyRzUMDLH21/gu3LP4Y02gR/
zlldFINb6IOKbMYMXfjiwxAz0Slx92sVAAqdGqxtIX+lncE5HHIOmF0nZ99TREpvMgN8XJoa+ZMl
0wukXV6glXx/a4OaeQVU19G9TE4yn7Z34zAfVsC4eEdX5jzYTdeYT9h43zSsTqZTaSGnwyO/5JRS
8wyVT27Zrq36I3fWncU2ObIn8d+WEwKsjMpv0Iw0l9thJZtasLJ7gqoUFac/DW1HLHLAG8RKqWSW
urr215sWAgVUOGxADYZszabppA3qGlRXMsuSXfj+QgU501SBThvYF300odzv6r7jsRQpzVKwko4A
p6SFLIMPqorwyBa+polM1JsuBGHF7++wGNOanqOXZbbLn/j1SjJ7cFDi53JxpAj7xkrfFM1SacUd
2kkuuZl1Jyn1I93GcAoWcJM6QpLM1FoH5QuxzP85ewwhgiCMUGi7fTowsthpKM7MOFKHLHs12fnn
I2CeGhBaU0ktYFQMBvt+SI68s89NQuPd/CfiDjJPmx5Vg+3UVVQWbWd3L46sM67DEQdz6P5q7qRI
ZNNC0aTwu6XSGXyo2luoBglHSEx3OplaRoA9WOusiBFp4qrIXpwMAIJDgjMtgzEtpVG/ENqZX1cT
wskv9xngOoHJ//UMU2oN3oU9XYZ2IzXi4wlWwY0WgbSoZkToi96XIvkDYrt+vfG/+ic0nMsmABwi
+JGr96/9bplH/X1a6gNm9W9ADmDPArpXtdhpnpm20Ky0dlkSQGX3B/e2GDTjMDvFjPyCxERhpeCZ
dI/KqActpZk2yhWuE86MSbE9hgkOVsoF1QJ0XdmF6suvVGtVljs2MkIjMKkP6WgqkFXe6FS5yJV3
CgMk6N14ZHHrnBohze4dm2aVMHOhvMzl2Iewubcp+uDab3WfKXuQD7puMdIqT/5mAeH8ZSx+Kfz6
rSgN9QpeZ4/Jl/sXElYmIH6Q7AHMX9Or97P3eputOCR9r2UDLE/GAxlKznyR9qM5zTvWJ2J5KdJ9
OMmrJz2B33yCFaCyvK/RRXXAZlfeZ4WybRoBYLq+PYh/I/fxfZNtzKZDQTpb0VRNH8BjkWi3bEQ+
Ye7e6JlfsnAItUNePNDy+yWfJy6Cq4RNqsR5L4G8pSpxsKKPifLGooMnbTC7w6dBta7dgQ3lJdhW
ilAxiu0V9Wadpb9jH2he2lJiwfMalkA4J3Hm/SZo0JmgmjeNlVhmW7iopJmycnC6NLX0hbElMhlC
ehHSIZ7aXWv4FUfayHLB3z6IwSmCHNY5m57qJnbbDpuKlQC+tRDfWCoHgiP0cEpd3MTPdJ6uqHH7
nTQuk2G8/E9kYp3g2Y8HMvBO8swUU6BMxLgGC7z+EhxPYnjOe4yQmJki95q/8gVHC3fWGNUek6iX
0nrO3Et3wfReX5GXjKIEnV9L94gkCE9RNZkOF/OZPH2TRhdf802H1KU+Fqhy6T+tMaI9kmvr0pnD
SISc7h+uHJo2TvcmR03xSNHps5GvQHeN19oPSIALmrfpuhijsjfFTKpVuef7N7xchC6ZW+ZkxgWy
vbI9u/oiS5BSuz/PdtQ85LX4O1Bx41pD8KKZJq93tsu8QMG/2FM+wb1nBwC3EQatl3pKtjIw8O0c
78qjCunZ/QRmgbeAwLuUVP38uacyhQhQa7UqiW7YgtEErk8jJJnp1nbOSquL7bGyN8g/I2OGn6KC
5gvTNh/Ke9YwFtChQ/ETrKFuCOZkhOc2zb1nbnnSmY7+G6SgY2KKJ6TmLF3XQFu+Cp2c1o3FF1Bj
szmi+gAYU36nimdr8dvAakeAQc5KN7uGMEAvzJdZ5jh5Z89r9rDg2QoNS2lVyMsz4a06ZbRGGYaH
ui2T8oKPgPypCI5suKZQSXqnyArv0YNfmKcVuwig5XyMeD2fX4U80LRy2R0Dii7Hay1qQ3PDslsv
L8enbrfZDzpGMZwVu8nmbsXPkb2rzScTXUHU1A8vGH57FZfI2ulVHz/mwoAzkGu65LvPFOUaDkBE
0WYDUI3pmUeqULQCXsKmLnX9lyUClYBOYSD4+Q1SY5c6kj5gGazEowhBRzqGw4Y9Mfs27xzChUfO
Kk/lepQVmEByfTtG2Wj10TBBb2ZaUVw+NtR7UkvkoRqyUBMvwTYDeC96VFAMZx/+quixMId5s37I
jpCT421tR58Q+tbCGXxMPBStMg7DoTAFdVYNoHbs6rEl4QZzV84WTSXsZeo0maFOwooAGdWaPHE3
Arg7vjEbRPStAMVI4wS7JwNfixnn4+bpoPujdFRQoQWormZ1LWPcx6zkPwMvi+pAkw4itTrg3sNO
jjS2m3tpgTG026Y7g1ksOQB/z+S57Apbfo9jFey6ofu9wxhErnObBDe1xkHjwsnpGjUjv7/DzTJN
1d6UwDAdyKIErmJfOMAtypkcuX5ZwbwBxevSKideSI2RLiKOhIg6eZ8RHa8uetXrEVnptz2RNaqw
bVk/cDCksGEbNsC7FlWpv0Wt2GY9Y9RPyOyn92i3LJQfa/Wz/2YNmYWISx0JKMB1zJr3NzKWdh0L
VytvsHgy9gjNk6u/I2rdQCbwLkXRZHSP7pfsvqf2JOTjik/og8/OM6dDaOUo/btaQnG8a07R6oOG
nS8mfvjUNifEnhYfApHfJuZfS2Yfl8zv3QtAO8rJf3sm965Mk8vtMqne22HMMUHaY9+bicQRr1mk
9NS8dggzhdAHIJpiRf8fWOZho+TVOp3vcmIfgNOzAINResAUa7ckAEApFEk1kl9doOqDmz6tVGgK
GEcnVS91A3cCmt955xagjAC7YnEyzkuO0Cmh74JisOjHSWIWkI+yK2zrImVwCvzGK8vZ4q6wOiDZ
o7jidQy9kADqQmCYgdBFEWE8Y2boLzDL1aSSsUsXLnsQHtHnt/SOqPrcCVgjvN8DueD8mTxH1ARU
h1hBAa010fe7zHyooXJMBYrroavf9b6uSiY8MScD5LVvEtt34g9bwn3HxFWhwITAw1gWnDPW9veM
TbpPktH63WGwwPlKbsRzVPaQzFt/9oJm3C+RvncU8kAlHqdyLs/WXCWNJ16lnO+oWq7x1Ai7KVFj
SEuANDbFvqf/ENDNWdbtLyl4iIpuLMmZrXb0dsa8QGv6Wos8GvYpFLqLzFmdGkaIBK4X4Jrcev32
DBl3qWJxoiMIARgxUR8sC3RGkovgxiUnsK1VK+1O41+lj4qftOHRxucwyWmCS87t4ftFEpe0KAEj
ttWeJ3MZF122hvZJ+UWhsDLLgLhGE8znLGmeUAFXB8Z811gBrV9UYUbaO7I3UYT7mLMN2XgBh7WB
QS0zGuWqA+yvsCsAwClrkA9scOmZ/zUj1AxR+LjD3RD3rhEQs4Xp3dng62DxeCNZVm1oIMLBfYy/
xOAwBlhrU69te+1QEUyeAPLPVM9/vYLdmRzRBLiBcW+a5tIdA40sMn3A2zPOMC/1xjY3WhTHKXcU
VR4rBSvISvJQolS/8qKaEiEP8Qt1toLmCGrMC0nSDiuR/H4lgy6FAwGc4suMMYPg3J2VzokBdjZA
7ixgMfQrGwjNmtZa0mijpdZuki9EKTuAqtoVA7hg/XEDba4uC1ONN5x/G35gnhfwjTjrhdLs4gsK
FcORxvd0xXQ4AyqYE4Z4JYgoSbxPaaAHEL+Y27wB24hlBCGrztzuUq7P2P95Wxyc8xRxibMtQRXw
PoS/ocSyCxzhXIVWyHgWq9vlybP7gEWru34+aiOsd1qu12zTRG5crYrpQYF4Y6t2WA9P7Xrguazz
kiqDL9rVEKf04IiPZighURt5fCtuMRMYPql+73bmySPbmoc0BOcwgDrx0wq9X6K2biwVEd5yydS2
+h0//70aJp9L0hAxnSEqaASesr+Mqolg4CVrbnVcxNLSiGnXEWeWXcWbixx6/NiTkrqM/RvgMHIE
OGqsyabCv3hg8vFx79PG++ozKJz3b2u3aa+/me4USaNmet6oF1m4tzrRAHpRFGI1qBQlybQkCbdP
MrzeXiis/OtFn3i8kZU2f+U2eCJLJc0OIfMn2XYvxwjNnNB5Pta2pUG+68lCKEphHrcqugHQ3u1j
8BOZZd5Cpg6R5HqdDatRQQlRp14oHSPXr92nUr6IG+B23NxLD67o5X3yCXwEeGKNS3lCppq7b6Ru
OJzZuc2acOsyv1cc5DqTbOdMusdVZlm/aZQz+t933zdPR5zLe1dQxraxMrnBdaTib8gH++O6DdZn
pkm/WcZH5I50ZjM1l7xFuouQBl3P3wgoRs3dfoFOTPMKMwGTlJfPBBB2Hq9Bsk16ECa4UVIsBQZd
gRaD8nRUmLu+P3Lifq5cGLmBI/m/N3qRr5dol7PofHhi8dlzjDcz50N1gu9/URFWju18460+ejlT
jyFD/je3eN2yR9i6xPWtt8+ZYReCEstL54VhhTiuJmeusP8LXzzL2kuEckQpsDJE+TpcrhcVYdwh
N4ruba3sgNcDGBGenUU4TsSXnARiN2wy+/ev0SL3DAxsHiVxPeo3MA5TU/GWVUpFrD2/lLQ4Qkny
AUWVHQKacDuV1/vOK7mnv9UAz6P6icOFLm+abcgH53grRWjGQfk7DVYqzRCqEsT+n/NuCwT6dYN8
MqPQgtaXwMAok/i/4l93KxxUtW+JYI2bSVnzN1eHi8DMhNbdSazTvjfBie+7FxWFAhCXQVIup3nk
pgiEzAHzdqcAee94U5DrH+VMiFG75etAjZIOBmI0lQVvIVrvTFU+7BXXWXUlXZiWAQEi0Ag0P0m7
y/JDKZyoelogjLnRKGLauOFt8tbqr0NJWbRCNQwKYgzDd4z8YSh71XaspFKzk5LJuDbMqONhVJxA
viDANu+y0xVz99rkxvJGHlgW3sVWlBZUOowD24AQsZpwawNSSn8AvvdX0oXJUopqjmLhQtFVHisn
xomhkF0nSMRBuiTisLuMyjGTF5KWno/KPpwnI32imq5MgDrRo/Wb6XhwNCcM5zB8wWBu71t998ql
wBVJjqr7HtLeQ9KInLNNGMQX4vCp6qgjwcVKFG1bjb5ICdZP8M+MKYmuAplkcWA4vx2r+uaKM1pP
9MITgIBmr1veYQAAZysb6XrHEjAnBF8on7MAmN4TwiAA84LoWplumRH6977VUNM5CS0EQ+2aWEgd
2uadxxzIDswigP+elQdS39D/Gzvo3ShMFuFGO0nRNy1EdZDODwdVFE3UpM3vy/9btePetxIgFTdb
j84NIpVjAGnEKLZuNmQq7Ss/vVqomCexYLvi9riqjq2sCQQymxcnYaHM/CLQTiumcc0fP5hHOkxG
gmp6AC0AAyi2uhl3F4tHKbtuDd1VuEXwCWZ1O5NNBgIrooSw+ke8jdnIRqZC/eGuPIADnIOfPOL9
y3A3DUbuY6ECO4WaryKuRTNdbYatEwSjCOMcTFJf0iYTSqyoZVfZ29Ln6A703GzAnnFWnSGZVKp5
vtzYE8nOARobrpPVjC4cL4TVIJq7MVPJ5ZVIs6GakmdGgd/aUjNfalwc318gvlw+TWzCg2ILYlRe
ROZnFlDNrad7GWT90qFOq2mJLYAbUrZmXSruqDgNAvf/+YVcmjYRc0NcLsuh/K4oe3Ja1MRa+bUQ
o1Qd8xmzqrGToEx3A7gpK5gCsIAy/w8iim6lSEdry4BbHWaSNd2LdGTgyf+nWDj3fKzVLEa3Fdt/
4JprGE9Dge9lCUCMq45gFElXi2WFI95n8cD5n9m7opef5fGIsnGmBH/9ErLi7hXeLogO7KrfkdDg
euLSFh6YH5OctnQOdIoUSMYRg1YkXvfFH0LM6ybYKVnY0++SsdHSbry+6iZLXbEWDOLFQJaQT94w
b0L94i2i3VUognEurHzeVjX3SgYd5JGWce6ja9K4arD8wbM5t3j6v7ji9rAtW/rxyj3whLQfuyN7
mCmmR2fIEzuzzrBj3wiu4awbE2jvWNOW26NvkgfXesugoog3+dBXLUyq8GayobCKTI5LVS1U43Kg
idFIXlSpuQsz8r8MIy2CeYJqjawz/z2DN4O9/raLyOVw/NebxZAj0s6wID1NGEGVwBcHhyfVFRcL
Ms6vamCvR5jyp4BYVkVIW22qqVTEfbsWjTvRRIGyxZlL4IQtmmG03rC/vcQ1xynS9RmmreQfAn3v
lsFOInjFZXhbWTTsyF6D+l14L2mD+8EZjB4yVnZHF76PHWeteMY5kftsjDfpheLE5QHujdLX+fpK
6SjbQJy8ketHcgLnPbIVemySNa1WZPN15cyj0zWnvvy4mJE+EVRXEwGqbmvsDqA4uYHdQ/6LTCsL
uhSvfx7gKkRIHgjI6f5x/Hd4QfiyQg4zOnqMcVXfHUXlik9E/n3Ba0YNFlrx6wj1Zt7GfGhGK2vU
ZKskY46WDbnDFWwYQB+GV1tmXQPQPjtcXDEbtRYJy9/HXOnUqeg4NqqUR+YouJjg0oUxSJKIv3DY
ynKkaDxFkhlHilH7AZOHtAeZBLKxmw5069Tx9Uz2u12qb63giN7/jAmM0keADR4m0Vm3AkKmOtzT
XHce8MoZaumpB4VRgxccL7aycJ4tYXqIWxNnQ6r6e3DngcbHIGiclaHAWGHYNAaMzsrVYaOszIIJ
QMqu0ACn15azookN2h8TvDoJWQCdSeubmYmhOUapZh47o0X/6JvKdcsbqZ2nAORGifnOsi1dejiy
NFWwemrlwX4mneUx1cTFqE98Cm6cLKkefjq/Uv1wyg54Axcgz0aadNg5N9ljv/fS5tBbXzbuUDBT
hEX7LOwOn8RusdWVSNejgWityCEzIgl/xkCrbe8B8uMMAUbfQJF9CJjeMqxPxNbsWG73unnWBSWR
scKkpQrmsBOAQS+qmXm406Zxy9o4shI57/ZeR3uiSdk3El7O/X7ynodZJRZy3/SgS9Q9HjYi87mN
OwYpnK1pDmqjpj+12VuU0BRHYNZvRyNLDnDiCR9zplEfTs6E7WiH4BKAx5pV/z/3DqCA5BQOnMQE
YjTI/c7PkknWMhqnQnBSge2kZLL3AhPr0GHLBDp0Si2cMz9cfNLfog5Xij7tZdSaWK920RJ4/0ys
qj/LJhEGR3iMVsLjaLaxG863OFB1TChpS9YTpvpg19s1PjytpIO709aVrSUelISRAvL801axldQQ
7Vvi1pfVDXB/DGH0eVGqlR66ZNR8xzHUzi3RTqpVFsujX7p8Xxkht0XiRFk4UEAmJ6PfAnmnIsUl
KOLdiXnLYc9KGH9XEO1XFC/tV/lHjVEZIl9srigwEGhG3ZxW0u80Fj3RiXOrvFaFCYzGl3lPj1bs
ZbJuAQTzEx2XwkoX1Nnul9UoTwjwcnw9Sg3ka9Kn5dV49wMkfge6PBXkrfdUhAmGhRo9/6kppoVi
T3dIqKEC0B2bQR6Bw2vdEvd9oqxKl2sxdk7SZnpKC5weHtzJgFXHXAXVVTm/TrXtsR7pcpSTMTsX
3ywV9bZuGIAZa3/zxje7WMUr3Nkiq85l3A5DhEUOUYLYHPoSOvxfQdM5N7rRBc0FGWPLAUpYGOwg
yoeQhmA5/2zEekZRr4jcJt63LmAABtRkr7IM7bKGoy+gXn9uJBgqRbj8FR133yFS6CXxjM8pv2tf
frrbHv+GK5wJuK8sP7hEUcGyUWRy3FLAIvdmXr37HqU25dz6PGKsry5qKrVdJFPuqTwCkr2CRqjz
doHJ3LnVU/eTOTpqScvYOCVPwi17X9XnU87HSFMICg5vDYERxIsI5PURS6T+XLks5fUynUfDPSzZ
+8cj9mn3E185KZJtAPiDrauzYMJ2MXFrnG948oaXnB+Bz+uhJhD1BLrNu5zEYVoEkRu+1AguxL/V
aNRVcCwa60a864+5tgmnbcyL6jhwMjDN3BLvZCodrk50Mpog+zWyWD3zwX4X+99JTVxzrWsqDtg2
/u020b2GfhxYzDf4nF+IAL1i+JjTtJ8EPezyW5Q/iAkOXLfnd3aHgcX3KqNc/KieYYF7On7Ndnyu
gkZBS5wWdeqPRFPzeegWvnjxhEKvWMCcJEXRxcRkHQuiw3kkcaBs7Xtq2GnMbNU7uEJEM0dznRLR
oq5rvBncBd/0A7/yzycf8tnJdLN2QeNPLzW1Z9DLyCxFVh8htIYUueWHfpxiPlffbXNOEn1Vr6Pb
dtKIe3/yF6wIuKiZNKf1LDMGZKxfWPTqXyTEsAvFlyELQLlfncWd5q5K/3MlhIEKmbDqGNJvN48Y
GxEXIwh4U6mzMNQZxUO8X39N3Xrm4dYuZk81MDuvhDOVNSw1VlZvexSXPwLliXKa4CHmqUqPJBvi
sweyCCFwSDc4WPGXk7em8qZ5XmE6gn0+1q2Eb+g9Q23v8GxmkX7+zXi/6kZU+BdjW5DyMWi5c6+v
OgPV/kTtEH7LnDQFQWZVXwAfLx3ZpB0NgLuHR5TYfTN8qJeUubvIo7cQJ+CTzIvzJHFxzbNWMQ1H
G6ZGmoH02N6nXEBf+N+plPAwfg7DErrXkzTJ73iwZx4bercsormoRNGm5KrjnGJZNKqzauu7/KvE
20UQTXWMOVM5pZ3EUpP4R7A0OajkhuvsuuhGMDqsMf+onwRamQe6gfSgECNnEKzUyhcgLEBRncrq
a6JQkkSP7KzW05Kt+aNhUSz9xbytEEE9uBztUVQEf8NU7rYfXisibqd2UM/B0B/kY0EDUgd91Z0H
iMpNvPQzZHOEkEBRZ5Kp5Z2jYKSQw5LB2ia1QNElysrBuG18pyhtzoF2415SkJWHPavYuYGi573N
BdZOmi52RGT3ch9EkiruBidfbfGOefPK55YyB5940YZ9znj5BNMfvqqvObA9esovXeTaumzhTw0p
AkQifYABQ49/rBwq45SlaxPgH42jCfdZSlmhVxLcoObFENhIYdCOm/bk2s0sBI0db3Sfjzuek5z4
rQMla068Kh6Gih8Rl201DLy3bkToLMDJSDW753GxnbQ2LXUCm3cpTnKCXl7wUz3o+PZSPuNOOvHD
D/00Tp80KtUQgclO7x8iIfQ8xTyjcMVwiYmYySMcxCRzNubzVz+FBuVck2PJglfoDSh5XGIrLYC2
QWr9XFnmgnD0l+YAce/lHdfwSGeZdz+JjMvHTJ85Ph80acMx8/RCgxgYhKAUN+kMlhcckPVV0V3j
hzoqXTiIeBSQix9M/+tJk1oNQv3JEW4SGHmvM464ThRSo9Gm+HGelG17f6hG7+l5AYHCcZHsjBQY
R/IqZvw7MN1KAkEk9N8cI+fh2yb314hPbVqw1g0DP20Vk8ma9EypMns5j7qXLETxuZc6Z6bCIx+Z
iyLxq/RbVOLSKqBpNq7GC1ppYlVfKo3RMsPidGz57gcdq2TNuhkChD4e68q7xhFbg3DtiE9k4EzT
4OABKAjgzdcYYg1r84VGO8clngdgRKhyTaGE7BoQ/5KUDwwiR2do0Nr5oM408aJr/LH93ahurVfT
Oi/J0cW8XRnFE1E2Sy2Sd1DYD/9XbntqJOjVXVWAO8pnasEZ0Ar3ixv7YBDB/o+xDDTmEuhFnRSK
N4KsNrUEEkztm4Ad+V823s7PKRN13ep3KtIA4SvOvsJQdVRg9GS5BtQXKyefJYFjpxIejdIeHhrz
W59MjZaOThC/zOWcpemjIpfne6tQCrpFdFi71AG0UTWMWZHLizwphk9NUtuQZH34DguLZM/oIG/e
qhKobkuDmpc/QreZjoyHlj6oEzgc1zkmYqEuYBrccXNVXXLx+2BrRXqxkM8FzBqWtp9PA9FW+REG
bnR1++F4XfRvjs96Yp5z+6Gf5iLe+aa+SDwgDe2gItoQLulcFKNty+taHGakP7D4WlTojpcxGTgc
PCXyvThiav1AAg0vYGZzZszq8Vb7YyMkPOSBAojVUQI0QtcvfJDqRompyxI+yD/Xo1qPFsVgb1jL
ZYy+NG+mwsd15di3RPjlyuQWMwMoS0mftbOXdkCyWX4fgBLx+SImnii/air/c33kor139Us0K1jy
ZHadx+hpCfLMZ+ipzJEN73hybXaHYDb5D6WSBY0OBzMJ6wyOB76E2uYMzTpfoPTEB73AQrryC95+
YDS5eI69Onhsa8ojPlMgKoNQtKTWwKBluXqzLTL9lgWHF0Iis4TiJYu9YlgQyXYo4Kei/nDgzAvY
BRyJMnPIwc/Yuf7nzVm4bcchnnUGY4Xzto9fZRWQc6iOSxmSi6IT12WlI8ljtamL3n9NZkHCsi8t
lGFAHDJF9iHLN/KykK5092scTN79kZ3FCY8JZUOrX2C3yWBsp5vFgzg27ZwWQS6v6UDyvQpQweTi
ayghe8ZXnJdi+fOhUsbITWwi6/I9RaSkYS3hLNiYzgEzx/xk0OECYmIvqyU3W338HG27A8g6JL+A
z1ltl4D7ZQ0eMIkYsQYRAJB6QvAh554La1AzOK7FVEURqKU6xuHcjBj0AjUke65gqYRRAwaac7MM
Af94lNbgRjO3MjLUvGvDeWdG1qkCZr4rNhx+UeUyWzbECk/rNnKeEy0RbPF1l2B4cvdlUEKDCdr9
Wp1Gwoo/WkB9AHDUtV75wWwNXC3QjR4F+P/CLvX8dhdzc/AUci1qyiuLS0trTpZbK2TXdAoBEc3+
iun/AS0BkekrukYLRrP895nu95j1QzPyFz7GWDZQBBTohOEeG/H3PX7QBdN09euGkANHI5tQ2qBI
uUM6WaCDLYaJ2JTSzIlhO2NwPpyyl7qYJG3+p1dmWklKyVTAyGEKzsfX7Troj9wB8E8c482GjRgO
YwUStjlzVa4RjU3cnyfo3UTJUAMjmrkNA5dUx0eKbXyjk/qd6UKhjbK2HDJmquuG/YaRyiPTRpy0
t/J/Eziz/u0886MZi3SJiwVmyCbd4WXOSkhZakER9WwkId4t22RGe5A0NaJT5w/KEl/UjuhaB/4O
LDpdp8wtLaBY+sec98ZaF49V2obtz6+Bk4LGOHePghp/frEuSe2qD3FqWk3BGhpoVQilXNHsD2tR
4gCbgLar0P2+06EOCuWPXTJG/S3U3E4OoEtcHdUiP7C8qbqClOf9f4vXMMswYGXLPxFrooWk+ftj
nxgdqYEpxnARzGpOqAv8ei76ZLZFXN1cKiVboRiwbILkBgNztbcbsfhCQtuFuugFkUYbdojoMi+m
G7FJbKKJpBDQxaC4ZA/bw51lHYexxdiEEAFwGYFN2Dkn4YHgEumIvkcRsGp0YrG1Ng1KffbsU58z
e57rwueVHOhJbz/Cqh7rFKvCRXEfWW04DrMvWFfxswpMQ7SWs5Wn5/FurV1i8S8mA/lRZ0hC2nYE
tM4znzlpAjBXcmxtagtgczQqvrBN4pBah0yqCs0NyxpRt5eZruoV4fezOdpDxIuWJd5pyjOAlJjG
u32a+949aVxg4n+5IkPfpAymanXU6G79Qxo53FTt7FD9NlyXic/vBlr8WvGSCFdNppplBIvUkN1V
fz6Qq+0ghnnCys4V9cGTzzLaSMnnoug4he04tsBGyi3sVoLnWMBlYDwBn8dqFCIpf4JXS0rZ+hOQ
ydfzLrKK+nNOwSLTrSsZVr6TVYtP9MU7qahtarpU6PLPii9Y+ljYJoy9uk0y5R6svZc5lBpSJIej
QJWGGBAUb/S/fXjKGyi8LDgY+ML4v/jpTp7TwcziVLtjv6kqJm5e0OXrSZ8UOQEp8m2ZVGDuJTev
uedIy55yt3Jyrd46j9Ti8icxMLK69k3ik6XOqxA5YZSegGsFKoQNd6HUKD8PikqkjvDzdgcv1qo7
dVHI++yzRga5L3MuZOhhynW5a6+NMZlgWEH755OB+fGSpGZgxiVCEcGVL5r2zxMmv2d9m03o+zMW
fULp/F1Bs8iaqgqG7IIn//Ya+bkvkiFLbnPmeG4u79V4QJsLPWBdvClyOTjgyuTW8kE+CPAa2y99
rDzTby9Fq0QROCN/cxCV0amyKpUwRySa348gC6PgJdpFk/9OyjTz/SXGY8w3nz1OK6rs2PmKh4Qp
ZFg4zHPQJOjE6+Yn0hR9uuTpk7kFy4UvQn4ToWUdJ/aIBtleQt2tbVM5vqpsGJWs+FHHGxlZrvQ2
s8ZnZH41PZ03W/ByoJGng7JCruaQJEu1twyd/L1vrHOV+FWTgol9chrloPvO2mteqKElOrD0SoeU
8NNho3mJAeXrpmEspmYp6oTYEIwsMqTfR0EaScZRqahVLgK/t+L/aJDzof2AesdXEWAqjZ1i0JLc
L/UfYPUWPICcQ/QAwGLuMmTOySj5pI4M8E0QdBChR+fi8YXDjWpeROrvpolUN6QfEXw12R+ybM2I
hzocDntQnw9UVlIOAl5TK5d5tVWYRSgT1vm+fHbvF0K2GgWqkHykTxuQznZaq164K1xAwafyTSmi
8ulL5f9m0Zo7329oCPt4iru73rtD1h9YgB/d/7Ee+vUjPTyqTRp0RsltVbFpcfv5HwQ5dBFtNsdC
Lwa1FnX+myM5VHLnwOvhYhX3RtBRgOj/AjlrrYHVG3OLlmZ+IoAGu59JXciHV2eLBKQtuuHu4tCw
9QY3j2UFG3nIZpmxFr9qypadxjJFVdBqW6ILZIdkzBc8MRiA8LUFQOd0do1cHp8vMf2g8A9/rpdH
+W3rfkytYfDHtxMq43MAGQiATkZIa4L95Rm0YiNnvzLA9EjP+0rTIRNH3jq8Qf6UG64d+gGyXe2n
QJOyqxr69jz2IuakV6Py2tcqpT4Z6vmV6PsobHQywrE2lAkahordyddbWjy5xrzQF2fvujTnx4cH
cJXvF2NIbtzGrRz053gbWCVAKllnmIF79dxfVGqmtaUFqQZLUhbveGF6qfLURxskfoVUsPQIi90q
2wBxXZck/Z6/dAAxnzxGSGxNBIQjEx/cc+hm4tm8DrIh5uR4KqTuliHozy8zlRZ9m3m5Axowz1z8
+22jXAKlxkTFgFkWw6PC7/sPsV2iM1S/2Y7yE3VcshohbeJ8MJz3HKVMJt2g30Jx2+xArHLBku3m
AbfWcKXPS3RpA7E1YI9pN+j0ejV1i/iISqEIr3t9RthMuQsrmTcORUBejWiefHCNtvMWSZ2SxKaR
32kLYfaH/1JY7OYzwq+Vd7sXGgCOxYUaMKLaL3YfZxRdOYJvORE3wSqaoefmBjv2AeitX4qmy+VZ
Yj4yzKtVh/R2bpZWqxL5e3yY0uamc52UpmF3/NTkw1zgpTSncAWURorL29Wwwko7KGaphmqSDTKd
O6IL8XqDBNe0k01jeij/iOwl7CnAqAkujNG+ef9sj1a/ViS9rxBGNuwB1yYmwDRoW3E1wzbaPBVt
6XwxhJsvjY1EuRB/PyOd7rXKAlEy98gbGktCNyPKHkL4FX2KUQXrEgo8tCAz/2trORh77Lks6rBM
75QQTsmKGJlvSwVV8DU/kyOATDVmjk/JstYQrWIqoJatzlxGca5+SiK+lMpobX9vbmQRz+lWDy96
NLrNYKTwW5hKKyXrH2F0dOHdyovaUu9D2wvOyCCrBbRgr92yjxNmd2O/Bs/4ioYypRivmozn/abi
pCuiboeTzbtVp2QDhVqO6zo3z3XdFj4ktbsKNjSftTGtZ+4ckn7Ctf+bVmBBAJvfiaZympYZhIPg
brOi6zlDSZ699Bk9grtB60sfQl6Zp7Or4nsEZGc8vXKj+puYZYj2yAoMaegq/+XxrMxUg9r2ijmX
bQjLD/xHrAs2ZpThRJLHx/n9Xru0E3Sz8ksI7GbUe8cbNEAeUTat++jyTwQOeJ3kyDL5CfMcuu8O
/PXa2fApa27WotQe+4x1IEmYcLJUFaxM8jIhzn8AwW4N9YQqTdSXdMqBp7xCJlCcMsdIgVqvW3ta
UAnJ0k8orfJ0mhAgJP1PubvGKKitFGE40Sc9qDHbQQLGh1xQ/7FxuUHA3F0B5lOk+lYpzVFf29qR
CfaOyifD45ESnazkLfOho4ckLbug+fhMH4fFyOzWsaFlh8x3oUSUibA++n35ej0qXorNfsmDdi2Q
sYysekEjKa6i66BeSYNRnIsKc70jP/+2YZG2Y7r/3XmuW6rB7GCvtx1OV8Wqj1EMd5i5ct6lGWHq
UhedAn1OtDwopFeRySAo2o6iMLu3GL8KraOwlqjwS+XW54+1u5ItzvlNuTc/AzPXJ38bKJUH9uAS
IVhWS/OsKNCMEkVtRKDlX6IABaukzK9mrn5hPs4VufMz/wcNyM+B5/L1kmBNEAriuc0ePOyHfShs
ZhUzHOeJviv8nD4ocS9lSi52c/pQuf6Y/CKrptL8p+p+NLsXiiFVwfQFIEX9udRiu+v0imceFUMf
KwmYwYen7yUGtgBeg8ealZJF53jNh67njMARHQ+k6eEYRQez5q3x2Pe2hRjTOWqkUCtCUeqNseCX
Ezf4o47HjfcmwRuq9jEK3jwKqepZ3ReoVHquZF9B/ITvC5FZUsBRWyQlis6KQ/0y3lBDisBDvqkj
hJgEFkw4jnIlc1uVdcFpGFr542c5cESivXTia31BV1PLYgDEqLV+kI/WskKMgq0DMVqLtzl81yx4
eOuXgyvKNKmIfT2m27fGOhtGXDFRSsBrYrPH9QoQVcZr+gf97Klp2CMWQBhTKLyrwyth09o7A2IK
7OPVJvrVrMVwMuD5MVbxyg0ZzwohXoUacWvSmyyh2XcSLfSGTglzTZuXilf59hAa8p/osXynA/8N
NTP7bEPZQ3kd2vpN1hFfm1waKePUxxSNoBqAa1iPKuRcYbxbDHgwwl69ssjyQcgrLWdzr/6qNyGD
I6mNLg3qOjXzhazMzKtb5/avBSgyL7pKO56veyljo/M+qs7Y7WXIEd233l9KICfwMtGlWT3Smna5
V9phMl4n15YuQIfQf7Cr+t8PMfJ8o441vInDWZ/5pTkBYjtNLq7cwyXi948IIuZZ6PfMBYZ3Ctbt
dyh7u9HXbPrQIR2BPelWzJfpmA1v+hGEUiPV8qvoas2pMNauSSacgbVBPA4GSOeJLG4sJFmiTz0m
AInvNz20lqO5lYbXsZKDx0QUOM8X2rhq6qbseFeLndHHfCkhxw2BC0tptSqWNScVX6MgJ7FyBYhe
/p6yFjeksU99UJEQ46o8mGEJ9hjugDPm0lYX4h3WEFFg+CeOD27N+XXF+gdbnFgIiYiFb+eVeyzL
uiHugxsNZYDApucUx2vJyxSj5ZQ8fr9AMPp/a7l+PeqSy/ojSmmnVrxODwNIt7nHHHEaSEcOScDW
YAfXPmF4+N5q69BIZ/S8f8GzZ80Z/7lx4DSx0x6Fe++/h/slPpV2d/yryo1VYENMYqsD81KjM0ey
xDSUXIGU3K+/jkHmINGeumqBi9m70Lwc1lCD/j8Do8Qrs+tklSuMo20DYSUilFUOTIgzbUZuWkeX
dVSwi2AzO9Rh/hY/+Jlhq2Lk48jI3SSDfY30KWzSmQq0fTwexIjmgslzh9FZi2pgnl/tyU8jxOdM
nU9D3CSuvx1CSn19PNL42E2BPTM/R4znYq00/B2aQzghlbf68BnxG3azEgGlnEls4NXn2dZwxVid
8szTe5FiDqdkGC+RoQ5sjlfFzmZ0fdLlke3qDSsYiBXBB92EJlU9FQzIiQ3GOSJzWOJc1X9YWe2c
FmCG29f84ZzTW2I055joFpLs0VFhMl1qCEiqc7zgBreUz6HxVdE738x84HOCqs4ol9HzBQyVlTsM
GmFwc+UsSnj4cndFsEtMIgiOtXiJ8sLuB0JvlrqI3OuSgphbDdeSUUfOr1AdI6P+RT4/pTYjOnBP
eqs/rncrnPe7O27yJ5SFjI6j9O1CEn2RFX0V8kiH9pF6gwx7E8GGoJJnDedYoKo3N4aRFvFe7Vpy
RUrqbDkcpM/CxfF2AAntq751/bvEd2a75Hapzo2sMrXptdJFpoY1iG7imZpg1udGkSt8MxglAa59
9JHAxvLc6iJ0BCzOxBVLRXm2OhmP+snx2SCznNf7Gkc7R5WRjHcoh/fDjwuh6h0Wyqtoq04+wRJK
ZW32yhbJWxJhVmX8OYbZywiIkZRAf4YqnKUUOj695ypSK20lcH9WyZ2s5fsULd2FPMx2jZDxS6dL
1uaBLIDUTVfx99MAJhKgstZv0gLum4MxK2PEv0spJPETYESiFgRXnSozwbTyR6mK2vmKg5pTunpY
Tjijsph0xzzL3heT6mZuhtDuQmiPVE6x+/9h9gztP/8wVz4/PGlidfT5EkEXcILe3SWZINKu7ur1
dZ4FaGHT2I7STyB2LbDE4wGj4VVqrK3ap54tu6i1cDyhrvieijbVYpnxFmYfDuyJxWRaKY9g+63u
OrLmVGrnS+rlnkhcvCKAV8cFUbwlNrCB3au1xs5T0zNkrUcqdKu36xUngeqd0fHCnyKf0wkhtNL9
N02PauTtAUMF58Yovmp5aFJV+cagtFY1tYihH3qMGHTVTzFBJVh472CN/edEXXSO9tIAkCOv/Ycv
EcsncLTl5bVG8tomtdkfwbRz3rBlL48WuwtrvGR3XbUS6os5tB5Fv5VHA7wYxr+Gr++SF8pGAS1K
ZUCwTzu03RY4ZUR2VcLBUknH1xd0XJS6Mm4bh3TVEqpJAprnrJLYRzz4bA1GOmVEp8TxyL2RALwY
kdndDcactrj+xwk+R3K9pgEMKOaopux8uXyP4TnXvbUQC3y4vi56iT/jFvKY/Sy+wLLAEDUwO95r
fRTqsAEiFPUeQHUyz5TZymlM/xHcM8TPQ/JOyiHCLBiOfatE17384uLpBctKAH1LMJuXXJm4flW+
9l/6Msmzij8bTvSH29o0V9125NGeKvzPQmR/D0PoL4eMKzBmLaNpO00SStWKtmV/PnSXbwOzngvz
1abZ5EDVbvXr2iv3u2XLbrJ0PEUyYuDh9wroJJmco0q+8GfAnyrg66qPybygZdQA0/VUStkSJ2Kf
EQ7P/X3SKkL5klz+mMncIf8V3mrbnXhsfTBex9u/UdibROe0h40yHkCmIOCchpupISO68eTCuIGh
jv20BjseUJtyTzcnX3RkIormRBvFoNEGdS6hrD81OMfeaftymGOxf5IxAk2QCH492wEBrwOVFtRO
LJ57kEQlsUSxrwsPVNjB99jztN3D1NNFRNMvAzVpDd+fui3zSf1CYFiRaoiyyvhvFXUkoj450nC0
0zTOLHfdyhr/Dh2OFeF7oEnk0RwOh9sOFbRTVzYk/lNygq0Ml9FgT5E7WNeJAKPlkX+8F7DvZS/F
7vj2JqYx3ShfcpSxun1om45N+gQevzAzhoZ05gPPvdhRXSSLaEUyDN8HkHZHqqZToOa4yTgMXU5b
sgCvmR9oGdiEoUUQ10dMtfwzWnANheHJr38hI/K5W4Z7lVXRPq2gmnhrpZNt1iyI7kbtPwKBXzHF
Fqoaxewrl9drEXjty/pPKblXak5sRxaFHyKrVSFgF61h6dsjyMIraCgVoYWRSyXk6iz7LFgnxScq
UV7sjJxYmamW0VJGAkC+10UAtTXOlQOALyd4k/YTeiWHxR9GIDTWZ2QfRkd0iYXIZUmTDSvxX6UW
Gy+ronnaaf+a1Dj3ETAcZdNl8tRwEbY8bk2sBDCCgoCrFhk8IZCl97ibvdJijPtIQ9NlHgcnglrg
X1QbC716O6Tni2U4xdPnvfvNMCWf86iv3XOZSLoSUlTU/B5US/NWlFhES/vrsHVV3AHZh43lqERV
vZ7eGrPc4uDOFiOIDGhgi9T0mrnJas5830UnKCK09GIH/b9J6QrPSLlPvHcqgu5MqERRN2c5haH9
g90Gu3Z0SvcmiG6jIENLt4pgpZEPH+vfteIXRVIa+dGGPsewkoyu4poXKFL9ZlVaV7bVqorQMM85
aYryEqXproMH9uvLEMULfXKOcq8S/UwEMV8Hh9dzaivjsxRQJ7kY3Ow3I7G/ihiLwvPDmZoG6CrE
UPVS1UXjF2Oo84KhLEoO/j8PX4cJvcMPjemMowdf6CK8QF5HgnEv/el3NPX4xENhQ6o5+s1fU0VN
Drz0VQctD3bYo9wNLBx7LIrQvCxUY+1OZzNSsQp2ZiHP0K0Mn3dJMsNbDC7mCW3/CTfRJNYpPiUm
NyRAmlEqVp+TGnNWSl6Fe1Yg0Z6sGCDY89CzgtgauNDt0cyGUAj6eMCEv+7oz7hIVJ20s1Nf2skt
Y/ZwGUuc4F52BeTxRxTd/S1XSf3sMvIVwCYNp4vqSK+BHaBsfUB/w3BbMfBpgglShMQCSYZXpwjw
xxpqFrwbWv8qr0c6BNU+LJ2rUPGbmU9fJk+z8eQhr2ySgbz/BbbjtnC3EhbV9ksdBZJKwX+XQ66C
XZtiP7rRvS/upGM5zOtfKL65c0NirQOGSDvbqNX4kUB/HPCxd/2CLmSzWUe996wb7p8lMn/viPvL
xW/H2fpy3zZQK606tik8xed1v3HVfB1cigi/uM2ulQkus4um7ratibVDYqx4q38p9Tgs4Egp4sRB
/Vx+2sC53eXR0g/SZdRxyZ9egnH3kh54sq6/7fsIYUavOGAC8BHRYOJefX0XFN+HMSvW9LDCzmqw
91wQA9cOM/3dSjiNMpPSk8NFTKp1pYdfXP9r2f4FflSJhIDI9G0vT1V+Z74NTxadyIz00JpvpTSW
jQTnLrSGTlIjVoAV91pYMeT+dI9SsbDj7672vRcIIvMltdWy9lGzD8/p+9mBxsgSAajSKJ2qKlou
+NRl1FK6+xMJvpbPLYF+g9e+/ZyorS1xIywrpDsbKX0EDQw09Wkx1UlY3CDVTJMcpX76Gai3tWqH
XH6AhI3AI3GdvmPgkdg3yYZY00cvRsd7DyVcXtU5LJfFJ25IE06BHl+8jrGcM0TmXGSVRMYUxGtu
YY9YlTK6dEq/owxuHdK+6zD1Vkz/bSwZfnUcPG6ToYdQIKJ7Oqf5ypRFecdGQWNUsZwrKsa9Sk3n
q2F0RFLdZq7Zy8Gm7OSG3kq8bbruVE3NuX9Tnv7LcbHWl6Ql852M/XSOU1zUN8qf3buFp8tt40Rd
5hrK/m6m/OPaYxWdNb4RKjon0l+zWtkuDv3dKwKHg7zsFruKWWtOINWx2slF4tT0aZMyJa1MM0cK
WuLMyXelxQ+tt7L0SVEL9FGfrPyZCdDngaYw2mkl2GD88EwcumEJf5NoqSpPpB0r8RF62PN8uUM3
rIVw6XMsQr8ED4Bko2nPZgM0QF5bVU/mO6R5y6tdrjL78XRNKUmLT+Uei95+kGB7kSNVIBJymi1l
I/QKrp8cwWNtiA/Owu2KFqyjJ+4rM/FoKhehQ5VL6N8eXB+qX8F9Zz8UkvGS3f0Pw+EkAK96sDRH
I28fCzM0F5KWfVPR58CTPdSaqGicmwpiMp5XfHRvzZY7Nhjc80Os4snDgst6syvQ8Si+m3eHJqz5
dMTOg9Tt4I2/gdrzI8FOtKvkb9HbhcwFgpTjs86EPX6xLbgK2WsxaSbZtlkHWhpkl4/xqQONgYG7
ldZ4Bn93avEWmKdbwtUIBSLh93JC+TsB+5+V9Hx72Dabyrt0BFi+fqS8mO73QQP7AW+x41HSD3MF
6U+Piae4SWZK7KnSuWzMf96IOUwvmjKd54u579ap6hdYO25Ig9LedaZlxJMSPXgNiQSUt+3ezUQ8
bkp2lyX21FFRdQy/ZDhDZPtox815BQ5Alfo+W3DX4fYVRRIyl3taX9kQWGO6hV7S/TlKERX1QZnn
DqgkDpSpB/i3sdgl9wFzDYuxEeNy7l3nuYIGnxmn9nUdQj0EnZPObz+UggWcyXR0sbiGQV8A8GrU
a+UHixPpQoFBR7peCJLSujFLYS+xjTdkzOlbW66rjv3sVzO3qKZ6jENfvuF6OYuJmsYeWssrChL8
+ejKgJ3Cw5BuoC7iRj4h+FpX3mB23qqvphGKkm/p67UaD/+/95+6spEmktxDTxziRuc5ari5p1ML
eJxRHDNEVy+dAeiMNXula7YD+GnRQleT9ztVGV19lkul3P3b2U3PU5It6KDYTKAHDs7QDuuTM9jM
7LRkESqD5D1DkDNDfw43ReA1/avZ5cVAvvSPCNwTUstlfg+f15IJdR/9pWUVVCb0J+Wf7NVfaGpV
QHgUMGjxUvLQedR/kCq2lZ8FnIIadq9g8Z9oWkVJ0Syue4PYbu4jO55E5WKGlD0Sr+eupMCJFuWM
8wR6LJHbbFdhpuYvOrKTEZs2l/gU7IL5esMFvuvQ+fdzWPLGczSt0Fa2HXdjFUdrFBmn6JM9S5d0
I4KmyIqAMY3R0ybcVhYBxiT4KRNbhJm8BdvUWIH9uCWLB8Mv1KA7L/EYXLlanPueC0HaVFBGKznM
DRoum+a0uR+dG8Jpnm6Vg4Rfr0lvHESoxqlTywxyVatFzuOOzWeVRdZPVLfNgOAQReQvJ8BZNkHo
RpNQNBLd4D4pHeX3coc7QqorqRy3zysPQ9f2RYpSHjPXW1tmyD5hptEeCepPjAN90W57acGAD2vr
ycbMSq2kF5WRJ+B4s7nWnjA1sTiyvf6LwuawAppYPgPdzP5UZNFeSFN0NZOAwBEfVM6Q3r8hM7pa
mntxL/LMygOB8HRJ5JQsVE6VW4kZj6EgmNI/NUGWYZI/zFcBhV5q59ZqDn4PPApmHyjHAaA9p1ex
O5JeKwSFS2W5ZKzU09y/pIe7BWH+xr0XOTYnyykvDLXxV2W9TwggtLUVbyfX4m6zJrdo9xFd9Fw8
W9zsjKleOMxVpPmG3rDymC+Gv+xJUArAZcMLC0AgZJBJP7vZXTCtrD/kHUuxywQqw+SfUmhb96kK
lj0vgcQwHazmMyWdUrrvc+b0nulOhr6L3bSZg7XUBPiqxec7hIe0ablUW2DnjjVBMqnZ0Gz3BDMA
eTbe7R7sletfrXt0SW9h6CFwKZjXvZERFF5ATBDpWRYkYjWXL3+qc9ovJCiUa40+KQ+LKqaFJKDV
gsuVbnbXXmsoRwaYSz590cQg3X6aCFTBr8HHlZcXd9rUYli/lZ5akLuO1Hz/Kg0GaO44FMZ4+AOV
EyUtY8FD+m9CQd1reUSP+1zdy/gVAY5gntWSkn2dCvG9N0FKkJfzmO76R3V1mBHGSOc3kqdRA8ea
u7/uoAfq+Bzswop2ikpxFrpx8YYdSeSyjn/c4LEZPWF2Vb44sgpywXNUO6XaSMz8Uo0kFlbFy2xJ
HIxj+xTu91Bz4hWFgoopwTwGu/MMuLgP7MhXHguc1aou6Y3hX92aMStTykjrkYfvSk+nltpoCWut
Jz7x+C7rFm0D3w3gr5z67UBLraVvMoAC+1yniCYQ3NXzg7A1aeDkJVNnmN4xcg7OpGcxwrEFTaL3
LYai3NKhLdOHVK1vAfg2hXKgWOzq6VsYHL/2FDyjK77DNxYcpQOzLQCCxcTmdo0Izs2EF5qkaaIm
ldCrH2fWRe5GDM04jVKmH7ughpLvr/TQ5p27zqPuBOheozgUWjxNwfodUtJEEfXV9aIGqgolZcjj
EPf8Sye4Rf3T3GRa6UzKusjtFgj5GYwds/ZhluX8OZ/Vl6XsiSRgDnMSv8Fn5B0qHogSEakdBKBf
L40kKbUN3GYbAcJnTzEW7bTfGGaOtpdd2zUOg4nMTcAOe3RoM+JUYZ00Fco36/neS+hgHi6eGlba
kINrU+LcNyLJ95XdvjW1NsaPY7+J8Q9eY6Qrjq0N+mGnKeskGoXFrPLU5QlQkXcSdQacU1mcleCA
tBATAwcImiNkztp1yl2vBmpaMYgjta/QxqSgO76v74kDF2W3hxJ/cgcw5zjrMnywliOGE2T3FJpH
Eamy9K+MWHi/XW+v1DbcyYp/eBfxRYaZQtc7YSKUdLIbEzER2V11ALOiiNjN94Iod3feiX/ppYE5
B+taLFa4QxvuS48LIHHeo6nrxeW7xKRfd8xeD2ELoJZU1vBTEYJ7QZiDkrXk620AFGTyVi8HRsAe
jWr6Shg6xwjiTszen/yWzzjUY84wGqKssxa0aYtvDrhVqsNwQDeNwytXgQW+vxM+UobXUu9Uunmm
qRYdYgYFFovct5RsH4d/M175O9J2oLHqWWaqGcd8PpfxMAwp6FMOtyKWCf3iKQitOTeNPVR7wbaI
kcjQaoiPhE/0mvpjR3np35T0dHZXpDQIMPDMvAM6wh1mwLw4yQUvJU2WN08sghuq7xcNmBkDQGL9
3N08opQmU1zUSdYXJut3BDHUf6R7EOugkSLfyuOcblAcZZqfdxwuyyNaqBJaLMc//FP06ON14Reh
GXsiSn8Thx5RPOqHKHgSKYIUt5IXIgGL0IB7+oO7VDPyXAd3eFrAjDCvu6Yma/mZgIXdPlCfSSvp
Z9mXYzciujHW/IglLKTbtlanh8ZkhGRNzdwnhDUiS7GxOo2NWDX49CSrqlWbdVUiR8NjP1c3Vftv
s4O02icCwWczy4E/abzoRwoAeYO4Vz1TNTEAhqHfio8V7ybbSXeAaNYb1XNr58O7apf/PupXD0st
mabmPwSRlrKB861qoVQ3dTjE/TnKY4S/ddSyAmsZNV+LPok1rRXUyIlpEYWkxQ134dtPq0UrC9ZH
7wOULW70/6M0A8822G+hoJPA+mes8bMxyaHZ8aTL5OkLCuJBK7PsHWCvZyZ1nC9cwRnqEt9FvDPz
aKIS6Y2GgiVZzxv5dF40mOPvqGJG2yz8c2RG3lcJgWcOQzbtlms/fMOEiQDYPnS8Gs+2rnVdPWqE
S8u9cr9Ij8Jo4rUSeT0+sNYonhcj//lMfXYy2sXTJ5CcsZwMN2j4qZ3XyDMHpm/hgbzq+d5D+ZKs
N7exfSL8RoaTo76s3zq3PeIlX5Xq1jBX2ILR2i9i1GWpvt8htNu/xL71c3+XrURP0uk4wLXkB5gZ
D2I/a/oWqAbSBpb5AMMAEhfZj+gQgawjEbfTe5ydJaZUCxTwuS2K4kBu0Lj06ydfwTRaFavNUFYH
zQvWabxiC5Dcg2fuFMW/kn66xJ/7kNFPTvuMvHZjxs56MNqrLgiw72I99n/B7GPJkcHSEFmq6dU0
97ka4b3AMgtHyVBlBtQNkOdg6uRz4A97C17wP57N5qFkur2euNtYOShG2Q0PZFENHv3wQtUnEUxm
fvCAzDpjJmTNR2amkYqq/UDdupjfcCeEJGZ0n035oQtII4zNCWbzidCHZck1VBF1b1rrJeLkEO2R
H4TFm6s5vz5PEvzXhPFmDpB86XdGCXX9ny+DjuAhb8fBQLAzohKOYuqoa+KQ2fnWK4eto2yxjz7Z
UpM2HP0/z4WkkQ6IhE1M4O+TevlpCoHrS28/kbc8855dQHaMRGVlEamZ4wSi2l2YCYR43epEJaCO
vUw891wBLWLnyR70xuqTuDzPdqbeMoiQx1owNK9xCNnXKLXxmWmL7BgX7NbPTgsJPKahFl3yGzvv
DwR/LQp6sMXRhhjyADqhi1/Ma6SksnGfs1H5J+fybpaaWITZmmxh/ZvFKf8xmYE1SVB1XiTkkY2i
TSEfjbuoBgU0gNhQvKy9LcZIC33E+VD2oF/sQEoA43jWESiRXb5rjJxof+w5K6dVvYV3dvSNUn+8
7ynC+QoDLCWxBZowL0Uold7wUjTHMAEUWKChFGKWvS+pLhHp2SUygB6F8myEVoZnHHDE+eYw1fyK
HPEDmPoVgAXn1tvGCO6M93jUfAxJuH1UDEHZ9SdB9aeTWPLfyjz7lZ9j9ELMg10WHRMc8ReIhV+1
FGvWVaeUzkgHlyqNzboHBREqoZTM8d4j01K1OBMxiyYIsNcc/NDZcXuLeVnCieHXP9u3o9ljgC3B
KAxiPrQDnORMLNwpqRFipEeMBthiBAgZn83h18UrMah56zWwMXo/CVWM9Dp4UDWt9YfEcLjAU91P
/8qW9sIqSxTLtz7VS+04a2LGubEOrv58iCjTUAfkIujnKVZY1SglhQC29t5XZsvYRruSLI8XweEY
HuZkclCyxjELq0EILGowKCtaIAnncEV/OZS1E7/a+3HwM3F9S2hb6PSqmN8e3ixa8xktXwsXi23i
s1B74XzLcu5miObmKECV8WMEB/DXMskWwiGyWsc55ibG5sCAWO9c2OsU8jvgwOIsXWWqeEXT4Uia
YoD6NCQSLlhkxEPg5BRJBOqX4BeiSaqbxu/WPy2f3dV9jU7gf+r55H4J3LaMRa1WwxcDPgJRM+rB
1b0h9E8Wqr+Tm7qs0EzD0bpc1aPTYbyWdSnDuX76NaG7BvFgt8JeXA/29x8ZCZfuHV3cMufB9JJ4
y2JW9lfiyTpTyHO7GkrsEusBuNYzac8LLUEuXlrlt1US1hh+/bwS2ntD1XlE7/j4WW6ixUANwFov
gU16X/TTsEX59Anj2YPEHl10Kw1+coDsqqX1yCygNVL5ruXlsBWseCfkvL2+0RpW+FgBjA6ME7Za
Hy7zP7NF8NuKouyxzy4yyP70b+a3OxAVe4n4srmHjTojknb2qWsh/ODv2U2INbNA7WLL4ddExg0F
2FhFWJiKGxbs2MhNoZudMNIPfGefvUnTzgQulNbC1XoMG/0LgmYi8uW+4aPif87ULNYUb1xqSAHQ
8uPU5IsMq1PzSJP4eIvgFSAYXV8WoJrm6ZH7Z0EXwq3kpJiq90PlVm9cbJf4LPjiUp44Q0MEIalO
YFmXLW41SkRTU4D5fNZVGiAYguRWILLe4A1bk0CfoMRS1EX2cRgGr5cbzJ6+RXTBN04bUuti3H3g
fy/yP9ZGhcTRDujxP0oAphm6FKxf0+U3ePyOvHdd/xrpcHnfFZt8flmPlZfLi6zqtygx/I/nl2jn
wwkvF/TLa12r2htQ9jxhGP9MR8Fcs/r/OHsC+nqp9eSnZi879IlEm0BaKfYCNLFMqi0jaVppRuId
h5U7ZiSSoHeTRl/k961GKpFlqvn8neYcFOF1oB5iK2w3EaKuFeAfICQ3L39FCQ1DrfC6l9Xeng+Y
SZwZIk5kMyWG5t9GRxeVLlGnDakrxn+ZDHUlEF8s+ibrwb3dARby3NS0D8MRnMrdDg35dZTIUfq7
sH6CdKelLLlRMZr6GYz6HXKJMnA2WPIIZEEv45CQURQ0l5p4PScj3pWHiKWgg4r8KNxSLfSB63MA
Ge/EKyIkTX/6NZX5ihV43q72R18NgUzVNDx4CU+nvDhU4BMquLfcLj8e9oxiG/FWJpY3jUz6sMrC
0e486YX3O+hWapyi5ipIghRGX2jHjK7qPbuVRjRYxb9/XPO8pkXLUBxiVHLKxltHmURybjRKc7wL
3N60LDDfdT8uHzzt1oSm4gDaWFR4OtLunHnWhTaM7kywqWbQHXTa4QL+S35xRucRninlWGF4fKNY
02Kd7RSbrOlqNHz9RkZnfFdmEQbus9OP+R/8w61N/5nIxut4CnzIicqK1bilVLNnR+rWANwQ+Hwm
ozI2oY6r4jYuY2jS+1O8LAKOftbsyNQGlm6ZTtI8ZZ1ohsMnwPhjf4LvziyqOXWnoHg3+dUyLsw5
tvp54wzi7pO+7U7P+BJzgDmwic2nsGTtXn2+rBYW+lpAe3RPTX48pNuycc8UPb4KgpnL9+eWvRaA
HlSqHhHo0k5mwDqLS3TmzjbtVK0vawFik7KlxW1yKDKZWASdOuWu0JtWomwzoW67Bz9oL+Gylm9u
6gfk3OMcfsQrrQ5lhVV4YMDEK5Un/M+6OJLq1XlBmeOsullTNW95s/yrT8t2IV8xmPFXm5j/9SRH
+eF6O9Sks+uKIXQcB/KYRwHJosWKNasQBQsKXj/EwRBum+zKi13yZoyIcnGaPJuNd5jnhgcLC9zH
34BUMElWc7B4gWniEHVtFu0lj6pbTcM2QlS4mFb5Wxbb35/oS6p5tIWY2pfomS4cbba7siej+zPF
TnKxt2uHGOqgRByNeKDm+t/03TPiPhmFktsEqSL0CbJw+qKGIjNphRJaftHKlyM/a9EPE72qP4mS
YWpbIpqPy9RtEtrU5mvWZCeZJ3PAntCxKZiDzRhD3iZjfr/plgeBOB1YucsWl83SxcPnnLm0U8a5
vny1bI7cCZBZOfA+nQqXNCGS/vqo6cZgnhVuBxqjPhwuvJmWkseToPU7a5BJspPEnkG5kc4Z8xx6
BM2zeINb0XphJjE7ZYVi5dwtgqshpU5lp759deHF70fdc7Ci1EmlQVNvS+szcjK4M0GMyHqy+8OG
VcfUonhQq+oyPHA3X4sCoevxuMtksJhfJV4ySGUHcOhasfwrhzMFbj3TPiGnyz6FxcPkj1224vsv
da6vVepmaRHKNyV9iT0Ytg8Al+9Ah5Ie01wOGXeBIoaK0N0LPXIQf8AbRcipFZ1bVWyAmyvmLEdi
Amsq9bF9NeJUe+4fPuQCgKPKDS8eKh8xYbP+TBGQ98XVsU1a3wmK6uhBS3H5BtNJZlAiQgTbV3iH
8Uhh/tSPckQ1qsD2Yj3KaVbrE6/9FIQjY6hz2/zboefW0ThmIFGZYjhPkJkgAinOozbvpUMJIOS5
Nri6FjK5WLBBKZLknJv8ewanjF265POuQtT7NOF74eI6/aUReHxlK4jopjIZFjzpGpfbZD1cH3OC
sYi/W2fC3EOGMFprdhVtdGGOjo+Jb7ObKCo4Tv6zg1mqXg3vD08zrZyCLGsKm62wwgqN1Gn7ds7c
SOGWZ7rvbTwyzvQrkqHNTwy8MwCf4M/XktUXisRNnl/UHx4cHRUX4UTb0qRk2jRdfir443eo/CM8
ALbCd2HMJFbPyUhzEu+0TRWxMbKDT2Te9AKs6NH0IIH7i4kkXQY2jEMlHKZcb0sw59MseBRK+8+B
aiGbhJqQQ0Ypv3aamiZXA6LtiKlJyq9eb66PMtsmx9CliOD37ZslECYwecQUpjX+02jAv3T5MGcm
UKOcoiuC9sCkqODMrdiivIISVXRfGJ9/WKZZNxJB3BUWqUxLClV3zKZlWJr42U1kTfvXe1pNtMZ9
c0Im/mYmRCCXGHZATuAfL3CzoRo5Ql880nvawzqj6n0E0RtpfI4hXw/3DXZD6Z3OcOPAMHYFMgWn
IysB5NdEgWOcaQWiwD38CvAgnJr0FHR7q0CzL9aQ6AJFwi65pXoRRtsuq2fO6TBOdVn9s7ErgKea
aBYg1ry23ClhHHzCBpxiKLSoJ3uWx3c94pyfeuNEHToPmyu1MQwdpiC46qXNyn3zC3FnkL4vweJN
zuufhPbDUULuBkfu+Ldw74hRhwckKoLvZE8KkK85lcjUQyREqFbXKKJPiSEI52nCeA1IHWMLMAnN
RmgU65pTFFYcEoTcKKg+QzkG/JP61wapn9COFFGbszNLlgFA6obT+KBVIv6baSZM+mRM6fhJ0qiC
cSA2ESIISS329S8uf7TC3yLcXyy9EUsmo5Yf57S4uyQ9BPcBveve7i7/NWCOtSpnl01S6xGiekgb
hwTibyTHGFO5g+h6o5oDbCdu0H5/zITAf7pNKtCC+x2rm7aYhV7MJZdlTWTfgWpy+LNUflyZ7yQk
H0G3QKrJyUXaTc00IH0Qwm42X6QvxR64eVqnbIeCzbhLLWRHynyUIXP95V+YwHG8EGQTTVNJ3E21
WBodW/k81hihxmLwUtv/2QJyPTZddpITriOCq2KGek16EGZm+e1tyC0plSQw5JIC9768XdnZYpRm
6stWAraSloLDTy4enJy9z0FrzgKCzMvJZ8xH+uJPwbKYWEeWg1jRLdVzeJOazFZx1G9mNePQ8+hp
nqyGAYl1r02Yt6SWprPg192qGMY3DaX3VILpPtDYtyS5UxN+yy4oAg/aSNOOEHO6lC1WflQ1Lm3f
EzJBhfFfDlUsbYnCHT8OIZ0nWjRd1v+yvEpHnKpGHoW9fasHEtYJwshYQsKaKvc+0VeaVBal2VlR
UJggJXiqH/Qpu1jOC2W5RJoIX8vgvAOlt6iYyvzNEhym6j3Qam3cddXZE7vpMpoZU0EhsppLScQB
mH3zQVvv5VhlcNroaug8YNKMTwmPpAjzaIcar96TNsp06i3KZ7RILV6iYhT8/BSEJNi1Tkvb23K5
ZBiMl3CfKBHC0R777eskxTXn2hvZ6s+cFfvZ4p30UmW3sLjUwRhdvjVVbc0A2GlrbHRU75dFmKa+
DAFbMtzIOHJbbavDW6T/oGm/SX+/sjYGl1MaPtcEEkBojnlTSbLPZqyU84LzGZDByEBOTzJSw5Jh
63JC1wVm6UM2NOxCx1I0z7l41Nm2WDQCmZ+bGSpBc0TckDeZvaUllExpZv2ga/al5XBIvNJsV5Ny
GUufyaKBQJAPzLDJ4P1TjsTl+jkbQGk/x05VRZL4yLyzLIKGTAye8mTWXiV5i7G7S5amhK4FqY9w
VPJlKiy97EJ38K6W5vc6wfuqwNuBPgMlZdiaGFbycrkdIHXTNm9vzA1dQYiJPmCcU4P4FnUPlKw6
Am/S4TOwNwmWoQGG2x0k/kmMttfl6MkbHFmC9lcFbC1KA1CnsEMWIyW8AH5w/8m3nUsmRKlcarwW
kq6Z7N1Gscb6KkIRiZHvmGp2QXJSWAnCsJ5/qoL9ywr/W7zSaAQziK29Ay3IuYJ03dury/+I0Hdc
8qBsgdXAjDMrKsUNf5L6PyCS+Cg/SOr4jual3IUjG8Gyx3pcie4m5hWxngjnMRuOi8umHLjagVcT
sRiOAY6Edx8qMNmxjbCQB37evtIFCWaRUow0ss2/k3YBnWCRN1CdNpsAEg+5OFMVqZfK38U8RrY6
Pu91wU11odKm0QAZ0KRjlDv0BTZ68VdnDe6jgZ+qYz74Lr/Lk0p55jSxBM58bU2rLIPjfdXVZyhb
ZNqL6mE2e2l2m5HXOGx+drQC+3OaQEa6HFiIbH4Y6wo3Dakar2FbvkFg9fYEJA74DNfgOP1BmyJd
//gAwTqDJcQIUtAKcQ5zOcTV6D+chg0b6oZAXOZL9PVAfPAsGqCPYzntW7bZJeGld/NVUi+1EMtr
29yZWkeI03eRydkayM2Lg/117q5hph2YpfCSbqi8t+oncY7dvNkr2pXkRjDwezRV7P4AkNkq43a3
73hi5XqV8HOc5Uop7om+ElQEtmzgP+uEVQ31+KdWMgp5faGjgpvlV2bTlqI+YSy9i+EUs4bE+rg0
aI8QgZ2ifAg3UDUS1YJATL3mMQrJwcOytVSBePSZFXTTBWti0zJptmU2ykSlr1xn12SsJthyDohY
4b0IlLrPjsamUgI+rDD9MoFe875OhCMqDKZYYFDcZCEiG1WOLWlwfeA6bTgMFA23amCaV2IPiVRm
abdr+iqWIP4oJgenJwov6dxRNO1ow0N5f2p5GEpNd+NmDfK9XwGkWnfs1VMMjS0pdhPU7OOq5g9Z
E7HuHhfx60VrDhiD2/z3zGj+/3/+bCU5JijVp3UD9ImK0Lbj2QNnb2Hskp0K5rOV6wCoqu2AQnX/
Ves0lHVSvjOo5MZKxOxfhIFBbbv9Wlk5Ci2mDw9nvy5dgKXpV1a2fsSj6L+bpX4pmh5DcSAHSjs/
sdow6epAkExG1bXutiJKvPhruLAO8O4mrMoPfHSxrG7nfN+6uRbLzyiOjvDx0q98iDrPf2Zz2g1I
icxHUnjX/8IUW9IUKnLFYnsDmwfCTa9qFDEKQ99YIFkv2uMmr7bqEiK5PphXxKv4coNzibqc6+us
/QSqLe+FT8WCvYuIhqjbYKIv545AFDLQDELuPZ2IFG6neuJ/M/82xUxwJyDoLkYQFYwwzoUIzF9t
NiG1Cwvt0YndY1TRPE8HtY/MRN30imtRTz6krkdvzzwyndDdPn6c23Pq8K6RVsCqpgdAbuBhQkte
cR1SHfCWyGsCBvXcyN9T13yVOO4Yx7O5ZDGmzph6L8IN5CfsXxtj0e8KAj1LkTPqrEKn2pGSxfKD
jQMpYvOubD8P38dQeIYwiDNWutKBUzgGzG/IP555MXLojfpe1uztgV0jMNWeqIVR4b5G8kwG7+Qk
TggtjZgmN8JxRWuNTchuGOpsPn6Tmb3EsYcf2bquF/clKs7W7ID33teTMUH+pvokIj8kXLyRVE4v
hb4Q6Z8iuET89HFo4DtuqE77nYhNjy/RDvRqzFwmvXUqb06RiTTML0H3KF8yEQXYwvEI1SL/o0JI
ILisYh1pTmKPdr8VXIO5oBxTDtxOOokhhgY/7PkXYJjvGGorvTiVWK2qvqzoMLQnxgp3RaC+hy6h
zCRM4HZPclxQZWi56BDvLgVId7fCZRHp9Uwlc4e0SXwgT7HHGV5CcG3z6lTWX3wmj03t2AMdQCbl
uRF5hFe6FuQXgd2HUxNYbafSFdY9v/4JVgc7ZDvc/JFnJvd/Rwg4hp47v7TRLeIE6RiJA+Z4z4yP
/QGYQsS4m95XB/WUcIaXinVdk6fJbPSvnAQLD+EYpLU/OPQO4QiRjcOC6HEJWmLuvwte+GI42Kde
mNy3FqZrlURdlHYiX0NzxqGrR+8GqywHUYCUD6LxRopaRNd77L5IhyFb7N6mjc9g0AYT3XqYI6aM
u75nrikcOlV0PDRibbsOb9AfotZ2gL/upBGSFGrqTdHsePILVgDdpIurtOF0pAfYd+w0DKfxWE/B
WisqWRZH5Uwf2iDgq+ZIJx86ZLreOGyk4P9GNBSNhRNFaT+QEs9+e3Hk/oFQKl0lNxRuzySXIMeF
wZUM1AHZJSQv2G/ilcirBOhWhPvfL+GxusJhdOynzY/unMalMn2dJEvN4isl2XX+FAUWU5QxbnPN
g35+dwxX7SAIQSUa+H+Q/hZOCSRGJ5hjMZJJheG4Pr63OtG7GXdn5FL/BPM+IT0eDmRehyQ9+aXR
ia1a/skt3kX1qjtxks0RBawCPGjSaIrMMTj7Ql8yJEuOFwe2cCmxCbpx4HXoNz76yp4yQ8qV73LW
KRKmDwfNKfXk0yQSlIsVdpmDmEozRQufzXVv07Rnf3KKJ+Y0r4OlmKedthuWPgwnH1P2uf6HprIb
Bc/IlJzMaU29N4khhtR3LNmKZb5d0bTqv2552xNKhRlUlFVW4W6svbG4YPEzd+Ps8ehoOnRcwqPT
9KSs48gJ78lunR2ELK8YIy4r6BWtcfp7orNQWHJ5lClbJmnDTUwOidxfPEmcbYke1/GVSBFoCL9B
Dpg/SxNGHQ9HNaJlPFeydVRgjXHCU2AupdRWF9vZnhoSJhzXldCbZMRN2AkTrI7s+I+6OpIzaqk/
upgA+B0kAIcCrtAh6fZXs0jfyTE9nLQ8YNXR5Q2HmPUCHXqopmFSd2FVaK2IkPtaUXSqTP6+5iFe
7w8QWhrg/4YfKujDeKSSjZl2SmPnD8MyWfjGPh6/UM7EDKZ9LQTNB6u18Ebl5/tICoNHb/1rV3QE
HXUgS7CjPgCI/nxJ7B/wJN12HguciM8SK82Z+3ICk4OHYG0pu6ZUQetirS28ZiF5xtD7Y1qHd+Id
2nh++jUqpvSIiP5YtMw1mUsdBNJRLGs1DayMN5G4+26rBMgFU+rstsZQ83AWThFnns+wbmnGxyn4
HwFNuUIXur53b4RFoy4ArAsuyFuNq4ukrcKwTfRXPKZuX7FNhgnkpfCJFZRwbVBn8I5VKcKQT90u
ixk1HU0hk4m6cCiJq3kfVxHxYprqsi/sazWxRryBJuh1UegeH1rBvnIkcJMl7JKcuCiBitj7uaxP
iTiv/ezBmws1GNWpVk3CdOmp3DA7Zz+5Reu9ib0TWo3oI7wBQcIYPYLJLZgo2DU+AICMQ9TKJcBs
N7TGNYTU0A4QWO91dAQzZP5vNuXAQ1faBwlY+HIcEtqYwNFjFfeqD/w1RzIQx0uG39o3w7ulTc/6
kZD/Y3ivsRNrKRY0882JwXXZIa8Kty9wvaqoZCq8Ig078xZeKZxJ303doFUyWHfNaz0Y68Q0//VR
uhwOX8/9czACNC2nhngELOEpPthA06TP7B0ltAMbdwYm1c8dJnc18bLmGL2a8wpnXWOZ8sR2YG9D
8BPSrbbOXL6lQ5MGfgTe/1XdXaKTP4NvJxzY4Bu/C2OlU8DLXq6Zyk/kgUPRCXDi974N1Ik+ZPoU
lo1914vtLTKCwy7v58Uy6J7qV+vrh8d3ngiVTG8ZWruEMNH+wXif181GdJ78IJW5AoZInHRHf83e
vLbE297cWLB2x6QbMcyTXJxqv/g/5j0WpiXeeZ6pUQqLwgIzdVYlFKS/PqwTz6u/7A+VLbYVAJdJ
C0CIlb538BU0JvII27F/IuNYEosBFbFYVPtGgJjj9w4zksoqyf3zaxbNO/UbwfpbGQ7+KRIgiF5b
QBSdeQs7EuS95jsqxaF5MYsMn6NEYRHal7vWi7DyCsS5MJGyxCoM1SM3aUcyZAzvJJneEipqeDPC
Dh/SFCNJGI577lspXhFF4gtJfk+gL/SF+1JfQLAWNBU/5eRDJdUlwviBsYsAtiyrOluK0E+sdMKi
xHDCvL6EqNMpfPqsPKnNf9V4q/TnBWog46ogxla+6ymcBhgDsf8HMLqU6Y0cyY31ewSohAr9CcxU
aYZXdTNuIt1YWBIjrl6XN+XNYM+bZ1X7lUtRFo3LBMiHvGKi1EqpJ23/Lin/5kSAN4XaJKyxjUCk
Z91NAxc6vI961qoGGVz4gVcSiQFKGWey4yHdjPK/LsZ6dn8YX8l4bv6pRvgsq3hpHlKNrYAYXfen
Fz8Ea6SZ8MM+Vaa8mUmRBy5Sr5B7xr/w58ICtGUlqjvOHKJFZTBZ9M0Ep4HiWBWY3S9Tj2BmnrZk
DGX7s8k187LOAnkMZkXCbmtK+o4457ThgCgMInVUAZBv/1sWreSyHEXXdm9YVH/yyp3F3HkAZNDo
u3hRilwPmREj7XGqoq34o9GwcQ7dbnDfLgIzwVRsSuseE0TX1B4xG9Ar/8zFc4hyB7ITMVkesrgu
JtYtMrwgxkBcW+sjEcDO7QYRky1qohSw/nzlkeHs8mE7Cge7mFT8UvmKBVq0gbw7/aXiCsljSnQc
RlEQesMowwWYXY/VW2cRWNg+MNtxyk4LT7dnsCVuyKVTt3d2t0zACFrqoe3C9oJoibVy/PuDithB
/jxidKSAdNNrI5cvHM4+FPQjm70XljRXKnRmeFDgc9L3TRxyoNr3kUsfo/a+Zz0VEo+S1pKq0W8J
R0juNI6mMuD65qU+p0fC5PRPykB5p/582F+qbgrEMUXj7IL5H81CBcVnFiGJHnA/S/myQhmUko0v
751sgkMYzxRGYPIxxc735n76JkXtxnTjcBgQ+Vzd1kJO0u2/qb881ZO1oIFQt28ErFANrzJ5WB74
9H1Wt9JV61PxNB5h5jHd5tVgJPE1EDZh2M19r46WO84IYsT4ap76k8CmgZ+MEWVo9o7zMFAppwTf
MBs7KslEKHteUofjVuEIccbunBg8elHTF6hginjdmq2pM8P19qNLeGO/MuU2oXMYBnoGOQo4z//G
qsyPYrCZXJU2ThwJNi8k25gzuXZNxhwqkmuilE8JhK9JCot3SmLusZSqWXadEr4YiMb0bbUJ5wg8
cVqjKL9BH4H1VvAFAx6m+mlJO1dBCvaQSeVdDWD+wUVYf8fC/vVDUXwdSGNvpBD0CFblLxT4T2hv
i+xjD03lzvG6UxJvk92kWFcJKsoraI4Au4I/pa22/S7dtPofH/TpD0Y150Q6L/Zb1dXXuV8gIKN2
Q857e6qhLIhuv/V19q6asmDNnOpranOvPldCylq3mDs/7bem4wkM6oCg+iC2FAy55yHk2ZZkbJ//
lxl1usgvp2qTvbvl3NHXNZMfunCCzGGltfTD/eL0Sjfmy6ax6S5T7i/az9Bd0CkdPk8mdhCpfCrk
JcywKTCnJ86ZdaZODwdjY2xLYwc6PI/NIxcKmppUbxlNV1ID3u9jY/HK7cg2ORW2WNAn8sPHJm8T
Fc+4u0h/cdn6BKUGkDBp/F79znv9OhSBXn/XnjKH68EkkNV3eQfC4yVBNe2Klgt8Fpj/ilaAgwIj
jL65RIufUvJ/Z3g92ymeZr8z3+R3/eC7fv6UV+Eg1WDpao/xr69YWOMXA58H8OQAuztUIVGqxXIY
WndyDq1j9zwAoy/TpFmEltbvzJr01KD5G8+UiWlay+Pjh64NGQ2YGCL56YhP8QJxb1tZ10KfM9/g
9PU/SbbA+beUoyCmRObNhWjIxMq83n2MNMHnI3xx/w4S96i97l20pJe+I3qBfb6/+GnAvj/H4fRZ
dUZTvAwIQW1fnPcVOmR6y9HB4otxPdGtSgQx7FW1yb3MaAeiGtORuarAu4606q93mwL01n8Hgdc8
yhEFt1ww9NSUeSAkz7o8wX44FSQXMFreiwhD9av5qhD4VGPtkHWw3w9SHynmj4RLwK1Kqh77ETmD
X0uhJcu0NT3HGxc6610pQ9G/xv3Fy7rrJH6qFe6iXv66zrJ4+VehNlkx00QJGzVL7/oQVWofZ8yd
/NlaqptWMjxeZOwj3sapuakQA8dqrEWO+tIdi8EXpiSDrwm3BDy1BThWWBNUQSSF4D54XE4WAw6y
Uh6029PLoTvvJ6vVHLVw9CP+S/6M7jDc1MUV1/PklW07N8emJLma2dIeAfO2Lv9tBeSvYp0V+n8j
ihahcuD/gAaFWiXcBt7vkuTa6S7Aiwvmq7NduFojLVakB9LFizXBBplxXSZ2damTxqR6YNxTtowp
m49iBaRhd0O8XHzFYXI5JpmJbuClDQLe/CWA/uHN7ndhmkcv8r51NQ+86jTBhofi5l0UEDniemen
0bAWvTV4Ml15y46SyIlgjemjF4ca/cG+oMVgiecDGGTVj76AeRjY+qVf1O9+/Wgis2b+yihM78fJ
WR/DG1h/wxqxVBxO1sOttJ+OutE5FurrqOPp+d7EEhjLzrKMi/X66ysOuuUaOfWl/0C05KcG3qEa
tTjeLBs/DcQleNm9otn79srTD9+jVt89SiGByipgng9fGFyqwGXslj8ducXTHKehULXhMu2mRU4x
g6x+biZSXfNxc9vSu7tfl6jb1OOi6qpdAaYE5yzKISkh4eYVeoOZKDbyNGegOkxqklc/BHWPF4m9
sYJsWCZeW3k5mIPCeuFbKhehSXPDhi4ORTMf2op6xtGsHpCDXumkwM6Ao0XMLIBG2uAYqt2SmHA1
xyakiQ8kEAL+hKV4154YRytmzJurnQFSkvVBVIXzcAClC8GeT4PhcZUp0MhVsnIXFKH1quYDjech
ZgO+ExojczGRyO26h25llgCnwCUETjPH36PAM9D6FxPzuxYV6my9aE8XEY2D+QIegzV9N2JS7cwP
IY7WJe2tNwp4lK9wrRYcXiHs5qzdp/E/sMzzkGGdVbjA69sj/cmhS4C9B0lf0n6qdePLkPGUO6hV
Kdiqzlu4Uz4y+bBqk/7UTjXZyrlv9H5yPScmjIM5VAN1OjtMwK+to8UlPcimdNp9VtyAWA3Stmkm
DzL6CsO2il0QirHW3Pz760NMtIfALfOuoUiXX8Um1aRNpwsr3HSukO68XrTPLvSslOflbkWdgQ2+
HiUUwDLaIG8zSCaM7aRP+7wUUbSp1Zz8a2a+21do1MgJnVApr6eTTHpWsw4z0CJCfVoAJPKuGkwh
16T4MgQQfktpXWvulgIaUuHAN/5vkIdOXuIq8zT73m7IX/sUwRmg9HBM6vwZjY2iKYYaItYDfOMQ
XJnCPqAurfoXdpGrrvEViiAliBwOlLKndue1HaXsFasv27l/nlNk26dfNLPsplpCxcWImaaCSoSK
3xbLzBFmu0jbavfNfC/JAIEow00p+M7eCb3NrbqGOlem9cWGQNf3kz1bpnorHJqwMtGoHuqKIFjm
RcF8R6dxONR5nDJ/36v0aYL5mUCgCG0+31+GOSxmvTldOxkomxEm+9X+2r3h5lD3ANfDcpINjDEA
xMz5F52I+VmL2GuW7L62tLEIn8wtltTF8i9Ab8bRoSBUOeIeLYY4c/LyFK5cCrOUwpZSNzTt7aIy
FKCN3Wu8w7Q7yDvaaupDKGGmH9romHmq83HyZvcWoCIpGRDBxphLocfxgPsRYMoxZEJxopJEGXU9
Jp8Ze3D3c9Zcf3siU0R2YSzWxsH4VDqZoeZ3FobaGdL0I3Sxvu5XiYt5R3TXLgOvB6PvS0NEO6gy
rteL5P0hCWyhXbvLj135P+ux7RXCFPUIInZCRrehbqH+avsthxXLCwU3sCwKA8ULLuEbElHcyFzt
ILKD3JdONBC+TmRM0XZV9XGdKp5uJDca8Zplw1g6h5is2WOgnhWnL06FuEpmogMbOAbPWfFghu51
i5URNF1Wd0a57Lmb/TtElvBy9gaL8dJqvVgvTOfcwFZjJvcsF0ZPrVdJB+tIFcDefluu1HyPYVUg
uEWjGfAqc++hFTZXzG7l8Bo94ebYnXOtujvYy2S8ATxPZOZ9ETJW4h1wfV+p2yVYFNjclNrtItRV
WIQVr1Np8VI4xU4vjqrZmMMd5Qx5c98nlkMiO0p3lgT9oSWvnRZ9n2jOhyaGEO+nJDKKHhvORSwK
OFyvIGrY7L4hjd8P5/3zGxfGDLs8HziL745z/8GLVYhExmEEszZQ/kcM48frF+auT7o9c9aNYMXq
Sd4oP9dlKK/2UqUM9lwECZhEMHC0gmfwe7YCsBCP5Z6KNOSWi5ckhSAYSlajfp8OHzexQ9f0zKlq
CUbmVejfeWH9Yo0pBwKgaanvFih52Q4hpGgRqxTHSKx7KvY2EAAHAd8WNXYh24F1zNYnOCqy68Bt
IOG3yPkjpjF4udXD3ued8DfCFn5FkDIjs4F/a2G6hre6E4khkKP1CL0XKjT19UmMM84U2u3c8fRZ
EAPnFbtnIsIENzYo6++jbGV4Dr8pIxwCwKX8dlTrU6PwxwpvQgAXoYJbk3OyxCbAJYVNN8117AI2
FU9pKMbPvBJ68qFfp4k1gBsEZBLAZAMPbK6atAUBWI7NPpH1UwQTgszLr8OX5BcK7ANnxoPiqaLi
KFMvT3ooFIxPLsxhA2IjmLNR+acZZQAZAmZx/gyikkW+zAFsAA8NB+M+9SK8PFqojAa7dC5tDjer
/HQuEHvcVWV5G20jmtmSY3KXLlIQkXGLCmHoiNMgC4/qSqbZKnaJeRw3Va2f8Qv08iytpMUsTeyB
uXIoLvFW5tgpoJQjrp9oMRP9JfGcpFg0ODrKe64B7w4kHdFd4D7pFdWO8fEx/xb4J6d2WkAa6wvo
/6bsm8w4dZphhWB/kgEq2KRnsHrmSbj+O2nB1xMm9KngIUHcI0c6CB/uV17bYLc2QLYz7Grt8jdG
BrprFznmzzalq/z6IzuAS4yHW4w+wnVbH2BnTfXFV0XVSNrGDygrOv1Faw6gSouG4olCBB5euVa0
La3s/RNI+NB9SRV+L7OSihlR1WgrzUhzUTRd14FzHtz4pPvAWu3PPuH7/uRNZkmJhMDyOaov6kAE
j6/DcNRdc9uBVHrS7pMAT3/hxJwNYQ2uz18vjUAps5V4sBrjgtrkfxSaHM5n30oBhSikieAaA2xF
DqrGTxP+mSXPMoCGdaUgiMseR2slc7yi5m3itaNO+4rKnjcC2L3xejSqIQzQrUME9m9QlvcYhvAU
oAhDMsm1GHNNNiPHL8gGPfyovWkpGu6gna+W6vfu2w/d1ku1HJRI64m8BZ4NqRxunIwSxAzHrPb0
63/8rcAFbGYNomEBWaMCqCbMftfInWkBB86m1DDKrR7R0amIzoWmxH0jlijMKbxNP5eJU1J7FYCU
XxEY5yJvN+MLlj4bflZ2ymbvPKDpNu6rOL/KtfwhXcFmIvDiv5yXKiNFqmn1sn05B1LiJMZwtSf1
HfaZmUBhoABdkdFJHIslso/CMItRxmvvvadmURLpg5Bf5eaykWJYA0OgHjNopc+66l+K/09+XJW3
y/0wPxfhUcKNKURyMf56izPRUizHuZXLrvsREwN3e/4IMXjbaqTcYnKWCtRf/AXVNuDkmkJ0MNIr
2PStlz/iNaw1hyBPqjAmIIpYZKqhoSEi9RvqlqSD0CkJe1wNPdi4ZOBfuqLS1zOJQoDNw5wQcNjj
Lu+7/hzUF5lUPHaFfJYs5lCpaF7H6rAntuoJylJqZs1T9d5HFp/cB+UniXBRGGYwJJPPFXp0V2iG
x0Qq1zHMbxs8xkp9hkwhv/oLYj7UuKDLh+lkNv1cUFadD8tv1AGSje2D/ET6QGBaAy3sXW6kTRxz
4pPl1+YeweVGkYSOGM5t+GWp9i8ks7n1zJLtXEzWIooArvDdHvgJCvH6ofEPt6S/qJGPYZTWN6XA
RoPQIPxMnyY3VUYAcilb8QaAuz0sZXhcadyUos6+EWslcs1H37h5f/W1/LdqQvTi77Cx7ELG3EML
TsGdDgfCh6jBZmERfyU37D9D4fVdgFaunDB8lSJABW9qpkexezOZMiFDgXY3sjcEtprXaY20/Px4
Z05cwZlhr5pyTDynjPx7Az7R8jIIleAF5Hc7lWysmzUiHR6r7RB2lFM/rOEou21SVuGLQg1EgRR7
q7YyPtuGThoiurRGTVW7zI4Hi1bvjAYCsBj70gs+hTafk3CNkft0Z0vq0RWLWy6Biim5mtUWXaMB
TXVofNR+YWyylb6NYwLGnY40KtywcPEFb5Dt+a7W11ez/Hj5zxroUs2+lEFB24Eui1/pm6Vdr6x0
xCNZDoKtdbW+9Rvfh3HfcZLKWqc+n/Qy7bY+VwTjw7E0AHnyZBEdGHP9XnkC9na9b0viFXddmeeK
0VWpsdljpM+ok4M1/2BFNomyCGwsFNiMPJ6LaHpCWu5bljwulhVfg/4u7rHVdPjy+YmK4fdcQJMe
bfWbUubrzoIZjlepgZ1bf/+obv4URvK//BWeDr+Syr7alCwDsfrcfIBnCvxLInTQtRfZI1/ofRAA
8Tj2t0m/ACKGeHBZ8bheI/d4WU7Oyt4fMIQzxByBo0OEuSaupW426E0WlVlXhLb9kSA8UzfuuvQ4
EbolC3tTqOuCwJ9MSi8zcOGxaQy36kULQYprxwUjNuO6kDVllQZuL9UFLwGqjDeGuX5tiAiySZWj
H8MRpPrVlo9r+TBBWNYIWWdo8VeobIGXjJIN/syrbEtRDmUTBdYCWoq8clfkhf2QeDDpie//5tw4
P9sDJamtkQLsMqgYWRg8qVYe+mbOWqL/waDCYYS19Qjyqh9OpkoUeaxIz/GZg1sV/gwsGy1sMr5i
jAwioFxarl1RPVngoVB/l8mdn0Ma1PCyybnJTBLYR1g1HzI+ZcNJpwBK1+MGHX5fJeUhDJHkQzSp
7hRNxTz3LT6IfCPjT2xhO0rey1MgFM0ESkOiGab1VfL0p8isUcDmK0W69lDzwHuyEi7ioKLLfkMG
ONQeFmVe1StekNNXA5jzQnHjXbNf27gePW/vhakHmXzdxkyme95DLUQwadVgz80HmjmZvZtlpdhW
PJl1XJ+mqVQ0A6culHyFgtzIF49FS6VljRQ1sExN2IekhcD3dj4s5/7u6wCQA0n/kfOEpJZpkK14
/h6AtsIbFMMwJv99zmI8EZVHlmbRdGL7BwdYVBfC4PrIfmECHSZrTtnxS/3MJZCHFkr1sKOMvZDU
U/sjz0e7nakgDUrYLJ1ff8mxcenrlVdv8JB43fukgwC402MsicjNEsKG66VEMYaryU0vPdccikox
dPTtSndes16g9f/vPSzgnb+GaMfWCLbXlSUXMoNagQIG2smHARxIFxL5SmMQJqW3G6T0Xt2Yv6OV
qNYlflcInL2SpxlKI/iYWmBLUf5Rqv7nmdcZu5iHusW/XVZU6owkpyItxeC00QX8Z7Cc5M4dqmuu
m3LL7yT7VLsY86k4BpnWEY1RiWR2IkGkyBMyAqipUcUJnqw8qQIb25q+Jj3aJstvOvBdG3tloNK7
Y8JhIhuK7S+hD/prV/dDPtYE4El1Uq+mDgst5Ce3C2MO87rBWJgzTQtOgZhOHzEdGCTupz8LvHNk
4SJ/kPcvlceHD3GqVrusdLjqz+mOYmshPWoTCzLaccFutJoD2xiIbMHI0wjJIJ45IwPAx3IPBmPw
TXlOEO4XUlNar4N0R3dd7HcMoVPopIH2PR8KtM4r0qKcPOvL0qcYdvMwVI18rW8iBgv4LLiPWiZ2
BBrSo9AcoNr3ljqXQW6KdMvHEF21ex+LziSaCNzBeZofeiCzEWfRU8YgSJq/Vxhs/lYEqTvd3EvL
SZ7KlGUpIEKLjPBP+uFopNAAoigV4k+oHu7As+a/FlhGdgIeLd6V/hp9eXgZbcwYzXFhLeXjidgQ
nwnKT/P2FTU3C7dHFJApofu6UqvbfPyZbI6ul9GJJrM1x2OnLeD1GM7+R9+tWOxQ+YhRNK1OhSv1
557VLNcEGVz752QkvtCkOgSg1u/5MiyCXvCPshflahebaCi/ucOI55cOHR5/hY7XeMZHR40HepIK
/k24m/QglRGeDMHVD8WuxXzS65FA3db7TCxtSikFCXBsqAvSj1doOJTapOWWcFZhfd3SY08dxm2z
6f9hOEQVT8qKYIaG24dVloBSPeSNRR2ATb8wIxvu8wbDL1LmyJsuTf98L7oBtBRZ2EvRn8e3mGZx
cuqbJjx/Gomb4oYFRoBgBcMGi4WWCcUnztC0WgFYb2sVk+A0zEjHR0pOjW8x3FQElFP5GFP12amm
2aH+ZS0teoNU3RRdip0/7Sq3JdXM3Mdfo4JxUycjmzO3L344yuGXrYT/fxrrePUNkQwcNtSkILcO
0m59hV0ifZi4hQqyveNCrMn3aaClYzhUeGM5RuaphJLemurwFpCY1dNMkcBbicsICfkX9VbIpO1H
Zn8to/36eETU58Y9bALdN3eJJxDJDT7/78slMeXOsZCNZbsSAZ5zbgZrNkJaTjZ6kIY62qQawn01
uey4cDly7wvoKPRbCYDT3vVs+K/bsRhAhytAi0r+qz+FjjJibGWSqIRoJVuJmwo1VJlu/5wWqukW
gX+5krHkBACYq+F9Fjd2b6EpCyxIaKDs5xWCOfhva1cJ1Z/iRqnPCePN60NI3mswIj++EqJupiT8
U5J8FZq/iHAHjL44VMImVPIkwvQDd7htg9DJPB7cpt3GGypWTmevuS0MOdB3PfhVkIZvFiMpXjQ3
KXUphPp79lSOLNKhaSOHuoL8JjCaqCAiEssPT4TRFmQANSrto1npeyocGlJvCg4dcC/fxPAuqaQR
w9v0QeSX9JFeZaPRHJ47oKmrKsvFL/Lu9f5knmEs8x8NkVM1ITb355FyeZZyL/gjs0CXUxeER6RB
jUX++6hzL6fObqoBtNJ05NFeDqoVqk6OfXPrCZ4tVRqD2+jUXpDw9p5cwZFwyMkwt2wLlBRSvRUn
EScJ25ko60vckuSKVzv2n2Jf6JKsjpKV4ckLASm5kW8Jvjvop2BTKMOLEzdk54Evh4qY3aXJ3Zqu
xkiS2GSz+FguQZ1CSIW6/pL95NsZ7MvgcgFxnZ9J3ltq9Iyy1dMA91AqCkhTA0vpBJVu9bl6/usk
eIMx2dozzsHLE/it1Z3VZuvPniZW67EBY3DRwvdmdbOGQfbz/FkIc7HmnsXi28N3CvEDhC09/NMF
JrWiCIICnKjtBCLdBlDK6ncs+JSKJErgNj1jKqor2w6JtZGMT8gAoFm3enMBc3b9J9MV4sb2vAxR
q7kv/UbhmeJrXjlkOU4XUcCbfh+MjDCWPNQm4abQYhROGaQQI2qG1oFfVbDhKO2UKjagFxQx91sT
bSWNrHmmMbml2alPCBCQ+Wb56HreS9lbPLLdORzOpxCG9nbEDKI3BsQsBVnX/JQBORvFbiRqS9IH
eSs+Wbml3+K5T3XtCBAnK+l+NBdNMDH/XFdesKedZyJlzesl5ZGz5UZZQaBPmoVCDn4I/AIzEjnA
+R1uBDF3X60wqPIfHqFBI+TnfxFID3kHG8I2GtrtMo8JQ5EHEBWnhz3Y5f7LGhGYJizAQ+eDBBmQ
YxuiWjfjROXpeu/HL4/7N+UEzW8jTedXwBbi5tg/wcGD7u5GLleo6lbD0W/c5TAgdTKuZTfEjbn6
zilC1zuMYFzE4cgzzV29TRrsKmdrpeGLM5z6tAPsLcmzViEjn3SCmI7FjL2JanYGc96i++lCz8JE
o3fXV0aZtUzLM3cG4Mw5CQBjpY/EaKpTg2LiVfQt+GaU46Y58BFiTa+q3fcoe2UWxueSQEZ8I6RP
El4TWguaoJIq82j3cIDYflZshAermVMkOvG/nllq8NN5g0vcfeSA34ySSDWomc++rKuu5fyPMllD
qC6e62rmZ0PAFyi341xwAv4mt5K0ZSk5OnDW3BJs1dvbdneXDxXLiEAjY8902sE95tZU//+vzBg3
0Dga8GqI2WyKMoCmMKA63vbt0Fjyi2XwbdmI6GGurAUK3IW1/viup1UVWefoOAjOZWhnrpB0rRd1
5D2Dng0WqgTHaTjn0N2YzGLbAKtS1Xff3b2xoDCk8YYulbvprZwoAK/nxdTxjScvNJSZVFn3wvJz
2U7W/nXJWhd6CNlGFa5AaVUG+jsRGJvMXyCyYHkEHtCkU5lpE0mNIvzZx6KYEQ7TD7xaQsk5oCEU
YaxuTfikUosvtdRIlSwWLCsTvTxz3mziakhF+iwfj6oeA71k71+KgCe7dM68GM/7kDYQ6nvdcYMU
/vwpOLUaZt5CzJPIL+uMZJ0a9a8vjulv4i8yqpnfN5tJp7ioldZ2TqJnZrqTFg1oWM/c9qnA2o6r
UllwfMA/BmCe8gHobRK1WPpj3MP+2/7RJ7kejoEFV7RZ98YNT9ly2QJ6pdCpkL72vvCf85CBSTQx
nIxwQO5xvDve2qDJYUj/lF0h8DHO6Csnz24xquPJ5V8AqsHn+U8Ig7ye8OJKSnmywIYtjwhDqfIs
GTUuVkQfqs8Pq/AzHrOv1AbxVKoqWlksIlNNFyS4EOHb5lpzcOQ75TipS9+ttB+kOo6P67kPqKoH
3mnAwBCSiuEIxVNib3TQlFY0dagP9dqUWUYABtFKLrsi+9ZOICcp4vlBaKUkpuEgjO871a1yq1Rg
b6AeTk88smrmVj4TcMX71fWiK7MP5gX1OpzljloIBnB2hqqH7qd0g+3SYe7GljSIuWiY502La2IB
g3d3hJnhKeUYVwO4CSnpIZhWreWlnzMsQrYJBVuwLktvS3xSCsszmBp2+qCKKW7DDyCSWoVeIYuk
J9eVSwvh8F2p27Z2XRirSXn2lz1yHDczGv8ywf4G0DZKWq9/+ZU30HvBLgYVX3fe6VfRClP0+mY7
jhoNnHsl8KB+azNVy2jpS7wSGomSSDTvMhVCfjnD5OH53x5EsJndnZKql5zK0TXuCDhT8E21Efz3
wRMBK67TQi5blHXH6U2f8VsvfxzhPe0kGEdsIR7wo53yLnh4ldqpSHO3bUEnjB5Hny2mnBAGwPPI
OQ5LNgHA1eTQIo/J6dK1WSD2o5/CeuhE1QimDA0EPxzBCakfYw2kPmfY1jEISTZx7EfJ18wEILGe
V8DavA4z6GYdo+fSzu/aFm+Tb1GXBeNhpOffoaUVFMME/RokfHFZwqYZXfZqunI0vISf8ePrMS1n
56tHQjsZSdR+ea/tGCBUaAJvRDFATz27Mjq4e4C6UYE49cnDEj/TbSQBH54FMRhlGmxVL48deps/
UMXzcmifPbGUeHoCojutQiPMAmplqn2Bju3p7lFKnGYLH6pet2WrvHyST0FdJ/4O2XxSkOAOgpeP
sT9O8hhNcDJ15a1EPt0n6p49jEbpZeMzQve+H6n/CdX4WvZKkH/JQTlHdh3U4YtjKSkTfH7itlZ2
1HtgiTD5xhYvZWW6KxCKz5BHbdIo3Z79ARv62Z3xH1OJxfv1j0q8+6+LR1Utv5Ac+BF08UaF8Zwd
KcoWuH3NlgTzwl7mBM84bfIm2JOVXm6/8ahC745eeq3SV81sujSfwGS/M6us4eiHM/5COkXJflFp
pi9te5BrokIirq50opUdQiTE+jrUZ3UpzDvGQKtToXETwhK9ei7wG+I7zbkS0z7ec7JsSfDA6ChQ
wZ/1Tq58B5W2Q8G4kKQpvRlWJUmcaTBTtBR3F8rF8oTWxjUxlzk6QSFa9nH4VIjFQTkTI3CxxiWU
NU1NUZfYGdmKZJgBcm9FfA+mVaoDr0RMKiYlMCpn2FwNTQlBktOAY8aEekSwOy6fVMryNumrWdAR
zviB7amq1kJlMEgTi/SeG042q1APNnJ+b28vhxL+cxty8jGL+csP37OHvzUq2pwI7VYeqvNoDDH2
9kSvTmCoNv65z2Dkn2iqiehDW/0YjWD0sINuSdnHhc9CJ0xwQWbHt6cOyo0zJ3h2nuyLnHwcsXeY
MSyYunZgBW3hcqhXMi5kNfcSHzkcThRqWJiDZX9Tsq9hbd/mCnw49Eq2oxeH9cpGczA7nyn01vdf
AFHfq7xkJQ88+f8XjVZfy6mCDSFSMgscDvgtyb5FwlhjPEwKpsY1sD25/wZgevsVusCk41VI+CJA
R7UQKuMfpCVD+SU6VoCnbxuLP18brJa0IKQRm0cJRaOL9+6BqbIyicIzQqut3Ko50QHb2+EJCQM4
jP3C1iW9MQTyAlxcUob3drg1EOsFJv1I4yL14wObKLPITHlw2lx6cTVo22mq3aEaVRZ3TGkZQgJJ
1bd5kwHIWG+60o2ZbNlSMJ1vRjU4vkrCJzestrfZi/OmcmLV2u3Q+UJChl2K1zqdaxsoo2FJA90E
LF10kHvf/ZPUsBxiAMRXPP54GcKKC9F7+LMOCpMy8TNA987UiIcsAHZPmjg/baBsbZ847H5nfQ5C
wT3yl7B500JW70CqCmaekwNFoyVuF+vrU0kB/LaBT/AF2I05pAUxlZYEDslPCMn/3F//GXWHUyKg
BQMQWWuO8Tdll328ZEG5+/szHEvGqWlIblr1ZrypIWxasVr4XYt7Q5JI3q/C9/cyIEsHQPYLPP7B
1zvEapmkLtZFfL5LtuFGw/RHUOBAMU7x15j76BLOvY7DlWlCc+MdSsdooiiAFHMbN+5w1acVJroF
Zkmugx/9gaGEwSw8lKAE8l0CEykwomyparFGJ2o0eTnXIALzyDp4aNzxgT+rYIqO4Ag9y9BOiY8o
SRxW7D/YAyU0dRA44S3TDW/umIAeD1NVxAacuEagcgMSV1RZBk222X4kGbVMu65Ex2awutFyad9o
QqFOM1kS81oWuck/4PgrM15LwG0pxugzoPPDrLtBuG4Dcw0YI22ImmiliEUByDc5kYop2d4iR9ZA
rOpc3egdcZeWWuUdbacv51vDD6ODMJwFIoy9YeHliFF0lKyZbrHOzbbuRzw/W6rkKSwwHqTQZVPe
j2iKYSZQxMCqtGHF2HZFQ5mKq8fBb03K2Tkbu42gDu7kO+1Huq/anoCqN2BF5SeXb32P3/JH66AO
F0n8vqp4gIspsxKAQBSxD8ipuB8B2YHbAGZ8LilQ3NOreqX+rDSdUAvd1/eGu9r1olCB5pqxiet1
Dyi/S7dhNpHqdlAgnGMRqwzjjD2hb7qhubKC1sxGhQzxG+PlPwhCw+MJzSEy459KzknI3noStEj3
Qwbpc7YYdCkgatO8L6ngcRli8i9B6YHYiELj1LYuQBpCKuJ/e7SCUJ7rsjKrUrhyHs3Th4WpKBvg
fqewpnJ+Zwuj4pLNzU2Pl5WwM0UaneyH7zlyHPRI49SjTLJA5CYgHHGuYHm2ZrElWMJJie+dlbWT
+usVnaGr92T8PtSEUU7BzopE9uHra+0+vMnfTlY88TkcrDNeaW8osfXK3HFDkk8USsYE+kMc1KKb
ns8eLMHWnaTGc+50VN1nddGQG/dBMaVVKOFb5otZzJF39S9fExwrNbIn/OI80x6zrDfWF0j6UB5x
6vzB1U6cRtMIUJVuUOwRGJR6IuZmw9nb/ncAz+Lze5GCLuZ1EtC66DBvQ6QulFnmwIA4hmRz0a5y
4kIvciZDsJWXut0kFosa2m1Da9z1TqKamcAKkJtIKV0MUw1KInmI29vf4PEmAlPA9X6I7duDZdr7
eFsxqD1AmqzuHJY1VATEN/3Jxrb5EO2zHyma2l6DAh7SwanMaxBY51xlmIYzrfxmXwVhWuqVIZrV
tisZE5wtlz5AyonOzKTTW47e7V1a0JagMwZFlD8tAaEPEEJWt+00R5oeq0nIVwUIaPaotn4j53jX
sjpfv01L5UCZf+zwvgMdbTI6dDB0+4rDXsrehhN+zB7gJhEhOni4QhTs5E+lGyMIgLVwmqliqGhY
g/PIMYq9KwkgLWk5WAxLdyayuNjTgAxD3ywRhNlvDXZLgPNSuBaFWbQ/JFhTpfe8nUjd7xRH8nph
6RQzJ2eX21Vo0qrVSQt9qdhZTkkLrg7TBhITfcQhFcs/nsxalbj9zU1RlyHVgdehrm8EiKB8fFh2
E55h9X/ERNaA8dma+B8C0X6oMG1RnxNhq8/u59S1/uHu1UcQ2dj/5VHMajqnyyqEORs7BGEmXBCR
MT1G7su2JAYnKmlNPqHFbfYHtS+GMZEmgK/iiGR0ek0wrAVTt57B5Agg3OisNYwEyZpIEhQBFiOa
i0e/qiTnDBHSpFQgE77V8Ntv4SLoKJtcFBkVs58rdCoCE8vbE/YK5yzgMgsoDmE4Ey68gmstqlQG
qLBL1Z/soyilMdOg9Ppwj5km51+mAsXfbi1BYtmzay/uPgVItunj801ilgWT8Kxf7UDwutPdcdYX
vJAtmKK2bHUpw6Haz7QZqo/OqJ4Z+/clsi7HjL55vau2ag5+0Ym4yd7uezBgWnJYrbEV6Ltn9DJH
Rw0dgkobFoLzsGSYRS/TMFc9zYll/oNiKQv8cUEIj9JoatAzMy10qpoFYkfrsjOiuVw7xmn01e+P
JO2JGRTgsWtuuWruTVpeHH7FhrifGVwZeSso/LDS5Xfw2AHUvxr/4ceK4t77ZeM7ZPx/wAFJmEuG
vR7cnWbOH689RFT9RlXQYlOpJYjtYS7g+5p5nM1JN6+1FFc+QX+8tRh6fTX1eg0MxczJiA/H/3bg
XTtzOIV/4wx0uqeDpQxs7nNVTv5adJRXjfXCKnVJRe7eZIP95pNNlBfj5WqiFK/dsEbW3o/M5Pab
CVbo3rGTwwfb63sEN1r/pfsPHZmTbm69m/CF/ILqQrecwjiDzBlrh/dsghLh4UGgUFSnc+y1u8L/
kQJZXEpZTC1yjHWvF7L4NLeQNsMKZXH+Ginl1eOcvbgCtFGQz8vCNqf6dEVkxYv+t0SfV5NcRLdf
8AgSYoNS4UV9Iyh1erD0sZPsF1xT2tmElTzp8HiTkMrXvcnZlszAWUVCy6ccxytrbLt9Vi/pO7LE
XFzFSrsFfD77txsOC2Ta/CTyAVIOr7aMSUKKyoOsEsvR7VMt+39CJUgQpxnsaAVAmNY1CNylqrC/
xKJHRQGXBK73VJ2E9sun9CLwSxXWNSWSH//pSjkFtp90Ajplg8GGgJjW6lZxtcnZSGStNjBV0mbs
+bkUnTnN8qzciIVLv3hjhujfDUnkOnt25vRCbQGvqZq+iQs4Q5UDxhSTGZnSUmCvgGnq2Fi0O6eU
ICaXWYUDIcv8E3/DVMqy3U2ywXVlgZXO5Ye2Dpmb2Q+sQO8F9ZaEKsncfl/UhqKfWsY4Fwn6adHv
yu2ULzOruJ+bWtyym0EwuuyOfPfJ4G4wzKqWhzLcBjhYfcmdqb279r6c9crQtt5rGKICZ8+ahE08
2SgoKJYztTYXLwSPPs3UWaLxC818xTc75Qu8Nz10YHlvDU5wtcbdpKv+RDuNnyVnue1mCD1qObIr
s26dIea/IoExh8R01H403IvLBvasjyfS6QbFaXMZaZZokO+JpLmPz/COO4jE857SfZVF1TXe2JLn
xxukws7I6ORK5DbJWeNxe+M+XVPed6kmIOr0TkR6JShKwJh25fd+zHRNnp4fc/Ekt1k3TDymxxxL
dpiLY+RD15AH7wzlsL1v+NVvLSb3N9M4QpN4ApcyhhxEP9UFrhUzXJGzS0ytnFPEB90wdRoNJkMM
RC1u+2YSSabL7MNH1fwqTng3TLwJ5W3SeUm9KbXj7nSP+eGgUQDA1swa2Oj+CMr0Ru56U9NzEJUw
bVo+8AThIf+9bMwOOgaKDsIGKUG4lds4oeb7SVE13tb9mhhayPJtl/2oE58RSOOqqASwRdG88VuP
HT1nAmKPAdCLq+LHICDAk6UwZgp0+NkDYvCVz7l506tcm/2LoOU5H9sMCuwYhOMvqRV8M8E4+heY
HhEsWwzfOocuDNyJ/ZxTPDmSEj5sUXe4KDp94CFbXPT7Ve1hUMW2vwi+CVMAZj9wHnWau2zmceBS
pq1YVceRwQZYgKCH2PpoCYW66caTxUIC1O38UN7MKifOg6/Lrp6ftw4PpbrHflh20wAT+NkewRse
iaLWyIZ7k57mAjKysfm8W231PRyINoUt+AFYyiAehscEUOSi+WFixhXMiTStFCh3/7RcvabYaqot
Cceg3ffG8z0spgaFW0+RoEo7ows0PyV393jFm8slWrQZNBCkswuE7vTMTZg9Vdf+ZxmcSuDqpGbP
mJMndAsWnTYzAtJYlGVpOe52wbhRokJgVYgLSoITdtdKN3T/G7uYgikXVl3qo8Fn7N3uIMVSzn6b
Js6ACJ0gJq0Ww/dVbZH/89i2B17HA85Iwbc/GcBDKICr5vHBj5IyN4SngJtDbN1vfm7AxURGEWJC
uPH99WwN/7SXe4JTKdCUgNx/ZTRMOJK5pvOl+j/7O2VPJJEefCCCJpfShgJsaBZvIL98Bt/JFbbx
p8A65k8bwWaRnZUrnF11HuedwPIUrA9jEm+UsTtj01KPczQyS25W8PoCWcqEhBIXrCQQ3hSKQPH1
r1XnWCKNqoKwLVso3Bv4VwsZJaUj+QmKuO4MxPg+93CpATo18hWd19+wiImrqDrQsK00bQmEEgLL
zWbsAEUtHTu1aOSaz6VB09JUxSNfIUAbxhg9l0L1pPuIzGf1ZypRWva7dGbgCN7BfS/adU2Z35Z+
C/XPVyJ2k+Zor1CRgYRwm8oFhUq+Ix8Zs3/ojJjtyFJKztoXstUkQN165kP+ZyhvPuaJRWzL+t7Q
pqPys8AwrueKYpbqTKtriOFqEUz2xW0gIWhYa9jiUf8rMQkf8dQcomM91mXyKliDC5hk/hRoZ7A8
+DueX1H1MzbaKOpe6mpcazj0Frq+VlriReobutzJEXp8thGz6YLCdx0HwEXis+Uq0nzmz66SBOM/
3knMfTjxSLGAVIWNzzV3FNJxKBbMzfqY+X2wZL/uru8fgkyZjcJv9Lr63Sq32CqCpRPjRJTZVxJa
Kd/kgU8NjX1FQwibTow0HCgYaGMVoTxpODSaNk8rhigBV+spGfUUXSLHGXk1Pxsjln/zSg3aB70+
fqBfdh7f8Yk0Sg40r7AzhoeDc5isfX/ja3akoN6jOdrSrFp1UtSvYJJI+O6/VF2sNZcK3PQL2v5s
hQUjZP0VDRvPX0lBXlCtxij1nOD2wf6lil8fc2mDnKf7Vy4nmglcPsCyNkA6D4WQVS5z44klHsyt
CpMQDYaEgupdwDKfQTxIev0K2yApXb7fgpTf85IR4JA6Y4hxFZfSQF44V4joVdhTaWnNm22kRBye
0MvynavdWL7vkI0D8H6HEAPMNS4WAWn/IzIPMITqNHunUOM4xmfVnA7ud924hyjxfq9hieNfw7i7
K6pn6mpH0jmxEjm+MlnA3tD4EN2bPev88gviMaBgku0CSlPMYJ5T33AgYsbHt/YkxwmLrwiBOw0j
24SGICoLrRhwK7mFm3fprmYtQ7TqC49TZl7Nyz9fkF4HYwR0R7UqWL30JmI3tpq3fc1Coi6S4QD9
BZVPTkp0pnsol0FOsopggvAgvWn7mWOTtcSDIuwFJY6QwZJFtCiyAr6CASjL/d7qPd0xhfO3q9dl
GXvDIVvN0WvvapU+y6o7o7EVZ7+//fUf8fAyJK1BeuHJ+nB9BA9WQ1F2yPc1qIVkk8vAlSqNpokP
MCCg2uvkDO+LVlUETuA8NI93lA08UXZm32UDWFGJ7LRFDL42R24g0ctuueacIfXVd55EgzushIne
LyUv84GZ5XE+ULK2fmtC/cwxzljzwuoYf7XtXk4X3II154tRQPiwfzZtBob3fsoiORzrcyXFWAXQ
P2licx6lk1BkBFjJ5oFauFuyLIFN6X8YI4Nhl0n3vxCvu3E40I/oxeb4IPO5QzdZ4+JGbeXPwJQr
rOgh9v4wCS2KRLKdcBTxCNE1hEeo9S2A0mtc4s1bWI6szT4FyMHwj4nYA7UA/yqeXUshOjoiBgA8
dmvkCbmx3hRVr+4YxyV4L8abjk/svuuMwk95qZjSGFdvnLxcKWnPhBiTZzKFa75aNv2Qivt2/q77
ikzCjovhyo7rqBSE3M15KJ07+Y0Ao0friyvMxwbEGA1hcTpIfHF1a3gJHKDyBGI7+crmDNLVDDZQ
4xD38ksnbGJIZHRBeHDY5SLQnK1BlZV7oRPeCJpDeZu5t14QifsNUg3UdeCGJBcYElMEiyctUIxU
i03He9CW54JtPvsMDqsWhkspRxp1LJz/0NgVNnfUnZGhBG2hEdmqOagDIZ3R2k6zJUiW79TUnE7t
RkxLszH8JP3rkVwfAJW7KtyW+tBCZBI90/3aXmTWLQF2zE+q50wWHu2xIluS05hwYy/xlsaidK6s
5rPu/mxCDq8i12uDWyQxY7ME0ZqLXkDqXnJUBfPiHSMRvBikdytJotcnoChQ4ChmUMHGUNobqxYJ
VIyqahOijZP8NBCfBqfteZMZFGV0/AHfQyBkFU2enVZMn58aG2UdKsmPZr4D8IoJm4OgQYa8JVQI
8kOLqsraxMDU9e5/YPMe6Qw7l2O5swhy51zjflT8WJ7lod1Q4qU09dgVuKKmmtAYhKsb8GdDQFDl
f04v27LyLTsL8yxvuHDAJt6gn0K6J3d1kcjLsmGgm6u9hwa+LXh9rZPivxpPY+MAohPSulicD1C9
1R0kx0b+J5BsqisUHLdpjt3yvZQ2mmRiT/Zyatm/+QVw0YdSr8QCBDedhlIJIuiDt1e3zpe9TY0r
O+ODZJi3EBeSERje7gk+YL7pZefhLhmqaP0/rZ07Br+HNCeE54YOyzmjREmkz+pgjnx2Jq7Hw6QC
7NnHYjLdVqs0EwHuK4HCYr83L/13J8G/jx/dbNfhKCg4TPk0ZPRm5vqY9hXjCbndLvflyQLl68RU
LBuD59hOtMxG3I0ph+57ug1rcTzDuyzZl0Bf0npTpoGsFjsUc2CWsxCExj4B2hSA8+K9QXrzbnBk
z1JnHdGTIjHYilfGQIJyi179u39ECfGu57DYKFkgqIec9hL/eHlWHVzk4ErlIi7lj+xns+9llm64
EJXQcevLu/lI4HA2iX1RrA2LSjIStEfMM5+ZL+B7DUBu9fpeTaiueLZJgf4pho4O5wS6I99XQEw2
t+1sYSA0e7n6FTdsaa6FKfSM/GHKY996etptccADH1PigZov23Lp9vn0r2WDBSuhbmzazYefUGgW
ab0bOV2mGwfNZnydxrHpgfoJzyTslTkK/C7Dpu5i4OC7Ti6jmi95+mOommpDEsIPGt/OFEWuUPmj
BTa47SOnrT9HZYiooL0hFqFgFFww8jfxxHIxJ0QTLNZoe2l/rngQ+1YyVShZvQyss5hB8VQaF9RT
BK+JuE2HsnJxv3YuHONWSoVDkoXRfBdpOF0QOzD54TjfNFGhsJk7epZ2mWFN5dqNmNRtflfN/Nu7
PiQXkWz1bMK0+7CMuXTP48NihWnuQw3vFTTkb/1Hc20mUCRbQzomzf85ZteyQdAf/jvaz9Wga3/v
yURSRsb3xnDcZh6ViCRLe0psvxC2LOiGop8rWVvXTr04kS0GmqmUEqVeJQkMRPKFfzjgjzImq9NP
JrGE2CrTxhPTd6s+BDUwTg9MwW3biKQpVMAWuj4bWONd2Wax1yuEKDt4nIYjWW3HJWRqMNWZMYB+
PH74DhzDLnhoux510kmUsiIc5DWPRXTiiUEEROEdIyDRAuTi2EFzvHWBr4u+dTTdEj6OyAss0Y1L
VZGkK5fO/Cm+PWlqGKwkDq9Dmo9HWVgvdaBuC6CzJ1cAM4fzoC41C0DAWBzHP53Ckm6KrucT9WDU
gl3S/5rRQyGIkLptZC+LRrsBdPdXfa4Ze2SR0M+76EkOkQut5sQRX7bIUCkHwDbRo+iYIeUcBjsD
qAddKDmnXNTRRMNEFsQS/uDWwQCJPDoG5aJOiLJHCXVk4TmtbQ748PIH1sH0iqkWi/TtLLl07EEm
ProR+hsBkidHunbKooTJm+gLwYPqZ2jTTgvt/Yqsd23kb+hrlT09RTo5sTO3ErC6TqluVH7MRI+8
xwSLFfHaiKV6RmbSSySodg/yByW2uVrYq47ytbZ3lDxmDvaR2OFun55rdlO6wOz0ISRBAwJ4MzK7
niVGsul00anFh1Q3VipT4lxZlHQYWp5z6irOR909evSnreHvEv/x1l/cEEBqvjNPJu08qLegALpV
+kxRMek51RxrWvrwZBLT/vQFbhBXbvzCpR4wu9S18Rm3skNo9uiwvP85ZKPWQ3tQSzaEQ5zns4hh
HpbLOhwlGJHr0gpY8YP6OBZ7bz3OcURPNjZ/5l/bgj7L04/UwKllzeQUr6LVWwccjOUEp4qxahyd
GLOvS8/8JGUdJGhi1iCJHGgYlHDGlPfsfp7SL1R8k1QnNrRlpLj09qoO3O9RUWDXwb80rsY3nVVH
ASxBLYyKQYzZZR7dAwfDWfJlHPFCTj0WEG1Cx62WRFyY4cUL08lARxIl0UNeEVDqMeIxgou4Mja+
yfr5BKN09S/vJUHUUzrVriSMVxyuvosbGB0GoXuDDX+DpJIF7Qg00DZ1H/R5oYEYmkRuXmvOj+lS
LpVT+AIiCIAuRrndugPWaXLJZXyoDgzyzHr3ns4/yYGB5zyqACyBaiOHVLnsdlDBsOIDCQGOQYPZ
FmP/VdMA7wK3UhwliGvwzGPLBBcB8rCuqKaKMYEE7uRmJILaRYENbu4DiBOdBjTIEKwDib1Pw1B1
sVpfN6LsJFjAZwGvyhLlB27L1LGfp90lktAdtIJPJyU/L+JYj5UK7wQXNLw8jchMQ5RbYs1a6itr
/rjNEHZzkwpkLudfq3QIeJl9JKWvUDypuanBAxSawBjkxDE/NlmaMt1hi9jtfH2OxjBGC3Kn6iON
yz8/fttKsAeu/ie4rm9XJSyV+h+PdauIMEUXquSdKIgqCzLUM4DWA7xJOWLJf9UFbIBZ0170ZV7w
P3cXGhwK5wBNqc0yA3A+oaTIy+7lUA6RMlxJ6jL0TCXY8cSUmVs4E1nF5CVoEe8OFkj1C5Af70gy
ARMXeWQXj1nX3hiHR0/RZhe8wl4udf5UxV8Ozp8GXkmVqKAfkstbKWV6GC7WCgGb3ErTtp1CfHJf
ew4qKNmeGV3VbOOqiGjeZWprCAE99/V39MWlN2uRQIyDLcMJBHcQPYo/aniz/B0ODxlfkw3E+GHR
pzCGy464azcW4pUnXG5YVvQTOtLMVkSH4+0p3YcsvOnhgfRDPXD8PoWuISoAwhE5ht01ylVvOpTO
IoZWAwKbLlZpB94ZJnZmLPzCPi+KULQ7qOE/C6yvmRYv6jFme+NXv6np9rhAT5MPYI7MG0tLAjUZ
FW9vU52gFUfBpULl3fSAG/xIV5ocMWWGL5C+8sCW8MBNtJSECr7zbhvsYKbt6ReY5srlz2230Ddz
r/ygWjlUquilzav2+whSPCTBjhJ9VDY7SJ7owcIcFfz9P7US4FZwwiAfrcwJyJ6UWVnlCpgU4me3
6ZTAWyeBl6c8aDF8VJWV0wGMh5W+31wvju2DZoz7xKVoIT0pZTfHKBORdHe0AHSoEp6ySkB+AG1W
NPmOorq30utu+Id2gr05B8hwRwYRlYL0vT01Km1ceOjIZmk6+11/KQr+2UFGS/KoKjh7eJUhNRCJ
pCkfEhyjdXfevZBxxRmIIOljxiMLu/VvDvaur0qzaILTG92xVxjMRoDSmAKoc4yytckdvqKyri0L
g0X+bMDjhO/ITUk5Uvorfr2nAZkwCLrx8HPBVKEOsPc3GNIfnxP22fvDRagw5PR2BX+BxLw9jPNy
h8izq/CIQqDIZQQveH6HrPC89joD0OKE8EgXEwzlYll2rOkwDRMt3GrnLr72hgIFiFDVz5j1QpQp
ssSFgtTrBVc171g1SWIrqCbq82jkcShI9OBm+7P8AOEIqNExXz85lRBkdd9/dzrL8Mnof7v7CGFP
sC2eZSGaadgTuv4KbhEug/KaTiGNck63YC4F3aAtk96ZOSRArKcDH1sc1yICu+xutWFPYAR/oAAm
bp57+mLWF3EMYQlYs/ApxMvecZEAgZr87yrt6dT3cpDS/Kum1Qf5ekv3VVRi684TjuOlXwbuqls2
7fXx23N0LfMaar/XryySNCkEGuQdluYe28W3GdLnC/xUSBWSaKqhE7fk9oOXABEH7J8YK7rrnt5c
GIOSF2w9MNrhcjxet4nsydF/BQwhwj8vfiv/QAPfNDGQNE8XfTzAbgBkfSEwTrCtSuRlgsnLPLn5
7Au7MfvA9TKlHbYUC5Bw6sS1t39xp4Q1gwJXy9aCY1aUpXle5j5GVCHk2N2QOX0hrffnqkdoQpym
oXx7mjXjsKcsi6IBYaaaCf/s2gO+Ym+ugBnulk27YCHflyQ4DeqbvEuluC2BCGBJlZcKNTrFsKDt
9BEn2SBO1JOL32ExTmrrUYvJlEgiAuj5Hdy3sssrfShSSyZ3OxALAecxtRA35clFvvpj525PuUxe
QqgmwnOGyACnhHT+OIBx3kXLoZ/Gn89sksHR+kWTZZMVWGEabjyDkWSIGttQeW6C92LuH19irLWM
GbknSLPQN44Y1+OjEVJiV3oPiRWYalD4vjeSAj4UZiFnjZ92mK86aZ/nr8/ZCjJdBOMdwdODrsZi
zKnNvV8U+kYv6I1mX/XtGgiR5BEh4VVTkQxUCggMDSHZkZqRKprnvnRv5PKlXOnhdWOVuKLqJdVV
kKuyriJhtj++Rm6klmHM7ZLR8Yz79SzAci/NVg4LCBL490EjkvBPDt5pGMwRBuVOdIUtuTSSF2bW
Hq9UTtHBcdKU/s174vKOHlAmYCqvJmMLtEZmDic1WED1cdunxd2GB7I4oO17r11fc9QxE9rvoS/E
kwtb6GXcpVJBqFV4ZUnKw0ev6rsUkcKhgOFfi6qzJSNy4AQc/V7V0JwXYCmJO3tHh6zyOyn9G7dx
etu8jRN46fHZtsZEM+IRiCyBqsjkBByjQHAgar2lT2VFkMRCz5LyaewbCkJeL5nTKuMJe6eLImUr
KA/KW5pU4Rcqf288uNxOVvwNxX3SgzlsmJcb4gEqJLMsyCBydUpjxvbIu9azama+U/5UkYE+jvn3
kbqBkm+ZQ/GIqxXIUNpH30GHjlKERaq25qb54oI7GlGNdF0pTwXt46PKNrPcwnrOityl/pFzzYIV
ZbQ5CTui+ubbUkNuGr6fsQQaq0cc2D64vA0OzWLzeX+uYIBmmk8mrfBJo0Vn6lz0IfaOklWaVij7
BTwhbHBYui9xNGYrOcl0aNvvI5wbNg3k6PGDjMYrO50ERjMWMOob21ibgFFnVuHh/iDI7JoHOqKJ
yxXqaHUF1H0KbwOT8fnkP/UnwoozVzQXcAPC4LfY2GePXE9C8p4RSVIZSIV7pUSHd0oosBLxUj1i
+h4jrBMY68Vca68WDTr5vP9vTmi+tnr1F9A5tUbbd+DBlp6/cfO4eEy9zOmkBz2pFuVQXjqmHypF
tyu/jpU/dx/EkdNdooHbXtEJaw+ac7Wbd1VWte5Fr4HlVvzt2SfrXOxAHpngwGaGOFN3TB4Zu04r
lZB9Cfy6cysBziMbJZnwHe6h5C6iWx8VJN4r6IyrJOT8IHW3nWNPyUjIuYcokvg5SBRe6d9oFGAy
shVt+GIwz/jzvYYhPSpH4ECz1t2ltkSiweuTaNudrde6VttzNWNwVfetMPTVmDScp9F6MerPqkQb
zeuBJ6mjq4YeoNKTwpljJD0J6vFnkEL7gr4Qqvt4eLyyN0tJsuU8UwGalQAcKYeZhbtLOXtD60DT
tMLoTgIPh1pjhuehL2A/ybdqyntkz/vC9rfpr0FNvHMkcmEctWcnPz5W1BtPmGJWlE3sPtveOFoI
cNv+gpOTwXCax5T4DVmJkIt9cMyRaNuiA76aqLuUXPvpZ/LbnA7QIw184ROqi1D9iV+U6GI6NslJ
Me3kKePHaro1peyWhPjX1y0XcyJ/TajyfFQ1dXhWa0K9sj5jOLf8tHGJRA8AJtRnzV0JVZ1QnlKO
b8Psf4S5f9GbXwn469I1lSKtHoIumz94vm6rCUAfjS51YhGQ0+WOH/jsllWxCYkiL6QxRWMojCuG
oaQk1s1hxKbkFwHU8U2H6lXSBil5fUHO8Pu0AknVPOzwpVeAUtkWKs+2+uRrFpWFXM6vm4LXkXVU
NX1+9kwtC/FHrQImt9vWpCmS1osCliE3QzBxHelS/1PLNKfqtBYrLVHnv3wBdcr4cwqW/Evu029a
fdhK/Us7MRQh5MOczfPDQpXQJHrO5Di3aDz3DreYVlu70a1rNTGWZm8avF2L8n5KeDLUvTVH63a8
OAxLgBr1kJS+8q02z/lYJr5MQY42nTaA9TXLHm1T+oOyELmLnr6jSN819sLqcOHuuPZ5JGVUQr1V
CrP+/Doc9W0KIUP2IDGD61g1JlmcH6iAdmUUG+in+b1NqnyTDq1yXrUDEV/xHK9KNqL3o8VCmxVE
CkaOh6VwZwGyCKYhu8KTJzgy+LRHd20IqFfN16byr4tBPtLgnXV7Ku9hD9SlK2R7StdJaX5OKl3F
1OMwFzA+3mTAe8nrlu3HwUxPS+YYeK75DDk0+VE3juNxJw+FNkCoX4B8mxmBrLDE8Ol8458HQHvX
dgs31biJyWfoLN28UgmSp0g8Bp4HY/U6DMgQSLMQzpCWrxixmN9RtJpwqxMRIm++jyrY/6c/W/UQ
djSuUoI1n12d/FrmLWiwwZ84vwL1wZjqV4wx3QX8mpYqYdl56jNaQDDDHO1WhrL+ShbGRqBgS85d
kYyQx6x7HdcC4UwkG5sACXlYKoi67OpOdTe54tXEzehP+SP/F1LRkglLvHX8DZayJ+qDwEtz3+v/
FyA2LGfSvyfEBvA7RLjGe/FNlJd3hxUUt0fvvWUUtQmGuNxiY2RVMDyxAbdH+GwcRIQKE0olt8LF
/HFSkIJtwqppY68Iys93KOlaCRfr+9PCjBzslSUR2K57pwTv9+NdCVz9wP3Pj1AOPLWyMwEwmkMB
k3A5+7mvileXznJgkDyVgokjQedjDceIOD4HH9MwWt9SZvnZstjy+fSsqiHFN1cA3zukuOOrXON9
Nie1walj/z5D8dHPre80uZgaxYEcKS3To/yUcT3VRva5S9DnCOaLid/wrgBBAx+aSPHIjJrTNqZq
yCe3CdmePvarjMGJN4qLti6CnWcTNg2TbAWlR/V619uGzoDBKlERdinUorvFqnA4ksvxWUESqyeX
LXfSZfmA9UcjBPYF48N5ldE7wSargaRM7LdVcplk3ueIpa5EtLlIjur94zqVbH6MR1bA0IJi6vKF
I2zEy4ncIZ+4HwGxg5uFK6rCFZp/Mu8mV6gNX+P1DUTM8zOf0HqiJlqEB17gxd99MY/Y9MILy5JC
7pvhQW43XG8bGfUl6w2ham1b9uP+cFXNXbQmUrPG4nfN5P6guPyJvxojmG43kez/cio7fnkd4oBk
qlDgZHULmyW9dhwdlvB2kMUjiP4+kxFyqvOL9xXiVh7WUhewkJsyDX3dic717FSPzZ/5x3tXa+fv
Cw3PG6Gc826HJt50agFCZ3R/a9TL8pavJS70jc2cl1kJO3yes6FxG229E85OhHiIkczoFZu9g0cv
GtmseHdYFfPJ8pV26np6VgNfPyYgE7O3iXEGXF92llFN934QozibRbXNDc5Desn5soOOMoQfas8E
3i1TnVXNYh3a7dtB//jmr2mbCcP64oTySLL9E6+iHz3cSmEoo66j2o0bMu3NbwcwFBZNLDrAGLA2
yhXvV7n+xbduuprPrRcqwvdjE0J5TpynwGWwJy6N0KBMTNvCi1ImQc/VPluMb86XDRx5E4kehPRt
C5M60LzzrD5HsVR+i1nw2V+DC4fh0ixStJoMuTZnkWFNATdrN/CHz4tIs0yd/JLX7oOujAk0bKgr
UDPtssGL3XqSN7Z3XGB9W1Pi8iqgUftdzUEKVq2b0017qhs4DR+K9qVK5/NATnLaPi1P8XUJP7tf
ChNiprsSlD05qWux2IB0wWWxzUp7VNu4LiVGOD3ALu5yeaTfnQ4nZZ1RaB7l9z2dSbhjhIQxImhY
YqDHXwWNmIpK3HSokN7AN0z3wQ2uUkI+0x3o1tR5Cz2gOGHnIwRddYQv3vpe0kRNkN5M2O1yEiAb
aW+2fzvyOkah8cBbDY/LtN6KqUeDAomuLRvqfItqJGqImF9HydoN1z9eHzhdazUiBf1WMd52EA4o
ZcmFtkZ9WdTuiCgoBnGprTf9dDoJa939qwqJZzvbIoYXErpuJU3MLOnZFHISt5TE8U6YodFWQk1N
EoozUMGvgsuxSaHQLn5xxbK1OvB5EuMx9NBlgIgvygSNik/DMhEIVn7bR7ojGzyQ38thmohV73pt
iB2U2GSqmUzK2tJMr+Ml5uT3DG00wnUnfru5m4o7n3BQj3gJFLIEC0wqoMIE7AO6wQDjU0XY34oJ
fr6ROgCvvMRzajMJkQy2NMNNDVPLu/a0CHtqvX8hoK277xtUnpgk3yqWmb5ESquK/4WY/O/oyQ4p
tZHsJ7c8CbeOtGWX8+ZuTGDfJ58m8p8yK+MawB8Nz5qhuQycn1Py0Qbopcb1wSrPcRvq2fXxLepj
o4qkvWJobes2RmWChfIzMXPeifuVcqH2KLZ0hg/3knHJgyriXRLwRiFRQZQz6HaeZGPMw39vPpbL
5HJ6vnaL9/f5gUh6DPlzFQBKsPoj3CtKc2f7m+QQuQ63dblWDgyEVZhfSeIyLqS4uIQI29mV5OxI
Xf+5vPGwEYQrKYi/HCGlxv1gPYDKhYedudFbfuqurudCWb3scV7Kjo+bw4DILrmQXo/ENk9v4DGg
MgMiPPESkymvYGQ2EHfoY6rkIB3p4mV6TPlxyQuPitTr4/u4TTxWySqeOofGo66AFRIxYhhPXaDs
NNwAuZbwnlUZfSmOw30t1LtSoCtqzaj9iznGUuZezJWbZ8fGjNF5KGEXJALV2lVCPBlDnUqYi0wc
Aj5TQJ+0tLTnw98qYMFmkImMNAJUBxvexf6pxef1gCuXcKprn6N2lVIrQW/785b5xUpR7ZxPwlsb
Xbyrtf/4BDlh/7TVwwlcsb1IF8hkN6dmU7+WhH6alThnO0/nsYIiHWTnFGnUoS3oW1JAShganSWM
z2orVtZj0lvKPZ+/6fGUl85QKPIGXo59pFrfLhguXyXnWPAIdwSRV/fXDjJTJRRBSVW5MgU95TWX
r2yiE3L8fE+SHPtNW2llr4ZDjqDoE/vCMljGfj+mvvzDjK24pN1NFHJRUU5x6OL3PtFymkDQ53T8
KwpcEHAIqK8Eo1qP4j3GgyDFIQsc5iF/Zb3cl37Xf2GR1V+admP/fDabkpj/aGU0IsTxwQvAsYSL
begY1ih0heqLh1aVkdY5E6d2Ki6NkRbj7g10jpH7ssCXjWr66191/kF2vmPNR+rOQTitaJGbxMZa
bbjJeHwZ2hqgVxMWdszb/SLPTsphS7bPxmEdFCRypcqgViVD9rWyzkpYRmczH4ijwcTrETuQe5pu
wzV7GZ53lSV0yOg4Xu4HszPDmH5Cl3PLihxoWXSoeLul5gbir1TNkJE1ym7mVPfulY/zjRG583M1
GYUALSHXqJAL7uj5Q/ywwH9ansptMUsMjM/jICOn8IhQ8Wr775J7XNx5HJ8BumRmEGR+MiwBj9Mt
3eaYgjvoMiTEf8fY3gnbD0jEn4j6Xe6h/ERsND8ek/ZeisRAmydsBFJIM0mGQzsTHHuhadNQU7Rp
pVXw4cC99SySJCTwaxhBUAlRj0iBVuA8+5/MpO5NdLNMWURo3agg/VhFBmojFOs22EItTzx59dYF
OTSdQ8sU4MjGWU7eV2PV9M9WLk+qhQCXvVAsA2B1JF+O8kKgui4FbLPQECDvPwKjVdl1/hwURnFf
OK7rGcXqKSI+70+e3asXzoDtqOzljiu2nIEQXV6Y35AOj7t+VY64mdC6H8wsoMyC8SZgedJALZti
ZXwq0iWP83Rz47cwPXJO8hLLg6sYvL1bBH2rSuAKU6gerpoymWWfhW4G05/vsH/HHidu+l5BNZx5
FnwIx+Zma+gF4upyT8MHldWoVZzHfxd3lNUXYVnPTvbCaRFRfMmoLNcifUpJW1bLzgdiQlILzVPN
InsMjKxVGbIAi1T4UQkW1HK4YjJu1OsGg/088qKr3yk9WCDe0xmbFeCSjsu2l1d67gvZ70cEgw4t
4PbbWlqz08Tt01yC+pXjBogtGaL7swc+yfpPnO5PWTcFf5ekEVbWb7/S4guLrQLEtZWyGKVUNupH
Yqq9RMd3nn9tIQvPBqJsK2aONLFqIw8iQTv2E4aX85VYTK7xZjOPISwy+XjgsWR5ETpWTzQp2HAj
FFDTp35Rr0QAjgD2h4PE9EDGuH9roTzmuz6EQdjzNFUluO2BG3GmAN4dPKenjE47dVlD74AflVl8
NmGp52gQNRhjp3tLqua2vlQ70K10fnco4ValQmvMR/tI/L2FAjpuRK4goYpMdnAphGCG0C7znJY5
eXysSFM0m8QPqJYGEF1gMSCo6jGTXhV9yokan5nqn6fMpehGtVGOWhC9lbbMyJpWn1s/Dv+JT37Z
eeCac9S13npolhWJUMtJgdhNfujgeoQ3jVa2P0WK0Jbr7TMcNnqi4qRT01q2Z0QgpYbIRxBirRS4
8tIlzpmynwEhwcb4Qs2VGCnVL3AWtBDjBBUmorVTkPsDq6ZHt36EwqNF68CxBkkv9dsZYHB6+l1S
vv77s6bfThGo2WJAuXqW4CESKV0oUXLIUPWPWv+10KT5PXigGkgIT+zOUm7D6uefZrVkKUX4md4o
cTKrBlFZElM92jDkjS4qygeTHU3YDkfucG/LY3jQlV8lyIONP3tddRHZFaXLxUAbSVMDfjAtVOl1
nmmm4gI4nDDeHEbqgvHLY1kHasDFzZ8PbQelnS/As9Y8AiHjUmxGnibPu3MaT7viJiVkJEvN3dqx
Uxh573n0EAWe9mwdcMkxdburveMS58QJ9AhQdhZPpaFkaJF5ItzhQHHL5vTQIyEuhOVyqP/ghGhM
x9X4FrDQ7roS2is7vqp4wFMmAFacao+DG+FJIllX8vxO9PTE5NGA6CuZiC9ww67TVeX11tFOM37y
I7nvyT8ZuasVPjbWH+lKlL57i4y5asUZ61CvfcyK6CwkPm7HHlRouzlWSS5u+7lF8crVO6nG5ocv
46Re8F2TXZxI8Y/ebRSGgujBfsZn61wRwHC1U9OssP/1ZDDmZOj/xX0uLgWO4Zbn3rdqtXqFyAZa
CSe9Ym6VHMn8uV9Cju2eeaqdHzq7v2aDqtZuOKlez7QnrTtkSfgCc7L/wgOB0jqSnKGF1Wc9ay5M
XfL3LSQQzenq0s2oh3UJtbv6FirVl6x75MBcrUbebz1obmJrljhI0cVIYA94hkb9Oi+7mYubwoHM
HRiL9EjiiZb0X+EtEe1sRn5dICPFEDjv/wILW2ZwvjK8NObGtzQmgg9MyFzegPczj1NzSgYRh246
GcvMr39aKJvTYra1tTzrcQUGfgF6cPGFWNBnVTXyu5pbwwx3dOe61Uz2ZviEqyR+Td6gsNseuK1A
udK0DOapK7zSjEp2G0FQ2IuNxn6ZxKXwkmbILUTIVY8OFrWBiMJsUdWyXGk6QbpZuEFeWvwQ2B2d
iE2vyTLRV1e5/m2ZDq/Kb+wN+4VJsaoBQzsgPHc9m1OAv39lnmX7wDdkJAWGAEzJZG4OGrU6HXsi
Eee7mIsG+qCdP0vqM4MGnnsO5RosbxNEkA/aYKR7RMPwwIL4bo5LEGJ3blGoWNiGeWq4+hgPKDoN
A2fgTASQB2IyHC8po+dJ9yD8PwyK1RmlLguxtPN1Djjufw1zy5vC6fug1GAFPM4LQUg5+GdWQBfh
XodLLXC7jlQs3E4/rzgPvRrRkDJlBXX9NX7eJf/itLiGoP20ElPDeP+S0HYp4j/V8bmLvTp7s6J1
IhPHCJ/eUGIwNwvfrc8qGxuAp/wCbkCNexsPWbC8zWnbiVnm8f+9dMFNi/rVvbgaj5rosjZVmQl+
YoV+IZUoNx9+KAvrQUv4xAgINAVVvtgntCkLywylrToKreflvmPvpP900IbuhVc8YWQUrmV/UOFA
PGZxTqtmcZJ01T6gpyMTey/VoP4O8RLTsQo9TUheIFfyLjXXV59nuafFsoQj6CP5GsAVSeweI4o7
MvyNWI/ROqRa84qB06344R83O6d8ZnI0P6+Pkq4dsDdP90dsWc9CYO5kjTxCL2q8usdYqKq1OYuZ
AxNhIpzYt6EPBj6KCwH52AVx8XB0Nzu9DjdrIbzsmrEdeMGeU0iBDqNnGTFAewLZWTn7Iseb9Jem
mDJITs7+OQBWufhya706wxrYMDPFbCxJJhUWCdSAishGjuDrzX8ekXrPEHA3pxiLQwNLGE3s9XMC
bDCVsiBOuXB+n9LvO+x1FlBrYHJ9B6qSyfmftUJHnHI1L7D9RxvI9wLVBhbZBP8vHZ3j1QUNUO3f
cL2ndBwfaud39eAcqocfICgbI9xNN/tBjRa4LKq6EtY9x7zmBivrHpe7qeNMaim0Ql2opFknCgWs
tjLvzIu0wxd+9rAfZQn89ZUVuRK8bykm+eW2bPT3cf5lOhGmJbt+hRL6QdFqHYu4L+hsP5JddwCA
3T7DdKGyCOBew6PMsh35e74+7gwE35pKltMEPc9b+f2UmfDFXCCQa24SIkmVklFvG1fRhqOZqJnn
FMIfehNYRYZcEbE5wCdCCKTFXciZeWmJGAnPqdJMuU3IFACZjv+r2CWCBKjNAKiz44Np9k5Uz1O9
5LQlUQ2QbZZxH00rBWPvOcQZiF5ATDpkXRcJNaunf7TJvOJYIKGtfVv0YO2kQmu2UKmQRbf4rEyl
V82NfVmQyEM2IDf0HrNrDWdcb8ntCDMcoQdgR/onxwzRfw750XWAYj01xog+rH0spJtzz68G9HHM
38mHMiAhGp5BTaqIvZLRiqff40Ct1nhzCqj4iZ8LVFXpXhDXLJOAEfJsnjMPK0tjvaXZ5cJ+gYYi
C4GPpzkmTWRQKQjVYHr6zwNth2lOTYU7Ng68xeuelJs8RvonpQ6WIzGytDuPCieE8mOxEHa1Nnw8
kGIZw7GTGcwTLf4yQ0+buDaUF8Qbl9EWq+Wn9GegjCnb41LfZq6y6CQvaBeLNk3jDueW8Sfb2YBL
+Aj93ri+s5K357PRFoEkN3UPtcjGWkSdvyy053dq6lgD1bSPp2LX5hRwiIbHg+ErBS/0dxqqG6lg
mtt0NP/L04sHTKwCJJoRY1H05EKDDBonZUhQElltG1++7hURmyNJQxFe6fTNA1ZV8n2DCB9S/weq
1R+NnVEtMz0nhKrcj/EQe0P5ZPsK0KUQ9IbuPjfVyoSx/eW+UX0kaKlOA1SvzLBMf1lCInhLNRnW
ezjUtUtcGY9k1gZvqbx+LCXGaJQ/P+XwsWjaWckrOzG+kOQY3Z8esQtJPAy5EoW8T4s8hASVLy58
NZuypSp8MFI6wIu97Zgt6sMgKKKoTw5hqEGgd/kTgOsMe9E4XS/PpwZm8g6+L6FpfmpWVDIvrxfb
KlNIg1Jg7k/SeIfOi0+G8Bno61oiQ6xfEzJgaOKA6vZ2oAPi1VzODTsK8rB4aJLNfHgz3Rr5nrht
7nz8pxC5knAE0rwkM3Mx2LWKGkfplxzCMjaNeeMu7dgNNrlisnWV6Kn6+IMAsrualsLAUPJQLZUk
U52TLvXWETr2yftNoGE/BSEYEca/EiAzH+OOXhQK02TnVSK7F9vqbFSJ2jWXyh8zaM1jkkmDpOvq
/Ij9sX1fzhlKft3lOAWXTphf6OL9XkjdBnZD84xdzPDNaMGDYSXM0AhuRIdSZGICatoNzYPxNR7r
OXiGxHbogtbAL31zk4aRBDej4U3CtTsF+WTNcZg0C9l1xTeCnYw16PMTYoCEjbYqZOYVra4YNve9
b1k8fWyvhkjNegb71boQpXc3QsoCWh3LJUBP0PM94uo3LhFCHye5ifdr8mWISSlotJHw58hGDWW8
gvykcXQYwelQa0Vqy0sonXXi9WnKFfxNcpIJRR4ayNHgO8mtWLjDPONu89nB1fcnM2jTCRrNFJd7
24Ftjk/91MxopavWJTTAt5EOMYRJoA9LtCxwfgLXhC78kGQviY2doHLj4vUWy8VglxYq9GTjzKPV
rV2QpyyTTSFk0V9m3oGtvuwlwutCStgV7FvSxzbNr33NcPA5LC37FwdI3LKGx0iM6I6CvSo1BxLp
Cw+KhW9G31eKdAougx1//9r5ka3uKOfak9RHF4hbu+M02B0D1UyP3XLGoBtRmLeT0WjbfPTFZP8R
kd5IQTURkQ21ewwNsgjpfQGDMIGtbtjaty4kUeSbjJdC5FEG4KP8GzGiwFBQHTEL6cvFatdQbNI5
Gujqjg23nr0KzVzR9xdLGF8dUnIDAxhEcXIzJNQPPHcWrHo1R9emoTn/O1NJj0S2qHkHNK4+X7HN
718SIt6uYM9IClRVjpQ60eQIarZaR9NscYwAnTeckerZL3k2gvLTmSY8miND7rpQbepqn7Oytlay
1EPL84uOikz4PU2hxwDjDPzPhdF9F9bhB1EHclkDzHzJ+OzFWnw3PcRtAzieG/xAWBNYvl9qczr2
il/Ngo566QZdzKgGGnZZF8HJ4tRb589pNTAKYi/a6ATKEilHqPK2/lx36Ez/vSsPWmpfdkxHJCI4
1tueR2FeptaV3vCePJdv7NW1WRf4umblcoWop2ROxExtHXDWpo+a6UJE7Vwn5viXwO3psGyfLgNi
JcVcoe0rFmBR8ma5kzuT9qSCoZlYVzYeGybMZR89jyn5YkDrQTaPgje4e8KALQ6jk85Zd2RIR5WY
HNzWUTGeOlmH+VfNsN9VEIt9D6tpQngOBMQygmnkXRxHPtswAGEX7KVFeYvKTBj/wUXPCJl60v2j
bzxW5EIL0jbFf8Ao11uW833BDruZHVGvjDdtALM88nVF1XRXcTD3TbN3B6vFjaE+XZelLhwuRsUY
H1nQ1zHKbFPCGBepB86fddCfVPThSeTwBhRHkxaL1/jDOqwYd06tWJwTL+lLHgP9b3CukMpCOhHw
Q5+PoDHLeEaK0vCLJDrJ0gCq6gGQpyHBPp8h6rSE1eJ1kL7UKK73+XUZyVjohAWOZkQf9yXZQGWS
yXrGP2iA+H7AL2ziTKLY+jCZCRDEhZYGLkcRFYBHYWu4fF+L76g7IgYMKxXlU4LDPQbwSOXgPw0f
5ZvNxg+7VtTXx0imjCUomX14SheRVdIZZZgcHDAz7sV+w3MUP64qvxrwEHLntlzSe50UmX45dA+f
6qJcn9IxezsL8aYKT7kNhPWp7+Ony7yfcHlQlYAVWjsu2NToJie+tIBfNPOB0sjRjMY+38V8Mv8G
OYrohzpzX1WfI5oAyTCUYmZCkKxzPc5mvut10hbUzStW+wtxoKEPWW8WQAMBYfPCPmzoXRSePgp0
4DszsvdVbA9xHjg6cbijx3KRPwGH6nn9p6voZyRE6q056iP6XcN6tJ+cBEWQIuOnJCmzsqRMoQuL
XehnV3oEkchXwQEYwfcwui6n2dErCXMWLjj8Tx02tY/pOV10p6iKLw1ltj5l+PaRcbvOcRBQZ4uH
zoUWP+NKA5JHuTANOuRGOfnL84qEAs3vyMMJh3yJfwd1XFhRLG6pU6IP4pR47EFIDMUM8ECUqSEu
232s93dYHW4yK+nwBeo1KfH+o2Zk3oFM5eh+IqxswwtPfLTJwPgRsC/zZrvp99LmYi+eJB65NVfh
loIcXfIk2WfKyUpAfSoVYd8qvya34ftBhPep5P6Xfn/Fl/j0Wejw2tanY7s1eLDXuM2+izRliKK1
y+nj/BcH1TIMO1AttD9mgR8cB6NSrNFbXP0S6IAEy/e2LIq6UmwEPEz4G8VNIQMdNb6fhT8ZBTM/
Hha+GfRgbBjyadrIPYDMoaW13tgwnTYzIxOTLqrPTzdOLL39gvlt4yU24/2pD8IlzXjhwDGm98+2
f8U5LipDZu2S9SBXbTl2eeAViTmtYi5VK11Ue9iFngr+ijFw5mPodyqeulPqwxps+FzrN52fvkLZ
Rck6gZ2cVBCC3yLxTiS1OmUYGTSo0zPiuo/x47sNNENLkLrA4R3LXEndTIjZKX4yIAhi06h+86l+
56r0ynL9HEv27YCz9ngJI6rcgi162RMtFNY+ReeNjllEmOUkHmBNuccI2m7dBeZddfKRkrZZyn4x
PGGUoyKeUZDkoOO48jSDbHJoIQEr8r0GorgpHA9H5NZwut4KyoDARIEZ7aq5sargaaF6SV5VW8iS
6uCwnIqqNGExojP8WyIUr3QaHG/RYkqFFA7rPHfRfKiMHLhD6n0WLuzcpFbu0qrezRLqtjuI9ZWQ
f0AFfv98W/Ad99ADGveAvz1z/xvTnB6f50xgeaCbbGtBw/mS+LOehCMzwzxXRgHVYqZiv7oRHAAB
iKgmbxz2gFoHReQQmlFcNyxL4+Q3Y4HxCj5/hfWfACz3NmGk7gJ3lL+eSWYMeG/HA2i6iqpvEgK4
nJxnP6TdryFD3FIzYoB72JMmNSwjiacI7aA0mjEgP9sqEyc8DLfSHktrrm4JL4Sr4gyss1nV9a3/
wUhC1jk/LCcx+TV9aRiFQqvFg5UtLxGVH6yuLJFnoNhN59cOTexubSQSZEtTjmjfw0K0s/BjEfPB
QJG7qB0XpCeCMWakgJDthHhTmjQy5Bbr2YmhFSYAt4CkwH7m5Ae206GgHWXVYxOgugEpAta346kC
K1NGRu16jWJXQjzS7roCZp+zlbJ2mBAy3fYXxeF1/Nqx9IvmlLNVk1FZfIa9OWhafbwc+g87pEDK
t6hc/IM7GfhkPdnmeIK6Nsag/dlWecKPfIjI8ZQENqEJbry/cCTxkRPRflAvwhkxChJ609XB5TsR
O5TQTRgR1E6xDWhjRj5Z1L/Q/7WPWn5a+bFhrDIN4zZG9khgy4IMPuW2+6SlYqyz7kha0sRDO+Sw
fm6lAO9jesX6dmJPBlUbhUBpJDQLjl/rJzWenIULBdIAxKVWBjizNGLnbNSohaQpc3/dkbYf77M/
+2LnugiZF8AnJZWm4wzjXqm7YtaF8ZL4e7lwllTT4hcek+dinYQJrJ1wS8ikL16ExZ9XcON+6Cis
gAt+qz7pto2tlDGtzMDevmueCZlEk6TvWeTVwAC8XY6tydNKDA0H7wkBlnO23qfCwl8JCyHQMjnm
ywIPp5gzI7LhwClvZACRJiGLMVEoEmUbQufSZez3kfLnC/wWYE0t5Lexnh+iL3JQuYoeB/oKAEOt
7meb2bNWcu6mT5FQMJRgKyhkwJQDc6VZKjshJ83om3DFguoU//w0z0pGv32LugvIRFyQOgtzdYNd
nSajlpi0XzAncwF1ts/eHiNsAzY92JOk96hngE0WbGTvgvffdwbLu1PdJZ7v6aeB9dBncngBn4I1
Dt1if/3ABfccOnI793KufJuGqHYLYoyFaWKO7oQxWSuuxf2abF1aJOz8x6ad2H+FUCb8nuo3QTRW
8j1dCzT5PJz7S9osJyG+IQwqD69dbp+LiN+raWV8T+q2UZQefSVTgMJWdBFx9HFNpjth6U4q7xUo
40EH2YGdsuh3T9IL0HX5CFj6FTR1jbsCpwqbbdlf/UKwHxfF4TVHhbVWnW7KiRcyEX35JvFu1D9X
MotwzQ8X6AYnY5gUx5KJXUC6v5U/o57cZe/5ciEZRiUgqJt+yatEaYwS5cIF0RoTJGwkfqaTSaEo
NNVWsF4VbdRrKMO0STrgKC2ZLIgOKOdblLlWczMZflKdrY181Cw02rrF0dPKb+uziI+lvGsOP/gH
/MBwAQQLe3SzeDElmOlM332o5mgvNsi7asqEq55EtHop9vP2NYjB10smua/DYDaWMqOFeJqt42k0
zKGuzTa1pwJ3EE7fbqqb1BK3MH+s/rKSRS6egu9R/DenSTzH1Jibmw/TBh0qMnBeXHau3BLVOhDK
CpdiiA20q0cWnlGgAcSoyCpFEucVavIynA/05KfEU44hV+WZ9BGO9CJU8d4YGEDPHxS+B8uGAhHU
HYQ0rWr8sPDjQNmCCos4NsuiRU/FVGLBSKTp6Da/TLh3oOVM/Y+jyKAfurSe6EdT0OUSVJAk0oR/
QgMco9JSYQakN9osrqW+QPkvL2FnIfheFOPNLD3yXhF4OpRgDMGhCGXnTkVKfonNVHGsMphpd0H0
4WexswJtZT1/qypIvihU4UJ4tbkS+iYNe3xhpHh7ngUtnOInZE8Rj74z53yn1ZF2Ibl2303tr7c8
K8IKgZyvlQrXemAFmfvdha3syYIHyKW/I0LV0uDBDLoXfny3k/7imq2/ZHFCCVArL3LfIH+gS+Ie
U+rd5yqg6de6ohg6Dfe3YPyIfHbU08djmQWkn/PDwMCwo6SIRxCC8qLCI2UeALOtl2jSz/BrQ1T4
KvFl0SbfFEzBOUpR1AsvEg8xjlzBKNbyTtC57gXgT5iReR0OH0RSMwutpS8PMRj+CoZzghXwUHXP
t3oqFAOzxu2w2o+AOKN8oX9/5qqL4J/CIMpKegR3j00rl3dPSVmF04SENeNsVRCrNTMVtW/kh5EJ
1VYuNnN7tdBDtj6Ski9/r/OiaFXfYFkQnq31SLbHYEJluEHoa4/d8wxX5fBib0G9tf0xQ9W7mczm
s9yOuZAoGs6M0z4jQeQ2HZ7GE1BFOi3F/GUTzofxj/jvgooDviWU3zetU2FnKA7Nb4mKdrthwkr+
HT/Q2trVCh5WmJOMtSZbXU65DmxgDuqb0wcS83io5mLE44DKoVjM4Hvpq8ClaaSE4C3sXICJRa96
INM3LQLptRmay1HTML6ByPpCJvC7PSqRW2t8b18vxde8ywQxAjUPP4EnxFAT5kntbuVU3IlDR0PZ
AazMKI8dadBNsBYuwCV4Jh4OCJWZn5cxc4v/wlVgoOoCWF7bDr6sqMs4mzPb1w95d3ta3uQ0aEiE
jV/Cjqs6Mv3qEqi3Yq5xRbFUAqMEHlOIvkvVS4BgxZKYbH0u5s/DaDm6DTpogb44NBHYEBQMmALv
PIwJK1miqEtxjB9H6S4Pg8u6Xv8DaaYxodwU4uE5wkgDwZq2Xh3g157EzcMm//5siQiMPu//H0Jp
g+LBdZun+p1fPQLCGB2KvxeU8sfqeTW9VxsH+cRtjsHYDWhEDyPCRyB0CqDTkJ4nCK+WbIux2K2M
zSEI99e3wymBFb66JGYCFiEFkOmRCpxISPoTCtlpyy3EQ04UvhEPuyhJ/4HLOU0rIWGY5Mdden3J
rX0jTYpVXfxDFbgPb69m+8tkeDVOJRyad002W/2VamSyk4Q9mH/z9G+Hu2QdbW8ca8dYP7T3CNM1
Go3vQ7Uoe3ZG46upZrqk4kjnff3X0mZJuKjoA3/6z3kUWB3+DeNXNhv2Ss88jq7QBvgpethzYI8/
a5xu+2u+GZLdz1ROB3fI9paBxw6GWKqGzA7lR5HwpkWhssCBbN1kmrB+fEWmQCLLRke/Pec/uoFU
y88b0Q1Fqaq7x6Opyvy7jqoNck171vjTVTN3PkM+3ZGcprliQAO2t4Sft7Am/V9/qTsqi7mcsojx
qBUMc8M2H8UYfJQLECESQhGmQEnZKEk0ZRLnVjSTjjLLtjcpW4jBcMjHPn8hywv1omyE0EEkQZuU
IcZy7+Ft+XXI8cwXxdBnM5fzB8Y/ydOoXLQArEh/zO9JLh/3F0m8a9xb7IDr8x4DYjARi/b6p7+e
AeV9kj7hWT31NjfOVTmXX2xf/UpXm66Qw9V/KjjHfiP7bEKGHzWEStltKFZPBR9bNS06hznexqZI
qkGgbga6K4QoQqHsY95QGHRNe98efSaXCLbxaSyQu+koLNd3PMo/Vey8h5VZp6Eh7p9qeNMLB/jX
IU6/g6YiybVzpb7HSt90Qg55hEqfRJ0LkfbAiAN6v+WTrP6BTaUy1trAAWDGK0nbCwn4qFQiWZpH
qZlCGxaddVGnn+NzV26Hw5DegNnU31LYC1ZG0RTgCaNr826zUn6zJrtCKDvnqvm7j+cRFO0y0vVN
fLTTGvu9Pekqih1PLyfjX7laCyucZY9sQDlezW2eLydi/uz63k5frnKw+9DSiytbGyXog9NQTA1x
As4S/0S7hhtk453n8wgWsk8jzPdY2SBrRkI6XvkcuugucYs+LdNk8F+6olN2MdzL8s+cCf+ww2z4
NhJa7Frl8WxiVdeeKNphUXkBxHuU03j9LnDKOEPjyZnr3FXzRXFGhEicLKOS1XAR8t+Hv9Rb8Bq+
j6ZRJzQk8JOehphwbVdg5Lj4PpeWtyZphBISt4m3ZFE1bCFFAlhBjPDiRcMpok0gxalOJ3L0ukzZ
MC50y5Zp6W1/awU+KHr5eeePlwQnx20szsUnltTmSOss9c598hyKXhiM+9irIX7CBfPfgjQ/65hC
9TzhlVl4Hrv35jRqcWGw+Ppu5GvXApjBRpKDrDfU2gS466M3uh0msDdysSG/pwefMAT7/f1Y9P5g
rEY6aAzfh/GFuCPdI1NZxsNrTGk7q5qjcMicmtW4jkXB7uNxmFK9s2pgTC5bEvlzVgT45WzJqF6u
ZUriSnzjRyoNDBasV+rDEyrPeCvv2BZtZnXMUdtXuhi452xJxJPpeeFCapMKx7K4iEtp9VLWl1eh
dHNbjWGMicO5NwP4UlXHt3aCcRPhV9OMYrMRkwZrSw2dG8VBe/TJUDkAEjB+jOqMQY+I0j4LTDQx
ZOx2Wqgwc4zcdKqbxco/bYABfZlqXAKt4qbIj/m0CRRPJF8RFuUli1MjSDBkrGPct8ghizZWN/WY
CyyaapkVwLJSSm2BazQjTgU2ErLLFoazp4HuL+EeGCQ2OixzSt2AZVvGv3AUAhfb5/Ek2JfVUbRu
uYremwJmNsB2tvxSeTcl90TBqaZNyy1Wg6Hqj+wSmNIUuatRkX6+AA8Z9elkTlpbxcAjuzZ/49B+
FI0ExeBRDIsgkhAdhzVmFXGU6Rm8QIdflxQs79gz+DNrw4Pd/fkhy8gdTdJ9HP41VUa+volEBZrr
FOJzkI/RZ4ecJtpOJfUHj1OC2SvLBiqP6Bqg05B9Qw5FApfcf1LfzvTv7f4DbR3riBOf5lmyzhm1
B4MkBLai5xB41yNUQGTtygXLWGyFVidKPWP8xdbjDGLT8sOfnWDsNDjaNp9ARiVhG7FusyDua4AQ
q/5/IJ98aD0VCDLBRTY+veIRmBLbEH1p++YkGlECMsHNn5d31fAZ/g10rExnQGaRCZUc8+tg+F38
TGOMtfXu2HYPkbPWdKO1SYX9/WCrof88QzDQ7+m5YLmUcQUGNTVvSQSYTNQnkOJ315Rz5Q/DOOOe
5wa/5fRs7Bym2HxIfWUs4CMiEsG+BiJDUK0clSIXZiccL7ZbW4tls8+jf6nl0IY3mqbDOetZ39Z+
fiTwVgES7/AiJ04lksr4+5nNhGSslAvlH11am+V+hB+/cP2MGcYPpvASXkCzSib8BYJoWYfRQ8ZE
kOCMCkrpK/rFo/VcopWWG7r/RHlCHPYrk86oGEKZ/pqGQRwLEKiY7hqPRnTGd/ARoVgNVvekQWVg
Ah+JtT/ulnKlkorzxAyYM8PsxkswBiyaGY55u5MlHrMtCUyOyJTuvfTQL6qEBtKW3FZaoS04QiKI
coH60vwrxIxabFlMnDC5S09KEKHOtO8hma1v7q0RcTbDLApktBs344TqIg2Lmk+Jhb0RxuC6EOnZ
rq7MUBMKA9NbO0mrn8SG6socIKXcuR/0SP0unyD2jrZdIWoHjzXJqIaY5cdnkMRSBRNre4AqZ9xc
Jz616UPF0xj7z4M/LRFCfGmk+LC1BhCboN8lXqGy2viCXZ86YT/l8lY/9/Z7nzMzBuVbUTprEUlj
XV1F/PehSt/zJd8ZdIaeXXwGEoBbRkTzhVif0E6YEgpo2Y8LCIfR7kSOehXrMcxozrw1Ryw5ACOx
OsZWr3jzLrK1O1W7GV/pxmXZ4xZf5SZdozJtXe33IKd5DmNzYBek430L+zdC62SWPOwIP6YlB1D3
R3U0bRqBtrqlkcx66I8Bhw8V7h7+DPKQcbu0BJkU3kbxg4QnL+B26U8k8FPWtDlVsX/pHua9vXd/
qkN46hZF0O0JqIlgwfyY9KQzLT173A9KboV6c6wHq0fenZoCdnIQ3ats4vvF58w2rW2dfLP7hF3G
qX5vlx5rT2lp8o9Wpr4oCQSfaMbnhOOABS2S0BmCA9sAneNOr1HHFG4G1/uvNf4v4v2kHMKeL4Wa
33wqK6KlSpGr18WUuDv5MIwVCb2ectT1rEzxkcndqkluHygSsoS9I+MDToJRGV5iyrNBvJ1vhgK3
s4Ine7c42YNyY/YpbiHnuwdsrHOOFtf1qZ+J8TZXravn4BbqySC413cm8uKtVjrBBuhTwOgmD7Bt
+n3whHN929EnKhqiiAG84eHfaXLkZ1csmUCtFF51vDQjWf8kJ5Rm5Fqn0VDPrXTFOtjLWZei3Wlw
YI/5S51SGI3H30+gzvA00YykEHN2WZ7l1ITIvg6feVWRNp7JQXSdUPM4/CV/2WZyYdRA0GOfkwpv
PbYQnIbspVqqFUKrAr+axMy8HEulElDuhKSxrorpwtLPko2kcpcv9EQ+nJMnmBSEa6Fht7XZDsSx
x53/qR2WXgF80qbNF1TgQl+4EwLeikpw9gSWiOTvYHLWL+BnEwqp7obSlPTD3r1RJ25YWAYK703U
eFbM49Y4+TrgQu4EchwMX6163wbaGseUoOpLqd4+b5yxJdbfc/hBsdG6zHPYVjG3gUDHjgOSo++P
MTQhch2xF6zxINEx0S3vzmjI54e+Y0VgLTCgPkJi8xlD419HkRzJ46oGR0hMyyLCKRHorSS/vDKl
vWITTrwQVzUu4f59Wm2xfG5Q7LtWjij0fr2/QgooSKnmQR/eRffRkPyJXgPOLjlubXjmA2raPmPG
DA7nwohDI7RzqCQQ/htk+7iAmVBT4uWUvpRT9W4kubrPwAy2p0bvRnLxxuant9XJmOTq8dxue8Ek
CxMo27oD/t8zmQT8ddmczazLvlwOo+oZW4rnr8Sv7fh2XJ8xeakoBDG2qsyeHyfT7BgFJZWub+Zk
F6Vyq214DAMLPryiGiDc0cB6+0+4sY38P4SSVELilFzgnF6XCYaDORF7oWQBAnjpSEk7v3P/ETCN
eWMzC3Ev0SdrJv32Fwrzb0Z9MUjbVBt1RrHL7zizEnt+ctE2Y388sw5H8Y1CGxX2nBt8m5FONyTf
+323oU8JknhbCwa6aucW7UftnUSZ/ZWvjkOTR6bgLc2wZe1N+NK5GxfjkJkVEzbshInsOuzGRzaB
woO9/aLtRofiPg+r4awedubd3EdgJCoUAFivUIEysFvbf8fC1WEYBuKoPMi1P8Si/IPrSF2tZzoJ
oZO821IjyvCM3lzlJYGmlK3cY8xObvPlJay4uu8zhjne9lE0CfvWUuux+nviZDYNzVcAVexLj2d1
kWnHpbxL3+x9ncb1PZSzNs0vQBQEtfBSruyNjdonh32QGI0n+XJ7lccjhidx9mlTwtrrOtqw2nM2
D2ZMd2bkAfnG5fS++YyjyOpV4CXYdyvNOMwZcGAJyErjZ+rUSUoKIklS8erbUvQ+y6VXKtlOaWSs
6SkCqSN3ZxKVCb+IkBs2Jm8ukkKnbMDn3ZSBpP0FNVmU1Yqfmnh2w+cmApk+2bCAk6Eq0gR7CiZ1
LgeVyyBxERKpz3M/iPrP2PkdVW+Ql/0xqmmEJvolsSHzurNoO2V8VDWvWE4DxDXmTDlCZ5RdXaC/
QzVU0kn9Q/cpfWfMYIiZrSuylWgJScicdUUFqz3u/bf4ON/ZkIFV4chFNWaE7F+dLLba/oUl02cg
f4FM9Z4p6EXR/I4d482SIR6VoYJcvQSg0wsB4IaIaH1h5fS7k20Nfymkm6goOEsjbyFecqW5D4kP
Lf4/wo3Qm1l6I59N4ULV0FvkVX+ML7xEqTHLfM1VyhhjLWdD7FjjBZNZZzOE/jahlZPHx3piHRRQ
qSDP/E4Gbtk/4aowlnEeqsIYmmWcCJ0a6rG32Omg7eoWy90MUuiRIA4pkv3yYaYwy4wXUnQNVmB1
ACMF2rrvoZzhB4Wuyc3aVhUsAoFVbhQI7ItFFaYAV+5hLVw4WTz0HzHCwueIkXCmCkzAfvxMuPca
QnIsCuSaVdrU6ESyMnje9TDJupq4cJozL0hmIA+3AF61VXo0jdcnery3mZY0eDI+pUrNI4AaStmy
NlgibHUWD1woQ0EGNf2pNrenS1YKataJirtL8KPzLU1ssEvyOZeGvby9MdwefSb4e2CwHJDFXbcP
65/SEHDGd+Ik3EFM1jHUFwwMtnQwVsVp+c948kviY9EpRnQDeby08gIgQWUhvW2wTfrUgqU8iKhR
UMDuJ2Q1usVQPROnWMd+5NQ23wICRvsysK2Gm/wLNYdE0gQDFCfBlKJ0MsjM8OSpPN3nYTqN1Oi4
wswk5C1z2wRk1iGG2scMupH8Wlzj0m8ghitT5NoVpSluiY7lk9eu9vuYtrVHxPuUwifiv6hsxcOQ
hctFa6wmmWo7rrMi+vy9idctXfPwpjyk47BuXhwNBkmYZgwzM3KnMtUUEBiDnDW2qSYuWsuq1yiv
IdM930wxnVqZda7S3vUEJalHFwV3PPKPvqWZTI7r21R39da/FclIEarJ2HKhDfdav1XNaT6KTeNc
VZZES31MdhB/EqS+VANWzT7vCVy2IRh/2HBkYOu8pi+4RUKmQa5ZKOJfFYlV9EquHU0bw8hyNFDh
0HNUvoXcas2HoAgRYbytLdEYFBKozkdBx1XCUIeGnIRMGPGXAFR6CozlfVyP5M3fsGPFQ2v4SOUl
jyPjr++6pcMgOeKXcE0Wmbl1TLrJEVTlOjJ+TajCDCH2N0meCqOOIsPblPojMs8jxZ1+N/Rz7rSV
0+C5K4lZcmqPnHL/WoLd4Wy3auQ9DDN76A0Myd7BtpF0rM3NAUnbso2gk9rPoDrNWJGTBKwfqVR/
880rac9RVQ7tA9jy/CmVZwph253+w7f9C2tRL76n9BQZHsp9Fu4XQH+p8Vtc07Rn096mrI6V9//M
Cg9oUNwImbSLmrL8yWIOE0S9ljvWCtkquR0TgRV5ycQKwDHji5lK3nusRHD9u4OOWcSwdEQiEgcr
wDs6r8DmLGOojjkKP1rVC0LbzD5kb4m0TtlCZ2Ch5kkqrGWrOHADts20GsLIe1mfuIa92BsHyd4y
wdA2y4kCbCnl9hSY08Aj//Yd/3Gw3cW6P+8GbP526F3hC3GKszXxF9LDKMspvWV/+Mg0OJK3la/2
uZqXXg0TVZzaKLgpewu5O6Amx+CJQ0ejnKSmO7VClA8yRHohJfmmIg0u/CZ1fiWXa0uslLVFoWmC
tFxzBHyXW7MAPEHjaKrbXWqQ9Iq+FaLg5zv+76McsdJS3Lfps9iGITW/57dJWMw/tEHh5SjjrQIW
FC+xxz8mRtoz8vsJtiYcAhgJbuCuw/LCF3QmIJ+daUrvl1mTZqMvBfmq7LXitJxYPZ7kQcyYzhh0
SAFK5hJAz0Nck+NvsCkYWq5lMjv+S6hOmjxwTaBpuiUv/OCHMqtjqOoMrqGF3P0tIYtKwt11tpdj
zwe9otW1fEwLJDk6uxDJwR7tproD2Bbysjh1EKD9+feId/FV5cEnVNtm3HizLGyE7Ml86QH7IhgA
z1bAWSNfmFsGOHmDGrZP/Tr+jNCCemn/20gaMjFLVNo92b7pAbnGcwxLYT8EVCV3nkAzaJvRWYrb
/0odgpjGn02Ip7dF9nr8sPH1TwaQb2KnzEsFWMwGMnJ/A5v9f1DeYMnlNLSrWtAxJd9ETrp4Mdgc
uiYii3rHzAk/bZa0BE5LzkKsTMYPB7CkmyBR2KGtp1nfRQlqerf4BGmf+2m35iVevxMUkdRusTcK
V5OPqly9hrRqqOdNBJWRmHAzshKNivBFqKDhytTUuXvJ1XwCsvKhvH4oQD6YSahPbTqQuUHkyffV
qJLHf3/c64MNKJCKkMS4GQGMerkwbscHv+zOHr1xH2SEKJTxpjyODE118yKVgFHttI8OB7Sb2XQH
izBwD1+JJYLzpWJ1dDn4/iOFY38pIkhUl/E+0OvNpKsw5XECFEqFXzTHNVnLDYupBUlCR32UUDD6
fpA3nqrDJHRndPAOPpyV2gJHMGLRlySUW1sDEREl5RHZ8dpUtM+A+J/xqKagkaRvZhRPChNIPfOD
gn3X1RT2PZFjgyL45aSG4jEj2+4CiJL1C8tuhal+ehbfKjoCYNf+vaKwtca86DuNqyqb9ppjC0PI
MpA7vrRUXfY2+lJEvbu+BwQSD65N5Mhte1bQRN4Jkb1Zuc6TpdVmGkUoYrSTRq0W3ZQU/xqGC6Yb
UlRUApxJQ+cvp/3Jw1kK6pu5LPaVN2FTDf5WO8YY6iyK+VNj7kK9Zz6+xghYsatQyxDjSjgbqj92
1W7ADzpHdYyoAY7W4Ne0DkbLdPSqD5Jkkc9oFDf3+J2KncRmUqbq/hpF/oixRGdhF70LLFREoNe2
pypYzuZPuEmoYST+GcTJwDn01PoeFSUfhxSdG+p+dxj/OogkfZO73GDGQgJC5FkVVbGe8s7uO9t8
58Ug/nqbJc+cIOKP1w+O5gRiLWE+vKh2RMACUUSLZjof8R1fqeShbmD2vPTipJ1CRaJ6zU1gaUa7
gCNJhEkYEtOUPNtiEbMZIZCZ9FmBgcCoqa2lcm0u/oAQpOXw3R6tIro/cV/ZIWPfBb9iooYsKVKr
h8QvFZx1VduiZaWB8NrdIFEdIFwXt+RhwSNzxIaqc/+h2xQL7udg/7w9s/S6bZWD0Q1s43LheL74
v8ovx8Vme+LLY0fwiViiRWMoqn6qm0jA1CRWWy7WKVVsxvEZGvOtaR+OAUYZbCwFOss0cXOICjDU
EP75Wppn5lQIVJHerYLl6l8er/8KThWAMDvm2vj7awUSn3+gELWE4QHI4f9emMNLVKkW11MFhkdo
PvIykNHhDFjl1WGheZfN8zmckHg1+C4Dtzx24PyXTCkJAyvV5dWaiyo3aXK1gJuMrsixl6EIJFKp
ToLqoklf+gR+kyEIU4n/0CQIaySwGWopih8U+gn1TODo9AzNjQGkSPUEK36V2D/TCNjhE5k3vsf/
Ktwy13Zi56uEazVqHezfXtPu8KUqhW2MQfUeo8AGZjrGa6366XKuTQ3zcfPNxe5lPJQyIcPNv/Vf
HcTMWYecidzaeMZvcM4RknRBJ9fnizORWtGGOot37guw4IT/byNzFJBpPTaLLXXCX+rKQ+vr3SMC
yLOgsBh5sBH7EXKiVbJur+WeKg2INNrxokDpDdFIbaWloF4WhNFI1ZxqvwU1mtX7bhls3Pm3Aels
vBZYWeNrAy7Hlv5WcvPyKyiIMAQwIbCIJam2NCE0CFhKBUowWDyMfgV2rY8vgBTEu2IVTpg5SAFG
cwIxNXc4Rn3OyL1ue4BIpUFzsW7lBhjxS+enFIs9KYsKud2G8RgsG90iO/uky3mSsUNGgbZSU9h6
4pKhUoCKNxWaz/fWulb1MdTg7PvahRTKA+4JPKNiAG0/XZC/dteytjBhKtTN4X9AfUt7ke8KcLyh
4vK40ksQ0aGpjeL2z3d41riNS5E8Drt34BCn478cXAzG2KpY+TRb1eJdglUrWyxhQb2E/pxBzHqs
IbTCXmbpQr8f5p5B09h+ZuvtCeI/g2Io3aZCM6Ay5yOVZoIDgD7hxiMjlBhLEn38xPFgIuOmUiPE
HjR703aaKAI4rHzRcWIm52SWZqwt4Y/X8wsWTkRTpWPghsA3ef6O3R7wb71gTyQfA+lUqxc4+mMl
84wPcW/cB1/TzUkOJ/tQnRA1fl2mRsZRU55OCz0gp7f6P8V/XGBFQrzk6jyPAEcEn6/eoCxyKsBd
tPhVDAfNUhGv1YozFLKIY1WvyhGnaLu3YiVMoih0mDb866/LczRC5pWgIhsHb+094IN5/ios+k2Z
aa0Fz2PsMwPazmVNiFo0PMZPcEdoJ/IjeX1crYYUnmDsZDoleVxVPXSPDhreaywsdomHB2eX4M5/
jF8/682X1zFDbqarKz5F5IQYSJOd5uMUfIdTxq/J2fxWe9rBhJV0EpGLOf2NxUTcZKPYk0cUHdNM
+TSjm8V0d8O648Pil6YzItZHGEkjSkKezIV/ouyoAVy8u6UZHDs/ojEKlDpqFgo7CmgyqWwDl1s5
knA4Z5q/SEPC2abIPP1jKJ3l2mL+9px3aaOLbR9ZS73QyL5kdhHbP9paSIpmgx4G5UifBCzhPWHo
OZ4YjkQ461Zr5R/pOdVuJnMsJ1DcoQ1JJ5FEEEcVV91Lf6z2eBfYRRBHzXuZk9GxD7p5azB3Yty/
BTuL7ieNCKBBG716VFuLxxOb2uiLOCMvFcmRbih0mTq5ULehl+4laj1CvPt3jALzh7ESCEu/usYe
Y/7/fdOyz8Lsp2PRBDUr3v5FBZCs0spTbX+26KAoOnCdoZqd/7bX40Tse+mt99VgkVlzQ8CAZWkd
dk5Cpv3ZfBC7dyo69Uo0MtDGGEHcReZ1d7Fv0vTQPuHxyjYiPK4nguMdBWwsOQxeGtKskpRfH7je
85wfgw77poNEjuJkJSVk2NjYxsJjQAlCJ/o2utIvtdF18r8c/j/C2UOKb/B9McKHnjG1+W3olf1w
VP4KMmkPBB8xeb+tB/kUqKCOFQgfo0rFF2lmH8gtfAOrRl4nFhsXMeuzg8y+duZ/0X+q9cPfUBfe
ueX/M6SINmzIQzKWK7aHXP8trcgMKcD881REzFMDcyocfqVKhCd8Sylf8Kn1Hel8RNkAJ9TNqZNv
ghl/Vtlz+DSUcImuEjxAow9mK2NfjnSArOLEXWzbE2Euk0smTgGDiBOHe5u9ycqg0i6EVdDlWFwA
lVmwXkFSiQU7+gPgmx1FKfErOcLK4FcwhVs26jjl24b3JvqxY/ginsuoYrNjscso5As60kpWjLvk
7OfeZ2JjEO3bBqVD5HZkksfV3R6MEaD8LfVBI8kq1c3i+cKm5xpu3afcgYRpUg/2RCkER/Q+NrL0
PMFYnaCeRPv+GM06VfVZ7fqpfFEUSZ2B9MJvDamKjpLObwhIV5hQ+PkteNzxzmEFbi3I02E1xe8K
fqlGkh5EA9NTQLLZUiooEOrcExTpVYzWtworzed1QfpvD7Bx+zfIuGrEY9vBnwVjTNio9REnUqCG
XZy+wr/Ye6mInW2443z2igZ0NWNO6Cu1qpqKqWVsqgOkBAiJ5sdMEC8LwrLpaYAbBpDCCyPMIgho
yZ7W0m3+2+4i4dgQfZDvwg49jH86kaeLNwIm7Mup/dxHB3YIEonWb0sislHckgIlv3tCAT9H9+HH
wNP6hoT2vsccqic/4BbSokeIwiSe99m4vyL6XqB0EvFFkxf38UMN3oSj7xY9x2//VE8OWT41301i
2VnvCr5adoPF9uV9eS/PAUKEqU9FkCCU4ZpuAJp3bF0nZ+GgKYVhXDNG3VGiL3LmIO075klk652Q
xAup9njmwomOYzKuJ3GTCzIHs8JTSfj+iD+5u3Q9mUn38vJqohuMoJfvddkoFMaM3aydCZZ+NuXp
iX1BY3H0hOOK4Psmaw/hWD0lPDuJ4WjRVLhB59QRkyVxNr5pT/bNay4RRAPaGuTEjrvqExYaopTx
Kk0IZ8I3elBjqHf6N+4D0QtHFI6wvOLZCdRks4smf01h+zniVZYZawTBGA3FVeWqv3kxNQd/1fPx
nsOBdINh67vKpUSLhfQOUDU3V7f/65VVplh1ffppPn3tQWevXh6QgyqhXYGNw9tZS0jwz+X/Q+Uy
bj1ZLt27a9NSqMNaS8kqvdf4Dia0m+Sutt6EIOgdLNNf2lhRlQDpwphNa9ZpTVeTzKIyfE1uc3zC
FbR+rf3HysYF9KAYINT8wLkruzrwsQo+B7WJCvO258v9sC2a5sqM92n38ZTArEYD23g2Q0hZWz4u
bfqB6/SZme5uibHUjilxzMN5FfcJhe8JPqyeKs6gR4c8ChRQMtpMoJlgs70jkth+oZ/OJztwDorl
QFv5yFuiXF7frORmJ4F/kCmeJIcttpmXBD83XVk6m/mI0v98Td0OFDPCTZor1AIKkHsDM1SULLbg
veId7KrkOm4DS1AGzoJQk4ijCXgPgvvuLzU99yAIFgs8MnmzrVfGECOCl4lbE7CpOfMafPWRlphr
hFSZxdRn5px6kdiQMTeriinWURg/a0Wo1tcBWEXKbwIDotQHsQzGOKwekp6DhtFUW/msfXriIgUw
4CACxk+zie52zg0ytRmymR2tqVG1NbnamU//zudMmMuyviDT7WWsdLJj84JnIIlSnvzYmAoKVukx
VsbmYb7vSWxd7+XQE3LhHbyGiHoH8rae6FJoERtLagCNhNuGdgz5ttiCKBKpmpIYWAggBCMNfCQ+
5yP2OSF0QrBwvVmOkVYOSJpXDdUggSWCq7GWBqZ0gw3rc9LgiU67F+7JKm4iVkTeFjkBv64HXNP4
Qjg6braDpJuSsZMnTeJXyFhuHw0xhnSDp43fYiUVJ2so69s4e6MyQpbz4WLieMnAsgxiok5amkGB
Fq2QtQ54tLeOzz0KDzkspC0Z108nzbsxo7mSxiy0w3X2Q0eN5wjcsh70S584R6SPqQg+N2bNWSzG
lq5Pr1smfwj4mbxjOtTQFPtgBVtX4jw5YHPHpNBvllIhdsxQYLtS9pqwDAa3vFZN6Bm9gYE6Md5n
PhwfCARIP5p1iDh+loFpL5d/YTw00dorM0n5rd1fMNIWx+uwu9KiluHfF6GxLAbD0CJfHShdYzzw
yii3mafJU8VlcE7qt5GNkxssKK1mg1tQGA2pw7RA1+vhq6AcVQAElJYVtt+WRf/PRBl75gTEjOZv
ExdoPMrasb8fRHP60JJcVNsSvrNr2jsAW6JdkjGDne6DtXDeiuq3YBb6fBD+ZBenfPYb8nMIBIHa
DR4D4Gv9OZ7uSK7g6PD+ls2EXpLOpM3STTsB8fhbr4McZXxDnLJpuq+dDcc7Rl6QJWqeHSrhsB/r
RVtWsOEV9EcwvhEUw2t8kPQg9Xq4P8Mijlf4xszj8C5HU82yZS4vn2F5F+Gucz/mz5vO4yiwz8ow
beJrCb9mc+qTRTFSacTZkYq8VbAcCSYznEaBcEL1BjpYqGTqxVsvpslVyfr8jztOXUKWfnAjVStn
cCU4NuPR8cswDLsWNvs/Y28IdHyTrL373jyWtRUdkOxf+AlrGy8E3J/8cTI5hZo/JfcxoKkgbhyv
7esyxmq9lVZZUC54tNWCL9Jk7hG1ALhBCKSy7RsGBlxRw/+4dVD1hwnhniJ/cbj3tpDSDfL0CNM+
1dHCwBAIKYOmFyNKQfzc8eLSgJlxN77delL2ySWAgm46Vo5EDf7JJrCx9NjuxxzzCABmdUyLFvrl
vO5jecyu80Tq5UXK6GJ8QLlvi+Ncj2OhzPUkxUFjR8e461kZWFqa55PNS6p9yUwHynvPfUuHSjE/
D0sk+SQP3FRGkOq73/GIhnIWS8NZHlMQJnTMUhbtlhnkAKoO7Ev6Ukj8qA8G8J7baQVn0rA3LG9M
9FYDjIcWC45uVIbZvIBjjpAofZR7ghwJY4QuRd5avN6uAh9EF78KqtkQSLMqykSPzlq92FVCvNgO
mST/Vh40HMIA3pKWlna495FmG8mpXT/Oe6+xn55d/m+Ip+DGSM8cPZImPExKcMzMnSL3wVT+76Lb
50qaEqw5k2QNi0JplqChK2X1lChSPFfA9Nuc/k+Yovk9uMuFe6LXNFCQVlkZRGZ9+4435e6iLl7g
xejLpqMqO2AD7a5FxJnA0KstfivGUok/1OHOkJGECpM8oWDzGW57xhihpnnIabBsS3tdSgYwtd+U
vYrkrNMDnPAMM5gGjJcm3fYN1nPK6W0ji1v8FNeoaPKI0XJNjIwjUfWc8+JdLBHHj89obTPd80Jm
++guAezv1o9CDsJ9fmBZvH+8pBtQPiJf5lP/UyouaRnglOumH5XYL2C0YvoU3HWjPqZUZRab7xkx
3Yg/ddwfknQq9Bi29bLGVCqTsPIjzylP3nJFsuehlusQO3CEo1jmePN1ZQ6V8TcBruzUznteXiRv
vlEjshte1zdFlntJ0sG3jETcZMlFHR4frUV5bCn7xC01hkzeqOzMRZGYlHVHxkwNWLBmKJDJcFx1
WY3x5mGChBEC6f2qz/z5KRY+EtQc00RqZIsjzPwivXSHtV+zjYPksl2FkskU4HrfYAKfje818jBO
/7ydy7k0v+zQm1vpoYEmn3YL7j1PfXfHQqkMOtAm4McOXZGuIVmDk0xNTCl8xyVz5mNA52SqaMax
V2tC7Si6A18aorZDwJ8bblQ/HcJiT43K/VQHLMlMJZk49Kd/Y7XS6/fRBdyHwyTsRgaL7M4fGeqI
JMdEQW76U3RLQrwl6BIBBim6qbLZJxyynQNU+037SY36F2zWJmb68tOoyR/+T4j3FVD/kLb55oN+
/tNUjoBqzuanvWtP8jEv/dB0KH+0upZF3GTZvoUkMaSVYsipzPI6M3IjZSJV2bwEXAHDqRyUjL7x
+3zN1JLoQrV/FBWj8oJMMu8WG8Lb/EPhzjJh7BnnB06H7O7KPvuCEcRIZw4aHwcYPRzT+q9Slk5G
5GKgIM7/i0PU6hR3TCGNo+1fkNdgV5N8A8tnBv2askrMuEEXtcSczfOAdULZ2wqDtOrbyKFuQowT
gAxYD236IENR/UYRorbhAkpg3aoZTHFi8PCtg+lfdXyILKJLMzKyKy9PcPl/Fxlj/RQ8nlAQ5ZVU
KI+EFmD+Lg8/Iu4nLimZOBLxVHWHG1L4DjqaPVDH1WhpwyQoIviq7iWYY8KNsDQyN2EO5vFFZBwz
jjEB1WPk93B25z+heONGQ07ZWUwUrSf7OV8HP9x8HLXo//7jBQmSzcYg5e2Ol5nP69sl5ZUcqQJP
Tf7wC8SWYKljqJUZF2gMQdAH1DZOMtJ+JSQj9EE+p7S9M5h/fSsidwRQCuXglH94kRhSDF+/FGNQ
+Ow2XEMpv925zFW7zE48lRpI5Nto/o1lVKRc6MBYIaXYwvaXcSIxfIR+Fd3ia06F8j9YI+97bThE
cT9GEDFCieH8MamagHfPk6F6m3qbf/QHZuS66goK6doMavCkovMDKydXW9PJBn5+WhO64T5cAa/q
RAsFJokC+gGe4m/PGh0+HrOjJNGy68jt1B5gevPl+k/YxY1fLBhu5UBYKiV61oRK4cU1JjfLbyTS
hvIizCaXGB1k9JRvuFsDs+DYIlpCeMGUiS0ZC5uoiMJbYRpQ9kpOotN82Pyx7Ni/0DnHUV5wjwnh
tF5MtZ+1ARKabQLllZPhAMhbrqEhdihys+Q9Mo4QWcqd1Hi2xVV+M+e1pOpLRfz4+TnpWiS1bhSW
PT9/4Fegx+AOLBXx05OezG1x1m3eMQ4MP827Dn2+l4ToPwIBvls+AmqPi3JJ8QVFDFiVtl2qEFpE
pibpKYT3tTdWKVzajc8i8QVYRTXr3iVCXMlZTm+sR8lSgZDuYvVA7iSzJL5lVZPEZ86qfp4lXBWc
ZcqiorV/cioRSnibYtBAm+eRdP3u5Te4M3s7CFjwAl20xV2l3BjAZvQOqwGWJGFYmoauBmfDjVKp
YjzT6YhwdzpLKp43acgsjZGg3KPlX6pX2cMHlRT5jWfFYdVKt46a71W+dhFkyl2XLsV5w8YrnfgY
chTjBWQ3u+hWSj/yAafJwA1Lnj+JYkI3Ub1hrvgkRIzCXKKfRrsSR47gdDD0pN7OiD/vhlhdYdeO
0r31R4+eXtLDvWaEfbxz8MwTNUr5qNlAdMArw8IuY/HoM57KXJdUXXjzCeWZrn+0F2z6v8wQQL/Q
oVEu1BsEVeMSzSlcE/QUWDQoawPhdLs/n+xcFScmAn41U5s0JS2UQKDw5XjNexdRZt5z8VzI3q2v
9oCSJKQD2a8LzoHRPuCbBFKTlVCzAYEwmPeXtqwG2zBoRnnJ3tP/EHjZWERl3JITCrHPvagpoAag
1Zm6oXfRTPnpZvTR0cJ3A+pnn78kbWA5QxCxDE9Ns56ShZUrYne/8WOHg3eDUV8Yv56ioBFrrTPf
lJFowB6mbrGu+NWymGhsfcNDubv+NcowPgx/mH4oxOBmZ3S0/X2Qvqaej1t8HPF0YurB+QIHO8uu
lxmIPCMmZKGdVSlvhwulvLrPEpohm1yWejaCzI5AiaVBsUg1jLBAdql1d8rahRtaMWuSgCpdcO4m
WuAO2LhtgBXqk6JHqzwJQunSvB+aNvoE7AxX/zLYaVMlgnlsjmx8r0UcfzNE8CLKCfROk67w0uvD
0M+9FHWfL4WZdCcQUEBK8f4Hzs9r9BLorLjnxF1H4cAQqdDk9Ds+B35GVP0x1DFjCpibDPObvZTp
KSkfTP/M2MYa4a2BYUHp81zerTVAvgOyj79eUXWvmnLLef/cVvuWSyNoqFOMr0GyvQlkdX1lmnm7
KzA5MDxLBMQjh/M/942rIkcokkRGlTSPm44rIiFmfnBolkDWXYm8dUKTOwZx89YodAtqlMyVZIPj
CFuhju3sFEebOyyxRqVbPrDLCnfnZ0O8Grgh8tSX/wWZwYHrWLCeZJnP5pqGGlffqmG+/e47t8xb
z9qDHbyoMOh2MBoC5tvMrxe+KxX0mpv8BYY1gPVm3sMKlQC1w2Sep8zu43pwzHG4x9RT2vC/ySy4
CSQj7pgFqd7U+Y0IqWIKEBb8UocmETuHIZfFCBD0/V+Ws4H+y9D7Z80FtLwEWZ9Cm6TWFIpdNKnx
8h+7TPQbExnIY17Q4zF/aNrkbODX1p40CQqn/stg5WNmDYIOVHdeSHA8XUe+dPeIsZiV59yU/Bfw
MzCNz58woXRKP3dnXDXsDqGy/IwWaTi81FjX3DMyZmBiBWizmgHJIzdiCRyd/XP0G5J7I32tME+r
hqTgqfhHydktzb8h7ZlPwG7Ja2UVdYYslclPlUeuphq6zmJeTD76JdG9bB/x3Cwl59yX1bd/qDXt
IGWUti4k0qTDMD2ofCulVMf8nN6WfhR/hF8GJkuQz2kw4up61IYKaTef5dGaJlIAuVbc/WPMZvBH
3SNNygP9mWzmYJs3u2JL0eO/DSfHvPpnNHccqGdAyGpG6/4JxSov+p90IuRGUK8B1HLbPE11bsOg
t7upNTlYeVxmPj2eECSOv2/GRbyVnckBPOzcjo+M3AAPwdTduqcjnSX0JeG7spEdWYwAuyrzRCie
YT6CqQAUxjvMuAVjSgA2HkgL+F0EeKs+upHa//MaqI0x/HT+4qERT1iALH+H76Y8ao6nTfIbGalJ
9CQq1Yt9LsGQ1uwF/UM+ZfS1p/h6BwRo8/TU4nXdn5OU3kNcSqzJ6BQuHnEyMLMiV+vIA2376zXN
1Ev51q/9/AgeyD5k+rwHGRm/sleeJ5TIj2Fv0p1/BNq6vd6VX60OA/9ci3WbVCND1yUtDrQQkEHT
Gh/PjA2aRk30A0009NdeI8pEQ7BQAfFHbULvXKcJC2sBQLpM1o9LAsEPzVmOKnmcSd66ezj5I0AE
cIbkYFXFzdIiuyNPOToDJb5Smjf3/uzde0YnRY7mq16wkEtENnwX09pWSv4YNlC/DBeyIkSLPmiY
lU8Yj0LNdjld6cjrAtbXAwfUsHfFc6Mu5Pa0J0tF6yUvlq9XOQYxJqwlP+1LRUGpsAEHeo4WIEqD
SFldUW7e2JRgMbWcZMuR/vFAF0BehYwrVKjQIiP1qBygRQDnKBo/rGjH8BgyfGydxVt4Ba36dTt0
qgqbii2fZH55BRJ2/orasNcE8SOlGWORxzT+HNvQla7bd8bJUNXKuiRl5TV0bC02ux6pQGhZD1f1
v4NWXEQZFAP3gYvuzpgyjxMAmUyLaHW5RuQNIJLLHozkI+gCYyo+aBiQIu/96hf1iJVEeWLWmI9w
BDsipko6Mhbx5lcyjPiXRbbWMFN+qP3XKCn9fj0f0L34pKepWrznkKKDaaQNeoc3m/fxGHkC/vJv
2KqiR/EXJU69BMCqCpK1pM4Jf+F4GLXtqBTXFfWOjgeBw0YQNe4Y7UZEbs5sCpyR+gVIwk7QXL2i
M37Hnh8/4Y5mNOEWN7XsidZjcxTlcrreaYxOsfaH8+ib+RZk2+U+unwWVxWqtg2ptwwRaEtVkras
r2Cgwx6IKYVGbqsW/T8tl6bk6OzObdEeWLarK5OCgLClDICK24nmWt2qObV+UmH0cRbJl4Rs971F
wp7aOvdms2ZlinGoVrAV7hhfWc0fhL/1EMDAeILwhqE1WbJx4YkbGVmNlqvvKOlKgnhRU/urkpYO
5gEZsP0mgD2UsGjn2cJYoW/CZkzRIi8mDU4cG0byKCAhQmkzDeziES45BvCQYO3AD/LacOff6gkX
8ZFcRfebkJLx6Q5Mp4vMPPtExqOqnEMUCji/1RP/TTApHvnJTiWVT4Uq42qnj7c4ccEs8Ne+yFJg
HjKD1bjJjzGVqqCii7lsVTDzew03W52nETOHz0XoiJ6Hc66GiHlLByOgxUx4xMwr2zl3Pf6kSwPm
k2gqbbltDZYdl54ntMPNcfy+riJhaWovYQMl69VibQXnwYo2/IPh3beZJsUg8xYIA2QwsW0VhRBV
5yiu4IuEr1iLXZzl3hpA+WPwVh75nl4/EDUOFuQGkPkB2jyBlkVavsTaTRD2Hs4o5Tm+LDtHTLvW
PcaIhayEW0u7vJ9ZN5UjDnlNNXR7gp96kWwsoVdzxJS3deusqRX5MArDeYVv5urGy8T0vYhVpA32
XCUP5jcan39obA8Pgie8/BVeMzkzcsrKa7INEBpdumraJ2ceVX88Mhe+ezkQA47urnvbOg+6dz4u
ZbWjUC78ogtquZ9TKq5G9tVQ6dQ0bDMcicNvCDpc01R8MSCozRWb6B9HEcaXkw/wtL5M+wUOS9n3
mGS5iifhg9dG7zB9oq6xdVy/7gaDQuLXVXE4pH9oIbMKF7YfrCq3OnRRywnFoIEXX535lk+oIE4z
G6utzstfB4YtRi1BMoBjpyU/vc027J7dNeHkok6i07QrPwUuI3mp1VXBVe9UWhrUYGha5jxTvlAJ
kIkZpUemCcmput2Y81IEDsFXH8w0jpNU8JqOAOnIHy+rGfOeeIbLAQsE98oje1rIZzqZEen2+MGW
W6HrQcJjaWVOEC+rXpXVXgW7CCLC9fpmA0ClO4rs+H3QaBjoeck0NgmiR0MxW91bHhzDcAAhnCSG
wK1G/c6O2zKYA2zZ1edVoFMP40UPUeAP61Et55smNck0ar2biFPvOH1GdBsPzY0mjxsSioHW4gNZ
PR3ZH5dMpl2yLa1NuRiKAREHcDRbrs21u0zIclrEbSY78cCPxlpWvseB2yEoM4NSKdSpBLKUYmWg
+hEEM7TML6ptFxaSk3lxgCkpWQX3ArbhwF2Q46lnSn9N3zElJkRtYX+OP00vT7OWLIbqWP/x1rAB
dXzOSdtQIYczTVHbG8KpYYjBDnpoUm29fOVYNiPK+uUmF+i/SfPXvZPp48qjC9z4ZAvPxip/5fJA
eGox/UDnbm45mH8iGzBuMp6acLVC2OOHUck8D8K96iUdFWztA2RTikxxpAAgzalerJTJb+RZtW82
xMvQZIFLbZqq0oebpj1obijkFWHxDqdrrfjax546AduDdhBMD6WkgxDedOxPDQBaI3puQGJsKW48
wK9oLQSzk+Kj2JrGZ9jKlhGy3vnDKFmm+xu3cdwlqkperaBVYhWcbJffV81c5XXC1A1AmYfIMXH3
BPqE+zWJ4YtZ6II1gZp+QwkK3ZVWuJUuizlORMHP5cuvnq7nW6uniWN0DYApRQeI8ug6QRi0mXnV
8CSKU8/xlJWKavlFB+92MXdBuSEQgL1sXD//+iv+4TQnRMt31P1Y8JqSi6uMWChEg3mVsfFtK/4G
AV2WUPs7LuSIrek5f9iTnZl5a47DX9Q3vn6r4mpw0UQHHWtYGkeTo8Or6r4I0bWeNwtpQRcvfVay
Fx5bg4KdcN1gY7Ov4mlGFrAN3uVGce7kHtF3sPkqInpQEPIdLRvfKYCHlfPZgfA4Ja4ZZMq+ZPB8
TSLgdR9XQzkBIQyBHkBbtFrOJMMxxLdI/ppwErfIoYrO9HrLIXBJqzH/57gwqPRNxhoPk4odx7h+
UITpOP7b3Z+sjsdstNxkM6Neff/VOFtJIwQOj096HjV5Bh4CfFMSsN3eK+ZPAfY0d/ca0/mnqorb
wytVtvM689tV4/3ejA61BSncOPkwSPWYnj+QayFC+5lPvjmqGUUWtv1etNFQ8Ju2FiNuUGmr3FuN
k4QfZfHgtZT1cIv+Mwm0quOfFVG6jkV7USIEMziLEwP9JFCYmYxcXSD178ll5LpAjK50O5M82HF/
sOYYmtt0TFSIcL2bpK+3/LDg32PfOvFfHkSn8scnl5YP99ZVVLbK0AFTNeqoD9AXPrS3hgqdLAzv
7nFFvSWHYQPyv11Tn+yp/vRTGkP3aAkEy5Hyez5d9RugptTfmbXLT3yTYbI04DufumTy6oZ7n6Bx
Pt9Z6haUl0q3vI5xaZLX6FYWgF4pPt/xYXC8sHH3uP9Fp+MsF/zcXIZr7yDTuDCODamEqgsdlLmr
4BnUaM4cOoC32xvPC4E6AjBaj/1KgDtA8MR5lB9P+YcZmlmxp0+7EH32GiHJKYE4wOSArhnS+TRk
yuz40HhDyp+mOK9/QBlJ8s/7ixt3hS6Ds14ySP+zVu/aLU0SD62b/SSOB7qig96HEpBLVNwMARYu
tOUBrOT7Cfk0Cw21aVpecQZ5uEyBUg4hPFzXqg+qlHn+1u0GQ5aesliQi+UdwcxNYPeyneMpjwW0
B98irnGEXMXNXPjsG2kXn6RfrTzXYQkgnN1etRx/Zpz2FFO6bIuzeljX5WhifaYiW6kJQrJvAgQW
hxj+lUCDh/svSkeo15srEkihRdLvUjj5g95rW4yKgBJmJ+CUdHOv+Dm1Q1JzHxGazya6ntWCVXF5
UXrr+NPUi+gtt8xtgXwKmppiF8Tv6sg7+mO9lvhorMtl+mlDKS+N7KrI/G7LtG8xl1yypuJOp4VS
Aq191YSsgVybJoZ3AogyVDoNFP152cLqb0z10arGO7060w3vIU1kMm2MUTXBM5PIjqmx1WCOU4h0
DBVOtGMkaUxdK05W9Kouxp8LKnQ5SIuA/7j3XdOOTQjKJli3PRwd4Ac5czHNkZ1zwaX6BYmrWpJy
o/2e6wfW1d3l8UkTQQTgSLh6CWuaWa2Hpc+erZuG3U6y8XQoCYZjiAoUxWNyNHtNw+BhELYmAEEH
Fwx1BP8r4Z3Q7ZMnyXCul5IMxJwoWpgBzejzBC8Mq2lEL7pLSWm61NnY9It2jfVK/4zaLyswpDyM
WHrEFKJ0s6V428WBRPaayyc+Xui5GD7A/xcM3paAQJTfPCdSAoeOXNm2DoutXr1DvVMsszM301Hg
lhZCF69jnlCK5vAcVG7hnlfrTKkvtWIHhcV7uTMukVzHFFaJ7zFE+/xU5976f9rLxs0bRCN6FRmU
JEUfjqSAyalF03j5Q03562TAHnbdMs4WuMpYusu2yVuyaECovj55sd+Gss/HqH2hd0jCw++KtYSL
gnOfIi1Ntx1L9bLVhw0QJka5EVSf3ts0DbnFv9jjgFemnhnwNqVPzYnkD0ORBBoBCzMKlJ/y4mHR
SWCzhz3FYMw5OzpLmvXBRN52MPPSFGYhTYIsbWskWQmdsp4RjA7B0Tr539nXYVra9WL7RDcTH9Fi
Trc1rUaew+b3n/fV/uRZPBSDrrPiWuooEJ8Yqha9PV2gv8C2ubRDGXu9P/qmGetkMh3JFTq6oj8L
8IMCcabGLNphfSjdSf8fSmqK8QxyBss8ELQKxoBOtvUsr1399BZFnzOeRM+WSNLirxrpFdiqHGBs
cd5WJbLwsZss5wg+qHX7SHHznW0NgME+8d9ZyKgwQfXhVAUoGlFmj3Le4eSq31KCqmpziUqyaqy5
FWB2nuL/lObbXpezixhM9Qf1eNtMvptZdcY54QK7n4FMAQqTzdr1JH0LODAKlB2/qBtepFIek3A7
wgDzpL560YiZE/AHju097m2qioxjEMT9qw8z34dcNuGoqMSvZt1m0hHWskccm4Y3uQkHKu/3rOUH
3o9NIrH4mm7CEQdJNCx6OpZoIInErITDQ5M/KO3+p6mWnuei1akujosqz1T5Q4dD+GI8AaqXomQW
oBrzF/VYcMEulT2hkQHSNcghhFa0yBbF7bCfs9DvSxt/Obz8jTYlPmY/MS/Rn5zObGHuqWc+br7W
osyBWVznqAJt6XpnXZVnuO23apq8VIAWQtnEBtnuP+BJktrZv+r5Op6siXaioJD/mO2MU9TREW05
iE8s6mZr11LvilmS+n/mkeU2MQv+bSJWYQmhju7FAyfgBWU1VIAgMCmlRVitV2JijTQkIzy04zvF
KoOIzfL4pnN2awpCGXcFUFy7bWCD+LYyn2QAU7mkHiV3YAiT8LoeAi3n8ZB5FqJkzTyoU1iqxzJM
5rmYeYc4bpo0TjIid9zvTioOMq10wTm13tSDU/4ez2OSfMuM+ZZe+REaNtIKKm28+Fc3QvpEpNeq
CZLvaBHmNT0Cx7KXbNQJEjt0RRsHUE4M7oZDbUKBiECLZnSqjEK7tSATeqYMohXZt465f7vsGmUD
6xObEff09QudawuFGX+LcksLKDHDydcyVawUrl8sgXxtGIAsLmjqS8jyEVpFvzB4x5R+ZUY7oCn0
5VSm4f4YDdy309KvB8GlukX/kfA4K7bRQqR81UmtyHo0CW2EhcKgtBVe48ou5IJpp0vpD+QvKo/U
y6nuvJu3Ozmndx15wj4cgO6kc5NPgTM9jdjr8/cIiPqiADN9jYtqdw8r2FTzPmTHslODVRRteiUP
8BtJyKvEd6/9WLBSBEis1MXVUMQ2BdSLRjciAMyN2mpFZnp61Fz4KoqHzc4cwHRYIsMTEgNergA6
ax78by4FryQzUIExNHnrvXhqOYhG8lJP2KabrlTSAeDI9h5yCm2DviHt7CnpX/Jb+kS3wlTOcX9w
++7tAsZKTPMqPKA5qVzrVVpDtQIH4i0SG+HQbJqmGSwg4cndkaT0xTGpmMRsKbj7doX5i03H1j+l
wmT/ysBTuPQ77L7c+RU38JEc0wkWOTgyYoOoO3d6sdboyyhquhC6c1G45g/+R3c8zzbQ6FkP+QBz
F6BH8MvjIxjbVL1axzmjiCgc4BfEgrQJS0dLpiL5v1tEUFnHQv6SwEEXy/LNM+wVzOA9BpJLOUUP
6njOIGx9tA1r67pWvGPoGZ7XzSTCSHXbVEr/ysIaXpchksEy7uNhJuEBUcGi/dnnXLPZRqaJ8Fa3
Vh/akLwtGGCxHTpx6xTp1NIRbFYXQysscaKR5bvUk4lpgMXAUg+M1TPqaf3+b611WSFZwQ6dzePv
pRBFgpyzQGlyLqYHbOZEctD4m0T0MRkGH39H/Wy1Nuhg49ugcznQ/uuq7HqcDHz7ZW1mFK6QeWMr
4WI/lSOnTk0Ai4oa7DPWrL6v+52JFWiXykURIweAdouOPvKiz13A+vkoNIvA1G/JgDOkKH8ilOd+
BwobGHt+BWmHxStCXd8hAGu7P5u5IUOMz6u98od5f+Qbn5oJ5iiJT0uWJOiZA9616GEpb/AOYj52
Xlbh8r6JOCpqnJLPeF7oED+pCJDj6tsWRO+A5Mijo6n4tqnswm4bMokR4A/wAcbi0gPiRJWskjcC
TQj7JAlGB7IJStA7ejyEfKkkyS3e6aeNazXPGv/38msQYlFMywgkLiCviXpH1cJRi2mfhPfliHWM
CE31QrUKgGiAXl9UrIVnCA3K/FIwYP7EzBEqbG8CAnOVT4tof3pEEAIf/vPjkI5rWsT6hcb/bD6i
ogmlZa8oDlGBSoXxQXTspsZwvpvq2YYzyvbKsSluasM7dR8nqk8Pho0zqECDbAcZvU4aEA2Y2GyL
jufp16HD6IxvvBaQwv1ywJRLw0NpqYXLCL8vILb9R9xyL10ZMnzTg2Gy7sIEc+Nez9j0OeP/HJza
skN2avpCiUB4KpyEs4k7d/WOIXV4p5klBbOjTUCMCqPZk4N/YXfVsVLAj+sW5D6e/BFuRUFwgAsY
PajKLw3ALVATyUTDPTrK+du+OCVSv2XHokkS5kWWirfaVZFsZiurcQjx6ZuneSpzP1G+CsyqzClo
ZqvIZ7l80RXriXFCQqjXrPNU9B28i8OW9P2AY6XFgLK3Qy9VHSxSd1baOtK1S1/FxvJs9bNFJ3yc
ZnJrpDVgBTXOL9s0miXCZwa10X9ZHIne63XH0H5YJqCqX5881B4ZlEBeuBY1MExB15EZRJUlRkA9
3HCZZX8PjLsul1g/j0Yo1ddlCHU4oJ6WiRuwDrIInncly/8Qt5mjCVKKTHDdcagReI9Htyc249Gf
gYyZRBIegecaBFrJVIhwkJi/v4HhRFK9znvTeLmuL5nIDLWR0G8gMAyuBmsCsz5U5KrLfU341Xle
Wb7c9UMAVCQq4ZhS0cRg/wQDq0wE2PBVdfaJje1smtaI8krUnXEwOBkaJhTscrA/ZWo6hV5irzHS
3T7Xluzdgj8rBRW3LJksMOmvk9jLwCK7bK8IInHf/8F3kKiLEQA/Qtswrax+j6LGh6W+hMOBhlUO
O/JlSw6apoaGz1KyQ1TpWELv8zcUCX/FZ6wT/nHwc0mXfKRXilT8Xw0jP/1K1p5/k/dQ6Xx1Wqsk
hJam4euY3DAFSylsXQXzB8qn1bhaFaUAZivRYLXT7hyIJH1w5ZcafHhCz7xhljbL7u38wCJhntfO
gkrQGLx1ZUu5WRj9YjkW0kcQIhmdPMg1N4Tab6PYoS4UYIKGAJsqo9w9z/FZXwHcSHaBIkwvDhS3
fBIHoNLAyUTpvurN4f3NP4tyqEiikvt5sWVElVRMhkE8nbaLoCnv71hNJhZQ2VcO7/J/1H8BE7yg
XUbkXVtX9cHjlcLiL+1Unjd9cdFDFIxicINuhglwqmhVJSSB2MVBh6SiLpcajagmEjXYVuGd3td4
xObTZiptA66TJxs4iWA8xtMSvDz5lFHNXfTq0Yf79koPogQTcpC/7rNYZU89R9/P6KDv0VLVHr7Q
nQnXXQ6JpGaqgAXX3OTd9d4YJel04APezBgGFjKzAjw+wiioKJy2G/UAoV7t+b3dOyvVuKiM7eg6
VhFnLIJCreEidFkkjqCtxBppqj/I7T/PpLCmkSwdC6YXTmEPMbZtBZwIqLxVG0721RCT1IvfOtvx
hOkluvx5hlB7uWCAAZVKgDTHMcWFGYBuOY2+84Dh3XIgr95H5wl4BPmGFVMl7Tq+01uGRdvrP6SP
9QmCcIXmdAn9SdaCRFiSNNqgATSLcKhmD6+1gyKYzU9QZzwjjD4YvfFORCo9Jk5uFdiBiEuiML8N
isCNY8hoypypow9rqtem64fS1nfN0apUB6xCBLK6NaK9RySZhL/QwWaFHxL6BZoiBxzdUixrAD19
c4zQGQ22bOjOtAmbwa8E07EZFujAzK0v97p2DpbbFC9Hnbvrk2bgRrZv6wkipsp+1I3ByeJJS5lR
LDNSgxE2LFnkYyzv0poq4zgowwxi36imbNa6J4wFoDKRO99WsUOeEh81BRCfgyzQvI9kNMIzzQ1s
gl+1DRYUPYoXDqTcno/vImRGcdQk+CgetCjQyXkFHZztnH6H8zZbSfn1WjMfPtj+7Ho2+9qdwbiR
bJfS6QjJkvZcmVReYrigCLnqTZzpzs53dJro4pw1EGv7VlB5JqhjIk+a0FogTRGP+EHz82aS18cW
nxV6kxCiHrnfF7CVoE91OC2tiGz/MR1Oed6As6ZfrHF7M76mg9ezbpKhTpgPX60Jx/j7vbQMHQtR
3KItOimE2sh5nwOS0diI59XGzY0DRWxebWOLS/n/dDiTrgvNB6859+f5BNH1WcT09tdboxh1AgY1
gE66kLsANRyA0bRVs4j2xzOO/ED8Q/BWRjsvFFmXeaQ9+zVDYRyEiFYh21jIPPEvWQYmIex4RxPq
I9ZXf0bx10pH75J+UTv3U+hDVdI0ztvt7uc23OJzgZ618P/HV35TgdY4Ml3UiIAc3C0+DgBcGkIO
TFQ0dmEFhYTdN9UCx8wNBU89BV7WWqrxg3E97tvfX93ILbgkhpjzgegJ2vUtIXIIPJ5emO45FA3q
3tUGrWiaXi4B0NGbTsvQxIjDXv6Wp8asObjtUGeHA4Gb8nSR4xUi/BiA4Yimtimwqac4A5jb1BKY
HMb9xht/GFYnZoyyw6eWCgv+sHqM2tmqSDU3Etv0hFvpLUdSTh3EGTquEJnLlFhVxMV0vjpccHVX
NHJmVBEoheZqpFNshecLn30SX6HR+aVRq/G1kF9eJVWPK99/UB4lePmg7GBfzuXwnPKAVntoUjDi
iR4C/QcLEXEK539dEdmG2r4kYcjOnSCNfEZfvlzRcPh0i/iK4H7Ftq9srJ6p4lbf58r8ow1jZttG
TIQSiR0nLc2PTCbMVNCMdELvX1MU5WMG9DYTY8vqdBWyzw+fZ9YL9/hJx4OnzYpGZek1Q0JhauAt
+x/UPPl+bL2BBd8r0jm3ZlN9oDACwWeLIENEUFWbG8kQiAalFTQzt/vgToIzHqbdLW1ZGKhz335X
hRVW9WESg6UgQUz0hvjRaPcWzd3GRjmPs5M31CLPzYEqLvNF3EWA5rQ5PqqUGawCd2jbgJ2z6jsD
3XyarruPjmTzSzf/kmJw8CdQ+/hypFqmrVndHDrooDHudEoRIvV2BHKIJylMmvurCZ2v9DJtOEh8
DMvKuNPOtqz9E9dOk+8PYhsh3EQtnT3rxis9JjEIUOX1xP4k3XAtGnV7o+Ga0V7i0W97nr/wPigQ
uc4Rtju0FvRYsii2YaW2L62Jrg3YHfY6LdYHsC7QzK8nNQyoubfkKciGVfLCJcvrZR6kZPGjUNdE
agOPuvFRBoMutQxV+fv4IUQXSagvvpbRoeKrkk74jHhcje5jJdWIR7Wpq0j9WewyRs734467Y0/0
OIdaCuDkn9m0xQJEklZJU/TZXuxpWeFpcm4QMFrIhPaJLd4iJNQzxiO8nXG+tg5lFoxKZ8cxUbvy
sjSc+2tS9vCuOFdUUaJGlVMYk7z79o7PGMdvUZ1H2Ywk5ym4rPg5ttym83sOQ5XDfPOZpLc7XZrE
dR5s/STohHiUhTgVTy8KGBehzjhWFe9zrK3PT6/aMFNY1Lr/68I2lOO3de3w/CtDHuoWqaJmolxH
LOERoCTno8zGukfi6J9rM7D5ljDEwOrW/brZ4vgg9GVbdXTEFn1CU4RCwdV22qATjfiChQg9nloG
quxRQi0RzGCWS1MRDy5tzGg12z58Kh7v4YJiM1/aLcs5sQEY0v0hZorL/WStB2xYof7STGw+Y7Xh
so5a4kg6bzIbXMQLl1IOa0TWzQzGXYzPxFZpsGXPY5W74j5GABm2AkilKreLHl7R68JJWJj+PF4S
fEWF8DI3+Ve6kpBjAitqvlq/puobMwsSKAvnYNylOTKHOWBWxWTBXMGd+RuLZEM9a2JSthohX3ai
O6D4Mg0q3AfifmhGJvWybsjROtvhwrwWCVJY+hoLBauMfql9ODFlTZSQDo2JCbD5t1hutNhPCgqV
zHtt78XJk6SJYVphCURWrQvWhPe61ixQ34F42XKaRPzgvM2ENXbdLe7goW4uoxG/vPDntAzG0ZmV
py2braX/QU2NTwRJDwHqCc4jn9KXGCiTZWk+gEwURHVNgaD5edWeO69l25ERTH5bxMhbCw0++BlO
2UxPWb2K2E57+yf44DGSjOa9xWioajWxnND9KFrN8pLZqhHZjVHK7rwr2gWt99qoU8rg9mFZrWUf
XTd9id6RnVxR5lltS12Y2zsTNPIeSdFSUUALDiaVKFXUCB104WGrtbpxe1dVO0QLv09u+J32be8O
QKoxa4QDDkCGeWG9u7mjO1u0IvK4Dpv9paIlQSPofGvqF+7JYpzKGBtXBovTy/U0N+GndJgF6nfZ
k+vh46I4eZJqM9W9GsdPU8jmAZ+sJ5pNsC74xaUgGR4nNxvaQLw8lB0rhBrQy/3HSW7Ia64OmIJw
jpn7jGef1kHufX4AuYCWWh2KtXuugrn7hSC2jnuJBMaZcDMB/6tP8e24Tez292Q0d+96p1uvgt/r
SrTrXuisS4WKhMERHR3F4yiHNpiEaqsgac37+Txd3II/DoIEcM2fqpcGZuNfpTAIxvQNRyL0dmi8
iKOZ59MMoNdYGpRKWBbsxsKuuabtRUmzGHT5ErbCRFc10NntcwXZkmnNCfT8btGS6WaZ5q5GVUou
d2oPWYvR9IPMYhCH/7alqnj4pkI/QpqIj9l3HeH/DAWuk83zEl+7uOFfDbEFi50m/gRlyoLd/VTL
npzqjAuXozzOTLkq9yq//5Kv8gZj7gCgV0MnYVT7Y2R8nr0Idjr7tKbYQas4LoQOV2ut/3XTUWW3
O/EP2I5/XIXFAs7kQUIXAsFf7Uao+sxGtA+yS8KH/uQc9LQg2qw5YTZOxkw8HiTEt4Xy7sfjN0Lm
k5AZZ51UvLceW0GuH5C8/dYHhCuW7+0+eiYAAzk4CaRxnIep2pW1rbBXgBiteN2DjpdNr6/NeLaV
JupsEsSlJTXi0+8DjtJKJ8f2IOcEsFj3PP3YAyzCWAmRXGZqhqARjDkZnzhbLY+ELo7e9U7IYBnv
00/QJyhu4yZ9k0ADTUTT50NIprPh/UT3xR0RVG6cIlj1QAv0AKzWNFN2jNN9fW5ux6ibq7ItAuxW
p9PWGj7mbtz5MKL1ksH6f3aZSjlR8SSDq1HPV8ROFFNHhwAtWswi/GJaj9m/aC4JgMnHsKdf10ei
NzHfsx1jp+n15Vz6H6Nts7NFcgSj8xb9FjtGO0Ml/QoC7iNeqwEUc3Y4f/5vutb5CQAfIvb4Gaww
oOfExXlKEQQ8NWYl9edJNcvKcKX3SlG+8ghlvSNYmJjrfdVGK/8TX4htKowwzrafE7HDjiLoZVFw
weKSCe+j/s8QHBx31Ssxu3j//QfP35dPJpIahYg1rnMHAiVmCZr85FaMmUV7pJYT/WNqhY62QsHV
qQM2kAxEMtRIjbs3laj7GcbffTUSldURDzxMnbppJROy1xdlgWnFmZSt5e2ZDlJfTGm/8acBX2aL
Iri/0h81WpXC/l13XnbFFwFpRz/9zdwzsmLhzyqXakQf/aF6g6XDfMpQKr+wnvcdGl1W2Q4bH7hD
0aJKMPtbyk5JLqhZNbXZfuo8wmAQXjWVPM/0Tryho3jdwHcT5T9R9UFN6Ao8QF2A3ZlS2dhcEvuE
UPwlgqAUnUWreqPZ56chsdKBvmED02nMc30qsveBDkHdTJS85EHKuhfjK0E5GW7scX3qDR6kbD4F
MIX8VqwxRRuwM6pry5hrjokAQ83dpLgL9JTn73Ni7Pvbr75gwcnldZI7yRRewpeJ7dnSn8H9s1dU
zqbDCnRV+Sj69kAvRb/U5juJCuzQk6BIs5/EQEeVIP3XQ0dW4ClXfi2G42frnssB0y0M314+npxs
Pwsd9f38rDRuAHYcQlUQTEAZjIsGxtr+7w1a78I0gW0tcLR7z9LgsbE8DbkIMZFLQmvs9vV5uOSY
95z60J0oJljndIGOn+oKo7dKyXdwh9JYVzA2wtY519w742ukRI6aI1OaIT/2ezoa/kS6agIfDV6G
psuPyNKtBvjI81JrL46N6yzCKckflZYTjQiLosRrFMpnZvE9DA5NphEiknOlCJBiEDerI5J3eAN9
UusBGYTDnPFWYDOFqJ2+AylHKernb+lmqRGvymqMgsUIgc5Cdf2GeQtTsvZJ3DMh98jHhciyYTCd
s7Zu9w+Rirp2ZDpJSRcTgHyoFo058oyD8xc7jAE5ShZMvF1bNdHpvIAVWnTC5WLx52i9Lj9fk4mm
rfQ9Fc40DpVAPYhOmQCqNneoLZReSJQo34urKGnoHawwzVSC1zQLQSYsMyN2/2DkgUG7feJXBVm9
oWsDxNkEi+VZ2swOhpwTcjJD5XiIHWxr+eTBzvrVIym9be6hQFM0GrK7Whi5r2mwRj099u6p7YQt
fC/el0d0GeXB7ycIXv26utBltSbSO8qO3deoUt8wg/G7Y4Lu6OYw/3ckDv19jw2lJaLpSuxT4klb
isumt1/MdAvMg9EInak33vuTywpL4mti/a66ISSZR4skU2eXMPIgsPzFBuLAwIMsBFq51eyQnc/n
7e3kWuDVs2YuFydpzl/xnfDJ9XT0moBTISWaYKLkGTWExMJa0mit2UUzB7Cc7fsDGPc7HYy4zrkr
99ftyj4pKrcX3t/AgHgTmGvUsT+iv0ZwRGcWWp00IjPcByybQ9ynZZxwYDr5PHxHfPUhPM+3MRYF
vk9COeoonO5UqQ68sjK2ZfBc4lzREXbeGY5ezfIq9KB/apNgmEdVdNFAHQaRKWWraxsxwQljeBS4
xz/vnh7EUYQUgjFUX7HpPecFFvtsN/7B8kod0T/JnDZaLs2hH75Woed00XEHUMauk6sAn8j69hwV
ROAmc+OUz5DIKHMY7nU+5NJAlNVSpEeydBLBvwWJQuluHaV6q0Y82MifaE4ifrFvgmbDXb9LryAs
qSJpbxzrRXGrAlvKjeM5P2dUdhnzDWG+s+0CIO2Q/QS0BgBTboaHKtIbxgkZ4C9+eJK9V6e9FCYO
vxWaqwPyQvnrT2xtWX34wY0xx/4QYv776uRqF1Dkco1NDRMRAu1KHmO0DphU7hN8C2JSr82qLzGr
wxBcYJmWd5mvQmjK1X6CK0kDgbWpe3+1rPowWnmmyry1BKzFGEjO0CSX3yP/lH7skzQEt7fm26kA
5YMDCLK1IUlszCFtsLBAEHHg7uukgIdBNW/hApAcMrsG4L1I/1A6iFK9Lg/v3XJjZf6N8tT8yexl
RYc0INj1xNzKa7/YcSQszl277UiJlUJ+hJDh0xjoM7IK5C5hCLcHnfWWup2+LqTJ6vdnqXZ6wsGs
lH31XrCn8xaikrDn8Dt6/PQ2uNK31pv98b/el5deDUhXi1JoHmWfeAHmQgiU7nTFZr6KI2PO5KMJ
D1V7EB+/wNfkTyu/WEz7LZa0uD3EUYWis+Ghkj7JjPcZYz9C4QJkXr4Tpz13EBtnEZjBCJw97Fqq
mQPlPv/auM40WbMJO7xrBo4GCV1DOjgSI5y7faytJ6YzYkK/Uca3HM8kSw6opPgxWEeazzGr8RjW
XUuAJc4475hYrA/Kg7idbVkk603hX576qtLNSP3JjoOgFqbxJ/sNL8p3sM3vWrpUo0XuxMmukhYX
LMfUiom9iN88D4izFWHUFC3YEucYn/6Kd8pri8dw83o0BEdU2btR1aAJCBU65xmsN48oMoq3lZ9p
3nh/t5zWEE3m5I+4WfOoXxucQZPHu11f7gprkGOWN9+pCKtMHbcdkNVRnJyh5xtpMbggZnJG8sZl
lnaSv6LajJ1p6Y1Ks3x2yafT9piUKk88gETE7lujVtSke2uViz1mGLSmLCgy1Qo8GUQqeUcMvjJ2
tv1JjVVsPP5Sr1igyjyjxZiUzCdhyZZq+XRMNYrhFmWzEcGJDz+pfC8fPNp6xA42NoDxkZXsURq2
rtl0rPFPUH3CjrQz8Zgtkbj0NnPYZlXyAcfcliy6yrpvomS0+AJyaP0seZT2/bliEvfbt6sLX8o7
PGGtOV5/ON9HzAPQMVwjIc6BsDmQ3PHpTGJyOWVYlLmPn/PiLGLwL69uUWcFHYC+5qXwtr0l7GSC
NFQTJKKSsSdS4PylWAL32S1yv+UPJcOlMato536YiJ3NBhUBqzLCwOdHlE00UAlBZXovdoPvQodm
VZ4zGNjHBQU98OpUW6Mk3F0Bk7EqtLLfwa1hJDrkg9Wg2H6tcuV/w1odcybuziEFK6S7omR13AJg
EIbole0m+qHMp6kBMaLkH/V5fgxZy8eETAbOIX9RbckFRANY79mgi7p0eeyAjNb6vxd+z3+eP2NO
iI/EKoRWdWSTYEzWzGsE1XtXQR889zGwOaW79vlDsdpLW/XASBfvbOvHqxvfyCtO7VgrHT91dSvC
BdDw+fRUEhZOAZUlc6GOafO2oiYZXy5I6Z/sKZSx1UDgUG6sM5eGsJteJnoKTHaAIdrwx4APzMQZ
ItCgMiJgtYzAt7yow+Y5aY3YWcw+T0O1Z3x1jNtUcZZj7LGSu5+lSHw+cc8w7W5vxjn2vwKeYSHG
Z8vNuW+0BG1MWGXqgBTm4YEubSNWF7KfRRHHbXhriTZ8MwRxWtwxfE6dmeRkLZr53xZXIoWarV/Y
axOvElqVbWdf/oAx4Shfmlc8iOspwJNG2zZWZsgHqpr7xS6M8mRxqGbXIKJYNjvqfGZMZVGJrChW
GGHboFcR/VJNl2n2eELxoYM2DeNa8ZWfkhc6pJk5o7Er0Hy58X3Qs0hO6Z2cqqzraYllBxwivrAY
PHZqmum7zCtYlqXEr6YlQ6g/GtfNP1NcmI1zHiNTVLlAuMn1sh4tuepmB+Q/WhJpLh5g6+sM29F3
vk/tNI5lXQd/bUTmIPPaubuyfQ3zsm6NWCgOa+jxviUYXi9xmEkkKXjWcLWFey0293kMJOUDqTXH
YIlv8x+j78OErTPgg695xPIn9mWJ40/3vOiKKX6lc15rOvpsP1Fmjtray07ZbZEji2MahQzKCF5o
Bkvo9WiQU3ZGEE7lgwMSWys2c52XzYOLyQyVVPTGAhcTruKBW3MkFEbktR9uGSxsutD8COhbxFyr
Mnm9e6OgE/uRCOvJHjKFDsKuqDhZrwYjSDtUG/6BM3wmVoeECrOJOb3b4qwHWU3YesdUH1eaqJLW
Wo4VbHUPOMzYt/U9uw1JRlWRjPFupYWJGFobLIvERFOEvU5rIwSFJhNFrknt+yNNpyh0rjH7m6Gr
qQ6YmKz1514wJrsjLOBrSOuLmX4FD92T4wVJDFdR/yFCfvEi2QQQMNsQYkdlTqqEgYy4gHjJ21Dv
e0L2tlPTCZ9BJnG6/JW8Oi5iC/xnU8L24fPnHE36Bxt8kvye0b4XAvzUGfOwc//QRywmF0NgY+ji
X9S4V4saEIBh2Z3aIlEnBPlF8aisBk5B6bWj3S9NFDjZNe/XX/as12FHqVIdDbV3KrGUdo+MXD/z
4eI4k4ci20bAgbSqFATIjrvpIyABaMumsBalAgVpDIrQfFFKpVxiXm8LwbTROa+euy8z/1C+/+EP
AaqQcafTe8fZllTJBOqK+fbO994LXf36TeFTAsoYS48uPz4hwCXcu0nA3ATyt/0NsgKxBadRzKig
a6P8mEijqyDLCJY2Fqhv01nReOQlLatIonw46I+HJGhigyH05X/tOZ37t0zaxQ9buj3dryih4t7f
8Q4g7+mbIcPDvD2EQfubPxMPsNEMaG1ypqO79lUUwU8vTr6cpt1G3ileuFwSyT+0P8E/nBW2WY/O
HzIyfu0rlDysIstel8ulCUOTtumGXjXuF4XPPeoMEOdw9rACH/7xzvgsLAfuwNKzB7pQrE8al1r6
JVS6OzHdmOdX3JeHy1c/va7IvlCRJ7rzNglaiHGN2AN9O7r24lSlzcs+D3PMTVmNFjlZKbk5+9Jj
ZUg82QuzTQKE3NCi+bD6+wSRM2jdiJzHxdD9jTnQORPmg/C3QxwCWRfu6nAdeRYnI4cjy7ASqEYf
ACDAXEagK2hMYC7FBieYxU6+3iTbUJP/whpk3xxgvIB6s2wKVn7LJqPI2DID5gko9dpv2fG1uc08
bM/ejTWzjzbVbSva9aj+i3EmOEXDfNGD/LhU0NRWr92qa/KQ2FT3xBGvgN6znwXodiA6cIIO8LGd
SG9QjxLRUMGtNd9nE/uyL0PYBG5m0iH+YGdOcuoBeY+ooohZcfw2VULgD0Y6M0o3TayCP8mihsiq
VuUfuWBiDj9DPZq4+wYbtV2sDvwPN38rXwPw4ENgn1nETITs2zKpP8knKhQGR5dbj/VRB1js3UlL
G/3IzgktRSGhiFL1i3lWrYrmOBlgTCIWyI5MmGThrl1ipUOqfrrQ7AHRxYFF0XXz1bDWE4j5gED2
XzbOxbS++EOk94IPzFBDvMChjy1WdmPUMfH7W8DOeXsTM/UxGRCW9aEiuKnO/9w0HjjEMlz+a6Cg
+IpNYHNmJvIT8LXa6e9nKdBIE+puKgMZsopoEEiWj6adhnxH1diq/rwfNoXjBkySfHJrAmDsOsGz
NZxSYe0VHzOJPSz7h3uRJgeAM5RjdxwUVlauDpwDQ+DI5EAkLm3EFnRljKjWlHqU41XfVClGWZ/9
QdI0xp1Rd5loMTlPIRgZ4bvvgAyqkP/4rdEOC4HmypcIhqeaAoFint4HmWkfjstog+mvPEq8ouU9
blKknDGregyWpy30BcDR0hXx+lZRoVAUk4EznhsFMapMIYH7CgqNlbtVJAxjOF6qGQi3qAMGF07Y
qdsX96HIL0dbhmaJbxB+XWtxZ0lhIDaBaSjWT9T9KQWrzE9ZxXHpa+l9n4Vi7R6F1OFquTrEV1Re
+XCUsBtu5VUOzuKnuUe90soeQtPJ92TauPha+902RyPxj/My9/3mfQ9YTYFfA1Qz0Sxa4SF5QsMN
uP57Pzc5upUWXefI1sYvqruKLN3hE/8Suc5fcftzqcB45XDcOy5/gMMxqmvdyQaIlZ7OWcqBIk5M
+/bk2GCWwuvdCB/ycqJ/DHFPkatfjJeuQRdzCAkRf2mpmcdPty9ez6IaRhkgiTmmEskjv8E6v6G2
KoOb5/Vw/tzxu0BwF5HkDH1bbefLRUrSh7XsYkXbQLqR+J50BAfIVW2yN40vYTCphSG6TmQ0CAOh
S24SX9nNP/xShYNHbeEw2BdcB6cYFYbCxzeqIkXCwrqYYliBmSutJX5PglQQkrJuNo5SS0FC1l7h
t4NfaFidLaXbCwvkC0zsjeG1I0dSOPs/K75JVD7tZxq5n/b3C+tvmkJMBAu6HSjnWZfulfJADMMK
6s8QqOQ9F3KOdxqwJk7Q1cKWl2P4ay1KGpXaD9+Db7QxU52LmnuOuLPrDeReS6tgTGZ3983meLTD
HfuPpXwXBM37uzj8Xv8nbArift66nYFuNAmczLTXlmZBSqlZsNyt/q2+0zkjLbRdkGAQQYNgTi2U
t0Xr2u026Fe1BhVSsJByWqLlLTA9tNRms+GgDHZNZJnyJVJs+YVeawtnHvQdSB5x5wHrzZWDrzPK
2VNQ1joIibPH2eAnjEO5zoI1QrkYQAdmJCd1C36jg3rl2XIz5Js6DIHwDJRVCfiqvNWEMb3+sKGz
nNXljaS+f4BkrdWWq1AeNlTpiMCqbpzrwQGbfsMM/xDQzQC6x4wIR8OEFf/aJbycXxAJ7Iolj/d6
rMfjOLC0rgxCzKnVu021jFdZ/PPh/j/wcf3FCz0EJ8EOwHS/T1P8DrFhyNg6sg0h/slst+afmmQZ
hQlTFg8SVQ2yvHfa7nK5CfQn1L7DR+W6JFksmKLqLyCCUuk6SDwKPu7RtT2B8/FakdIp2FYGt5Tg
E+m4i9nNSpuDpTyljDbyeFUtIAKtUMWjYhNf/eTnzgaE2WETGJ4RiXERadpotmdivAndWGoXEv8V
JAZyklVgkx7+NrnaaG94Z58xBFW3lK+wgF2UQVs2yVinMwufg9WfLi5QlYSIglyPtBX/uesqEr7X
Kpaq2gxI+f3MquwOWbrd6mn8y3XceA185cQRq1IqMrdCl8SV4EwSQ3p0Z9/x2vRLxwpAV51C6ymg
l8LWvcXaFEOKoHMe/HbuAiXVjtjqdXnbraliX32xUKMZsHtWCuQbEFuHfmaqhygCZ2T2dnZYz9Go
acHKBNKhazM6T+oO7MYIINLndeaHNDcnmRdHWotmzHtCw3DzuvNFDZcb3YzFjLCoMeMVyKRZ26LI
qRmfAgRvUTD0Vi25rwx6X+Q5Ss0YjD7QAEDqEwJOt3TirKGTgymVHmcgc3Impvji5oiCs89VZxaH
PovQL1z12SLV58EIZXinSE11bbjePVUHaHbJBHEsbMStd/6BtVAGiivxScpEiXd1d4WFkS9Qnusx
bUCnog6zrsgn+sgUT18ZRCmFRgajM0PDJ42lf8jjcwxcfUHO5gf69LEO8DvrvX3mKGCdCRGmIHjL
98Nm3/k5ALqXGwfCrE0u2DeMiqZ43rJ/SDrKH2JAI+lYL3IppTIcPc/3DXX4Rj4FfsbvN9RPHiJc
A+4Jyu5rZ2Av9a/X2lNGKCZqaZQe/jOfZg4TH4XpW50RULd4kUqacnsPBp1zC3RrL0pzWqAIa9kC
0LIS8xEC2n7gfLN9CEDcS87kI5k5y7IuF4TBb2p8jv+HfrPpKKHP6vkNQO8kVYzEvA/qk1MbDuVU
ZF/n0RixHFgucm5eo7BEZWyLjudhp05VXOn8bjrkCNOa47MQSbGp6xwCp7tDc0hJ+5q1r36/76Td
jfSZlGh8TzO0NjPv5uOTt5XvabMFTtNEJdA+gV016PxjbEs7PU3/lSmFcT/rs5/wwAPgD7mJezml
TVazJ53TsDaFA+VqNN2Y/aa2RyhT9JuzhEX5DzllNDO04hHOLK6KNqG+I/Lp6CfPfq7M9kmSYx7s
em7iOhL+U1PxVmZSFV48U5vjSRZzy2hSXrFtMKv//ZXAtcjRQ2Jo/tqzv8AQwMtiA65RAADMxKee
+o8kCweLstR6vMgP5X8LQzGBn8/OIBgHNzFn+ZEQlNT3sCNHIejr2JcDtSuld3VrwYlC/VDIJNos
JVFnfyxFHVmO+Zo8dMNNWH7qbPewjMnwEPJ6nUDMnp1HFmR7pNCNVkHoL8750Yi5b4kAT3+m6sLy
vD9dhSzmc6THK3/iJasUxLj+bs1dvEtnHZCJdyIYlr4vdRoNIcjFY9VEYoYAlbHU3KA1QrXj7415
ROL5OuQbHQjxS8u2hYr5JiLphyW5+jAkG0HMuBiXXmBZJ2joPCGbbSRYOC+RPChyaKMHj5cAsbwI
WDlpYafMPdVwpUqFFlIuNeFerX/+B9T4DlesFBWHLfmUPQsf2XxwHhaJudiHtggX88WkEfrfn5Y9
daD6PaAgbsFuVHLsD37nTxyIIfLH+2lMxupFksFaiYQ1LZMVHaqP3hwA9fKfOJKv37VWofxcwKmh
N40vXgN6XMWt3+gm2YxFJ16eqEdDucGuCP17bIIzMG2ZpjwllpyQAc0smarqbtknrSGrWrXC65ph
GAR6/Q3sTROv3AFroMIbv8OSokM2YiwyyBmeNZNkDaOY6J7VgqgmlqKLTx8pVtArKqI2O69KRaJM
U7Nqg4wKXN7Vr/S26sWpQAoKJQ6ns9UlRkcgeTZdY1cywoAXNHM1CfhTDegEexRFrzJxBCUwrpe5
2mWwbqxoUnrsM0aOezF4m6wy1xpDtNe2f9gPNR1Ym/ph2aF1gNPhe7MvZAdxIZorqLto2QQmd2JT
UkMxRjygjRI3etDJwdP6HygMYFS40NHgnXK4Q72LzONllCTvrhS5baOICH23IE+uZzGAyFWxGRid
1gLv4KpErKF+RmD8N3Rs9oNoLqi+KZnEErAjEQwifNymP+k26Yr0LNxmz0Ha+J4R3u4e9RV1Dnnd
Vbrm7Vs8bGMvMcdk/COIJHrTZdNjeWcadoecPlyoMJLuLfOabGCRZVO8Tjp3gPTiW5Bz/+OFlcTS
hqCGVZY8WkuZ3a+8HnQ83z9TFPHtoAORZoEJ14zd+b053LIR1UdVRWqx5xgtLA1jR8Dg4BvaUy0H
J9eIBZdJ39K2GR6vzEXH9YpVPD0VYVrxJ14701ZgYrKe7zIlE2/guR2UJobwSO2qKEEMQNYXcHlJ
wP5xVWzggVe6JXQInEcW7AwRWW5ttZZXKhwlZwix6GV1oxXIx2rdSWFScN4QNxB+/MfSNOFi98qX
/cIimITPYesjea/b5H0a2YeSSwRVwD6wAWVFZf/8A0AkwX5GW3Ki7SvnPPh/aekTvV89nNMLp7vB
+YAOsIdedcafL7H57TnytbybJd4TlNcv7x5/JGnllaeP1DWd773H17zu+ZCoNDK/e8UQYkVpeCfa
6sOMQRSLs2H7FVUPoz3xliDzcbvkDUS2Qk8VZ2Zv0q+miYh7hfUt7zGZ95B/CENOf7kvH9fS5ChG
3GJN3VPIHH5xmXPmmnS53no6tGRaC4HfPgEzSKUlVe3DK7km39mWnDPE0RWR9s23MgePJU/I7rpk
B5anG6gj4nHzVmW2ItMPFKHYyu4AdzG5xrgjTG6Q16gX9S6gMfO4gZpRlpra4uEFKOmPZO0+vP99
LW9mtaNIMwamgaC6Wg90bflfQrhzu6P6vAU7zc0z/ivxoFtKdTWiOGKuQEyRHdD+N3devPCv1py5
pJFmfSH8QdbNqCzwftZB+eYjeUjtpO4eOnQNrU/a4H5g7Y8EkF2Mv/klmVEEMKXYrfwWxmhOzDPZ
+Nt1Gl3Bkbp8WkY07dGECt7jucp9d/ZMX/k/5hufCHDxM3lrNYDueWYguEJ20BBvDeV8MlVuWuiy
c9elxeEzMRfifObLvgkh7AnMJmhdtJ+Gt4n4nRNPknDC3R570t8j5pNntebp/ScW1MSRuTibjOSE
JSPVW/7nt1Nw9ru/3l9rwd/g1h89UdCDE2ao7Ji2P/i4UgI0hGrWOfMDqmoItNWxb+TAGB29UHu9
l6tU29B4EiiMH0JHY346webczBCrT1/zl0rPDPimA0m2nzZNcLiPHgBJcTQALX3Yt2L9an9gLq1V
Usq25e+il64xo6RiEeH3oLQ5JOiGOuYeOStqdBrkQeQjiJGByCoxr+L1nyyU28leh7ITlaEagDl+
Is8bwhpFGL03QW9Q6ughvPHSoQRaSQ8D59m7Qr7cldj3T1uAjPb01KlWJWaF4vTqfFLMkjrVNUYg
u6OZ9fMriaSJeYe9cabBZPoI2TJXvrldAIdj4iAEg6L0T9dGMLC546ooqoumANUXP/LL4iBi5ROv
GHpPlQ1gPBxruwZpVtJI5fo6I90Mx7uWsZwh7l71FFUKI1i2qJMo8LE+vSxEMD7+jydyzzZaKRVU
8+E/eYTtnVNOy6trvVASoPkcxh6mZZNCqQxuDCuBUNrMmkTeAwmepTKt0Ov8JwBgrPqeelt5m44x
Gf37T8WS3r+nRHVHDFRsp01I6P/0YsMNM+UhjKa47cZ8xZOgsrtWtVqJleW3f5cZgtvHCOaLnK64
5GsBYsoTJBktQBnelxLmzbIQX/cXbDVDHAQtDSMRyte6iXXgJdspIWXcZLnF3DbOQJ7d1xMqvDB1
3mmgVvrRGx7wbOXP+j6uCxnxP0zxmYLZA9adlslbLx/DPYIAzSzTwZLPnlu7hINtuegxACHBjmfB
+ba6SPjiA77j/VMQgItpMoeW+NtfKd8NTUtsYsxV6IFKdO3UX1LZNNaJFLpTqWuCdXswBOAZRoI6
zP3Dh4SnGsoFjXlSA7R0ajt2cR36fbawZeaLwMNIvuJEws46AuZQZJ9X4lJzneVoMUgGH700L81D
OF/9tmbK1N+dpTZzjtaMIyRvNxhXSo2xXyIvrGOzKfKoUFLSf3byIVqObYiNt+CvbvREmFKBhThL
5V1JeAZNfnz23H/x7HVyLr97E3waRIn2y5fZERFB8ZDOKPJ2giY2Fl6GOAvQClwb1LaZkB7nG4VD
XWdKY2jjeOJH1kqWnqCQg5iDhLHRX7y0wW5l9mcSemYFTIuURX6IAvhUcJt8Fytb5JC1EEq9z6CP
Kc2ZKjFzHmdpB7Ax7qykX+dP6+236v96+e8WZj9kNplZo5h0QmBx05d93OBdox8otC6DDlaKrARj
RH4JmG+dv1/tMWhPfb3XhtboccKekz2sD5gUaF5+V/EcGgNauikPS8GDIVX38VRwsuudssBVZlhd
cxFYWMTwYFJXIUclP/OjFhHpAqA/BqCd3iQeMcN+1GvIpqoD9uH0Xy5bNlURXOcKy+0BE7RfA1WS
BHffBjFS/K3/MQVlh1MMdsAW/5OSkTNmFmNTz9vC2K8vdz5I+tlbT4c6kCOGek82bxQjxdj5jlOS
XRfcHuuJFq8LgSzw00xJ98/g3qcGIq3bYHGWv+7z9kj2FkyG8+imHhTEIRDEIk2fYFceW357MVtE
BbNK+YZS8Hch/qLLSFjBTW4OIrBjvn7gddjQanp27spnYWh+W0WbCQXWqtd2YMd6e8mGl0OBpy/b
EniBXaZi974y2r/ZN3o9k5RyZSYP8jRhbJyof9PisCtHJdQc0PDsIULW8ymD5sPZELEFzBIkrS4r
J5PgVziuzAifJWN40gFyJMK7VY1AOqiXZXgP2VDhXDESRjWqz/yXi3FaiQ0wCEUryxNpDRP3tQHt
ndnONRoEMNC1OR/JfjplqqYtYlDO35YT4M06h0hOOgQeRW3g3tqov/1PS7ha32/NAL5SF2bpLPwD
7c6gY3fnmamgRlkhC9SAqGJR9UqWL7M1NSKwInvAH6SZUrPkc+fQSyq0jDl8FJa5uhPRKSxWF1c7
vb8mtFQCYvEM1lE8YXCrrMLC4ZAg+5p3KTZuZxpTUicnDIUqBVynXXQQheJUPrrswVWrop/XEW5n
Y5QqYDvoznVd8vy3C0hdh4ehWFPQhqciKlbfg5E1xhUgecEZYa7oZLsR0wqWV1UJ5YYT4xYaAVe6
F9uGM5l4ue9TMXKYo6nmHizUGIEJzIXxA3UTZo9V1seiy1JSjeW5b8IZd59VzmbfnaLuRw2ByymB
ZwxC6nszYqx+LZpI31VBqFVYbqUOtk2W1NzjsDqGRi4GTOJcz+Hd32Mxv1Zt1ycyPWfbweTg04G9
lE3ibSGcCgua1VHmx2amAAGZD7z8Xm736sfbhvfZ4kTR34kLpWgzWnRTkU9S+38JeVTEJtQVLxt2
dY9LwLpSgDmyA1o0uNCfHHzcVabfLONKiCQa9H6UF1vEFuR8ZrgOV10C0mSLyG/im6Os9cjdj1WA
C5wRYYu9vk4m5LxdUJnFfKO/Otc+Lccu048W8S+DlONXcAKS9jNXMzZ1oJxyp67P/d5aihjtYci/
T/P+Ft2057dByX041lB0Np+f9efCkU62+y02321UAPgGuEM1JHYx2roN4VuomvTM5dsGyLfX8xsO
tQy45C0Z4OAj7SvCb0/XWHZF7GEPjUEmPDoeGlrjGmxyGeqSP0T+Q6+jUoThiBwgzPuUUybykRjG
8YPT5OvNQABxL9TLT+meKRYiEdBpUgQrpu7G0OGhy9vN6uXjtcH20cvdUN71MQnr9WDdAG0TvePQ
lwKWJzKaeTf4CJTm6vEKmJNSraaRRMumG7+dIkv7VPUK4EC4PK9OZ2CMn74jpm+SWUefuMHocRns
eKI2G+ERqmliJhkc/jYNbtc9c2om5oMBxz2wq1QF5+qMri+MJD0wPVB9JnOjr0fdHl+ERrGhl0sQ
okj34/MJX0RHLuDgVLwF1hfNdRY53usYHSsiPyupskMeXuk+qnv5QCTHx1J6UkuABsv0uwwhx37h
dSXzLbxtQGonXwZ+dy+miPiflotEHJO0XV/GUR8E8nWYWrQKF5IafCHVCQpNrdNlkNtWtIRwCXGQ
q9U5j/g7ZApBvhfh6H8y4fUYLp1cdOeOEf86x0Qj0RRN3bgi0b9TEsimB5DmK2ZDd1hKww+VfqzQ
H7lOjMzyBC6cNknI8F7u57qjyWHOdOGyrYYuNxT+W3eVx7pesP21Iog2BC9XX1ZInMy4fLqsITMw
7q3TVFaEpCLVGhh+65d6B1uaUs5znoZBm5MfDldxDCSEZK2eL0UDyHObUhS3gY5KxKMVRHWM7Fly
tgDfKUlbP9CoJPfydP89Nxja5jQfGECCvXpnKvzp+C0fpmpnRXjTSeg6KQsqQoSooZRiD0O+kuEQ
dgKI19QY9XDaS8eWc6ppHd2aVglhDYdusGD1JX0uDGlpWE2zbO+OrdHT07l/x0c2kN7fkAC6LceQ
Hgi2mUUJ3H1VRiVJa6T8FDPOR5ys7o/mOxqiBOCWL6MYBPNBXzihO3ESJFnZ4OHJt5AkC/559I8o
Gy5xQ3+4xvMuM7ZwLNBKPLdJVWbYwIPqwqGxYeF7n8eRoz1oCC0ny9dzJxScYAAD1PlqfV9cvGSN
nKX5+XAuSBaeMz8flOiObjpHzVqDSlc5LypqF6+gpOrE5ZqkK/tIPYG0fp/OXRh2n1tc3cvCxq8e
xBzWjwP/VyAOAVJ8I58l+sr0nDbGw9OIVZQxGknDAExyoPOOdDD0H+6qxAAQkIq891O8qPYScEw4
h4DBbK4TMAMpptWIYIF/wcXs8Yi4omVE0AlMMh4T8trCEKCg8/6s6vC7DrNWWXP8rVt7FpfT9PQ8
ZX6zoP7fHeQZFwf8QTqGulQI0MB6rLYrJdntNJMnDBozn6nsjWWSpNY7tBCUik08EexoAsI+tDk6
C2OaSFy+kTBCmGSUeTv2wgQ+hxuroFm5T8B7SM2LI+ryYVQYw1sguzuw5dYl1sesclzn6zeVwAcY
dpYc2kL7YWAel90IyNoW9JF6v7MP8WM23WKLXNRZyzsEbtgCpeIO5Q4BLwLNpL9829DqxxH8hGME
oIqbm1l1UQRPoQOm4RGej/Y89HqbRJDu72aplSWMK5LZ6XMCbDyWS5ZzB0m7E0CdJ0QR3H+HYkEK
G0egWv0kMZLvU8gScp5eFjtu5Elp+tPjQXlMhIIJjt3PQ8wQOs2JLc9hoT1BbT2S2hCcukIE9GlK
u6e7wIk50XbhhOqv7bn0GS74IIMZoF3AUWvF1lJVc5aCitDiWxDL7c6fyksWX/Qmpjn3aGOFdydc
+UW60bzObFZR4WgKigb0TlQpJD59+48TMa4n1d1h9MCeVqCXQatcEtLRAgcIdIF810jLLuWv506Z
g7YTWCpKQ+Zd82zeLJjRW8quqYgLcYfZLiqJgnN+UE4n7E12p6ulJ0AxNHmXmrc7YiRJ1B6+ipLS
AOCxUZeyvPZkTxWugtp7zog442G3JMSQRlkqR+FqbFZA1ad/vyMrZYfPmOIC1w1kP+u0p2mjPM3o
9K/Yq/JW+ciabxTUVNekqxzhhCeO1fUSv8UHOE8+x+eEfa3F70CEKTWemkfSq0j9gqJaQ3EL9pcS
4qTCsk6T1RQjYfbNV7PEZtYkFdKvFumKjXh2WrUH4C1XAQFxALcXAQ2wbAHKUE5wfCyKCSkxn/om
6E4gv43b2hcI/Skzu+LFe+GmIs742h0XGh5KRpV1xPad9rldn98uSpdaGsQTnd5soPB1PWdwgEB0
Uq1mu29L1OnklGBucNFhFx5bQzMPcSwIz8CDrYhj2VnEmJVewnj+EIcmSxXIWbiuLsAGsfI8mwhw
xcOFEFedOFYhibYeXDbYtCyJPIQxjsCMxEyHcL7euJ+uEvoGEtMyixSlR8vOhSefWyddvHJaN1po
wTjFNQB9tFiLtqcm+Horxo+Q2JFvwTtY8Ql4dpvNX0p40EqKqrY0sE3aMjO2QEd7VdsRh3TBv6iU
dyB5fyXd/vMcJTMrV/HkFhfrPCo0XYiiXDjmNQrQRf+sSRI2wMB7Wrht7/ALmc079f42jIzRUMDO
Z793lpXj1ZMPtCQvpacefFrOkhUwOMzaUR2CJY9GdvPvU/hnb1DAM+wDTY3dy13dwPYSNPU949fj
QS5Oqnj7vuq+ytW3VdhQC0WtdfBm/czpR/TB/g9mCYKzZ3ZRUcwNEbT3WkSPL0aM+XIbC+qoN5S7
AoKFB+LO+44xZ+vZWp5dI/u9/iLw75NYP8f9ibxE4mZGUrWM5Ccgc0E/V/7FxEbrcq9lMK1NRTNY
MMdnwmc4OZi3M252sCNd075y8Oj1K2j7F0iPGGh/QJkYojaLo72AwZu1s2hhhdaBifxwLscJFM4n
geDHK92VlS6HvYBAtgrGKYjZuaVhTQqR3qQIq3VI8665Cl3eyf5z6ygVvYKm/Lox3K+9CXSjGWrg
pss1x6mPErBISqCqHuMOQC2OrIbVSjSgDw428cw4D128xf6pyFj3iokZPQgPj13Ay6LOpQ+C/rD4
hEJwx1IrD2VdgK1ekiaX6IsR0ApPwajdnxSmNW0e0DegPvysCldtoP0dO6rRfzpxuqSNtr7BQ+gi
j/10vzzfEVzeVkVQ88aASFu8X0n+XRpPXJgEqzEPS6EYDUsRBOx5JvK8sw0S1D2ADV5oYTbt2OSX
rC5pe+5gh5dgl1h1dsgZ+8C0oXvF+qdt0CMJ2ad+GIX+RfJg5l1yzsQotprcDbaDu2jIpP8fkUN4
4EPadhCkelk73j/xCBaea5k0qFtJ2QmpLoWntMyD1DK77m4DmWNLvHVsF/DSmbzQH0Pd9tFUfiWT
CWd+DWZPinwJTeYOlCMh9eyWbrOEMzaAfa+NWwH7hOUyyk5dlrix0gJddwU4dbWdtQvA5g5ifvR9
2zyHf0+f0qkqkrhraAM64ep2AzRanjaBI8m8Yja1LcHnDC+LTYp1fvesAA2hYVfmldbDd8vfufxG
MOkL9XXLe15h8YqNRv6q2N+0OVlPwE4HWuw9MW88SAszE3vKK35oEuxKkduVuG7oWpgcfGKc02gJ
a5TqGGpPYXZjKXzDrWpSdjN6QBDUQ/slqc6ybiq4GtwK5WSchRaoIkXrWnlbQdqUepOZHb7MlIzC
Fw29lCCb+ZVnRb6/KjayzBirBwg6NuydqZr2NWiW4MTTYqh19RIp7vaFybeJubOgyq+5TIF3EvP6
3sjJnHyZHH7T/EtzEFK6+zIWVj2UUHy5AJu/coY4yUzGQhmsD3YZUB1TGKDL8TFVN6OTOy2dUJl+
vsTxRpeRkyd4YQ2Q3pK2Bivnrb/adpreW1UGGbcmJgDnPzZJHKYI79qme4SelP4JvoMmVnCfyrrP
9pH5dfwA68IQQHtTpG5Oy5k7ndzugfg9D3j9O57z5PKAbkVq27ziE/o3PLNoc6rJV97EH3CrFZCa
zYhV5JU6inYhtcUM6bfRHklZ2tqlWoyEQeAZo93jl4BtjEnBBk2Vaz1YUeMUVylmMRamB9nxVdQI
04aEKIbKhI5WHWNHhoHe60WENDG/zE6wNik9KSCDLD/44c60O5N1/1EeJPRRK/nb2mORyjyNJZxi
hagxabZ33R04K28EniR0KR3PcqrUuMfjdKjWh8AXEiVxRIBx/d/N2yUpxkZV33FlAf4XJOMZ6Am5
5rYbt5GHygy3n5I0C+Rw2so8Xo7LiIO42xV4V2dlscxIMmegdTBSI0wfw0WMoAWp79XFNIFtyNFU
SdrwC7UKoTkEbanun4ulYSXIDFB1zI/B0uNGTjSzHQvpl6u6yVUsKyJIWolB+QGL08qRoKP82BdJ
quLlut9k4erKCE3yfHtzOV4on68SZLQVoitX/zjewvswSMRWflu0Ub9V7kTScBRae0tRlcAjNt/q
aNuodw3fVI+BKhw/LLQNyU6IQxXECSO6a8G6oWMm24Y5q3eKVKiygwHyUasNJkBpxyxfahErv+kI
7vLrVnLQQaufsl9xTVjuuOSaBSLrq5hHmGY1tT8HpwMdFG7RMPBYUw06Q2UAnMGLXnnDTCIGw5LH
cFtMOMuj6BwUcxtWSdsMLcK1ickIxuojB0qU7figq9uE2w2PdxNzJkAx983tdbXctHEZm8ZISsoq
vPBaw3le+7YVKMznh4grggSSO4kDDr1PE0RDhuw1dvk9tZnvV5SM+ry0L4ZDLhwTTDj4vzuSMGrh
mDi5w9SGfx+83Z8JV7SObLGawzgx9sEkXEu9hB1WXoy+NHnv+fUEi2cN2GgjwAQut1J35K7e61hC
Q3NNXrYmiG+Pd5Y7VWFbtbtBA9Ma/Kxz/VBlsTH/Axw+ikebLsgMTqLDg34BbRyAJvIpYMJaOfaE
Axf4VjK5x+yNWdJRuh4pCSud8KGPOVj4OT+JZb9ePxd+t0x44gGmRd74YlHFsFExI+5+Mcw2HK2c
1dHYCxITER6xpnPfbrR3cWJS4fAa1RcyYYeqbCZ41mwbcHc4jtMimpJlpXvv1DULQBmS7mPwXkh+
H5ac1UfnfYwaPPZlBjXzpFL2mh+J46Rt/dUiJrOvU9FyVldN8WtlPYJQt8yd3Meble8UiYJKyiXT
aKlY0RYFi+HiHO+zC3EPFKaEq1BpW8asQh0u0yMg1cuHdOw6c6gLlk4v77hXcXvBsv54Djcvdeh/
bY8FO+aWiTwkpwKvAdbzdxakNDx5jxQaFCXSnEkiaHjOvHhjkvZJgt4b3KLfE9fph/of072c0CyF
jmVATEvMVCpyURhYbnKOqJpfbRjoYxCr0OpMgDJT/IEbIorPlEYRywQhbadfPDPCXpn1mbDzcHE3
KuKbipFysyVM6oS6qP3x/+cgsCeMXV4vN7NJv5BpcYeqvBV4M++vev1Sbg6HnOV8aoAwBmpdjkgp
GCIDVVgusuAZyejmo+QYfJZTC/xRgWEN9MxeIv1AjwYK1KnGqswpOMH/kJKpJGekHQJ+XfKhez+0
/EmMB+7/gy+nuG6DwOPIc7yvBnxBeTpq5vLT3nju+kHb1Riz7Z+buS6sPBeEzQUf3NZY2gkDJzW3
MPa6d3C4u/6SOA2s7mM1KjDuffWaZcZ+26OHGFSzx+9HyBFud9oP1C5v6prl0UVyv4gPe2ryVt7e
UOCwdFgkuvyQwqvq7Tb1yGoKOyIwUa7VkGDR4AGjfk520+w+1vNa7OBXDZasV/glodD65nCfAdRK
0f3GovAKUefAbjaZHxF79A2stXXhRZIjiFVIIHr+V6/bQr2YP+qcF0uut+JXZUS399igiskca+8M
ARZbOqJpxXaESnaNdx6GJF/aYRAE1AlE2phh7dB6g67GcQwubdZay+9/KvhGAxHMl3NiZtnhhVlg
819D84NHYDVCnTu/IkeRAGlGALFWKNp1UqVdYfeYMJGj9xEbLx613ckpY6BdciOpz21oMUO+50XP
k4A7Ti1F7jlfAwNiRw52/FL2B00jbhIdMiRU17mfIyotRK9dYBx830mcm8SstBNNthOJxppXwYhV
EwapDAJEiMx2wqfjB6rOfY5PkF6KPrWZxP/f7rjqOFaR1x7NeW60DOhoECWsk/ICMWjLQKsaLvMR
M+izA75uuh+Q9Dm4xNK5Ej4rnMQCIMK74aDrtzpRklgGL12yg3mJDdu/ur7vZ2u3uwCPC1JFHolJ
eiJDpU5qeOePCR4Q4VOJPuO3XLUdIO30Q/0V7ciBP8oHCJrPWvkj42a+KZhbfVZJ7llEOQO2nsVP
DkddF0HLZIfjEVJGfrp31ZrgNxrXg3qDIMGDZq1PitcW83cH/DI6omsOTeUZyoFuY3tZJ6KsAzNk
AOQNPPMFwyBV/RrW3sdJItxPcpeujOkUCK3wtmuWad5xE8EuRBnVAJbCBnWf/6XIJZIfYVGeDYx1
uwotojcStBZie8uKKUFNfk+HYtlNP2y6ogmEPFSs7Ikic3+pODGc3/X6NZMcQgw2W7hXEWZ7GZ++
Cgb6FyGN6N+H7OcTRZtkY+xHGqLJWs9by6YtdI7IJb87DHaMd1uzFeBOLc5qB3FZlkKODbA16ZBM
BbJdH9BA5axjXWtLoivJOGAs5ZJra9XfUs77Lw5iNrizsMLJmDAywNzvEp8CflidMWC6hLEAnJvH
AlaBswKuYHpmZdXlts10cH9QHuODKmQV/aDKidWtue/3mle9FQH0I0t42BRlIYJbm+Z/HockPpl5
lQY5tGEEeaGDAg5fMXRoSjFJdMN9lADkF4Ph53HpBfdwQmXYuCHF0OjByFzPzZXDPu5yCN5JnPnv
0Et70AqQQfF/1M4g7ELYvr6Mj3oNgnTqaS/XHeVd4MBtuhjEuvJ+3l4b6igF0shDQamSh4N5Waci
06fX+oQy7zyogrL9c0Xgn1jWagdJNvBuvA7eGDNCaqbNVqJm24LmotmaU5sylyZ/otMsSzux2TRV
u/K0uwnDUp1RhHgLHXJGFYKf+pL7m5TtDBMUrfmXjb4IzHfQ9q1TsgQhP9SYBb9ElgKoyaQy3UdE
GnQ2BDaPzSlkk/jXcpRcKjomzj6DbBIluSeUBtuYmmH+FM0Kcq76JBQ/c7YphKgiKJEUiubrZLEI
LJuOwidwWWxnO9xLnIn22QAaHpvxRElfJSxYffUNaJoPPzUeqBaq0jZXcYFEMZK88lmQfZd9ZT/H
heTMnq/uZ+542qeOSpF6GO3EnODo82U+DE8mZNuI3vwr2iOYHTNwhzUJyELwpVyuMHb4gapQoUvG
EGKpbCjhhL7D7ArdjJZojeaW8Ye21+mloncAnr/tEH5PB1TA/beqH4+MhY22PZP+R5M7YKu0qc7x
gPyVKAUHi/G3pUW06ofJF8QrT581MAeR47BhUPx3/AmRoxT7kT0r88D1E1HBkvNlPFGbaqhNXqQq
kfr+vuJ7FR5jZSS1jwt+rOA7dxDpjcYPz617GQsleI9hwwqSzIr6uXkFovm5HLTX+3sv+hpHYJCq
262xq+NDw54MU0qR9teEUSV4mXVGmvFSfm8Fejq0WHNVPKdO0bHGabvkURBHPYzbCI+6XlpvpQdm
rdiNBxHi/aaN/Mau6OgJ3nOjo0kJnkD8gNe2UBnNxr/OqOJVH8KGo2MYO8aaGiRWMhFj5UyMZYWw
m9n5xqjJdNkRq81lfTaHYvwMm4/wSej17snuSaJIw+1D+Om43sgDU7a7p1iIg/pAC4ZugFs7qYKx
mtriHCeekBfct8RVPobQK30NkJA9gI05Ky2kQA8zH03vEu066CJ4afvmHSTWmsWDX0P6cc9g1hrJ
x+ewho/edl32EjkQLTjdb0eW6MKg76XKt1U8IpsXlKKaJuFQfBDu/R804cO8aKI17eiM+x+SxEbc
GjIXs+HPL+qkFjM7J6Kz3el2hJG+hWoj+J8zkR2Tk99FJvFEww7OzCXJsnTew9GeNJj9oI2wxXPW
Dz/xaMIGY+JvOVGpy7jTHSSgdeH3tfjEOOCWkuMI6MsPkikfHPVsaijY/4iMD8E/Rc/tITpcEOAP
E37Mmv9FQ/PX1f+sXTDsTeiRR4C2NaA6/m0iy6hJqDVugGOJ61cpUWvvkeh4x2JTW67RpOQ15o2Q
HELsSxCRytBol3sFn/O3ImQ9wC48pTYZnyfrvuDHGliJab2oF04YYCfBILbwVJdW/glEYG0xS+lK
WfP/e31kISe1Igjf3L9ZCEcmxLrYPNqvfifk6Vwrav2ZSh7fy9rvlTkfg+0gIDxddLExTepE8SgP
p1LTMzbhRPmuzPEhhOhfF/Y8QPEiG8pTjY2HwLbY4+PUKw6/5JqTq64ajE7EUfLHpMKTZsFiwpK1
TmUu8JaN91nZENGhqD45GDNCykpM4SHLWXxtmZeflETC6ZoyqPOZ/K7XZaERo2oB/HQ1TyxAA4Ls
YiVBNfv93QwqLOkL3iAHJ8TUVLtbuYRIrVThTVTElawb4fw3vlLUHSCqJ0MqXnPhkXLji5Fi6hK8
JR0SX6OpKcyo6w+YZ1O9nEgGcpGLhujhX7/cACG2KWCf3zeUos2Dd37G5+rUaUVUsPYt0cUHOxeL
oeFFLuuvO6kgtvFT9KLT3DlZzzEkgtQDOj8N3zD1SiHOCcxvQUfm80QOWktZaGreVD8Njcy+SKY0
Qmj2JIIrSns8XYWHBV3yqAWbKI7svhnEJXJ8flF0bQ6bIRI/F4iLsao1jmMlMqhDD2cOuwSI7C2w
9OHixbkwwsMj/zyfZAYkuLvc3qf5kmlLxNuBoXnWigK4eLNqPVffkpA6RelP19n96BPXNkBq3g0B
v1eStHjee1yRxPcuDOM1Do3z6Bqou38Kq/mCQJRg7V5etEvUiAMLsooy5hYVy8sM9dCyPFuQuBia
R2wBKf6/RDXQ3X9TMYkKJgIF1NkldTTh3PEoS1Tr8hTjqMg1ir5A57OK3IMKJjHeo2k59CPBjEDc
ol/tOJi0wiWRJT+rFkJNqleRUGLH5strdiW/BAQq0hVIuyf5PvdpPMLBh5mANNn1P/7hWA+kkhD2
aTy5Nmhm/qy1lSwFK6GkW7Y5ApwUZwS+vjPlSIIFUUHKx0P2GVHJ4qTqSKBciIIC0oGqvKq54zVQ
U4+5kgkMkdePubBoj0OLGHGbZAfdI9ionkyb/5NjR4uAxqAx5qaofmN/gF2DGRQlnOJEakAL9+FA
k2qhZDKLTzav0Y8J1cu1XAFMIbnHI6q3mXlklbgSP6/Wdfq5VHT76OU/8/j2QKn0ty8oydyBdS/U
uyVrN7x9SQPF1FPrjR4vhM9u73m/hypKWWM4aerJQcs1z/Vy9WeBVfNhpagVp5quwhVGZfyB1j+c
ntHHH54SWfMxGNv/vtF5dLtDNIom/P3TShbBHb0lh38kHdL78zip55PcvWW1nPIRpWII2m0SrL+N
cbe7h/lP1dotH4B8/n7BhMEWJobIZv/oxn4G3sJ1vjz5OQTgAmRhOcc0qf5kFnPuXtyMwJpg01mq
BcHqNCode//urO7GNCv1KVt3Tk71cfJ1IfyOgl6YuK2e6cnGsglfLD8LENDkD0yFe2285gqjedqZ
Z8sz8u4KO1D5fTUW1g8+OHrry3edAXhTIFgflc1KrrrpY4Bk0djy56ZTTEhF2v5htQFDlXRnOkiq
zYjoEdTY38DGfkgsyNHevNNZHoOmmSFRproXtRpqxSszK+6inNZuTIebcYActlTa4emIOJgl167f
ndtviuHSMeLo3pxMgTNl7HpP+OF6uVJ1M47be11fE90gQXAHNrFrZGuG4uqthdZSuOnOvE4FC5+l
+Cp9Ho7nYFrzw8IHfEsDzelpnJZpmCXoALQnWsbjsTax9nvllEP8cSE24qKQaFG3EkCyUYKW7BgV
ulkjs8g5O/8v/reCMSeyTnWnQ02qZQ8/1g81PsectlCi312QB/vuzVHytyslg2JBIzLdYo2SaiNB
ArvjHZ62/pSydiuPT0Uf37Dwx7ZMy/gqvg/G/f7OD+cXIdSfWDL0WrcOIK1DuQJTj5BfH07CHPe0
ArmNYVeTJZ4TsUzq29tscYw81saE3DMsF4wlZEWrhB3IDDDDyZOmEQ0d/SjtrhUbxWuGuED89GD1
EQ4HUyf7/kuDmVMyJW2Mzn/CBC94c/hOp6zRlJCwCOJSuZ7r4fPmOMdpcq0jVimyhBlu2aPOGtF2
UH3hcqK3gE8yCVAlAAl9yT53pe9EAnlh26hwDu7YnuiFa4GJqZhp1xq191hV7oC3+XSXrjot2n7C
5w9PVaQhjDZL3dY29VkXCd95DhcPbyZFfG7HceqDsvLqjtD3iPPaZwdOh4hKargeW+eGsEy1u2Uk
ib8LD1vF05hYuGoHy3wqPq0zDA+TZbeWUabywjJTpNJjilS0joWkQlm6JH9crEbjwq48CBRj0i7R
9MfPSQzc6/u5w8Mc99tqGSUtqtZVYafTWHFQL1a+rNxm0fEcIx+XanbvfOt1o4/zQsC3D1t57u5W
/5l8u0VZHH2h2kRdbakqrdIubT4De8rMKiXmRsZSrf/+98djQ5IXm43pBoZ2LjkJKeiB1sS/89XT
Lrn8EJfnePnnqpFiucno50IBTwuAUn/QS0G9QmeJvpwZ8ocCJ9Rqj3WmS0hbH+U7mgqNXBGar74a
D13PPHF88x/xLX+9JyLLy8fOJf4YXHXnOM061Kou7XQyXQFyyXohbv0pf/U8vsVm5a8rSqO7y9XG
l1Jpp66qJ4T5dpgyPXi8JAWkp818jTrzyjCkKjpnV53H115iyyar72v0ZLlAT7nl2N5mRNay4h2n
n9Dq95FXtwos07IApm8GSJb0ezeRaREYhUv4MncbMpZgGgTyTI/cQVx6otyv43DvdfARYPF8Fuao
voqGyQuCwIwGIG2SbIiWl+E6Le4MbTEQ9f53kBJdt8YuE4EkcgIdZgwRUBI0yW8+8R6wUaLxyusa
NjAX1KPCJ8v1/VDZJRFBlAgMIwK2IDajGNkgFXGO8v1/WruBpqnxIOGDCkVUN5ZTMiXg6tmRpbFi
975ng5VsjMXTDj1hH5ViaE/5zif68DJTm8u/bEg1yu43N3NVtceVRCc+Ud2LZKp3p3MkV+lDj0tP
GZUM2bxq5RawG0fXpyyU+ckJm8bmJsw3bFzoZd3qfmMcpn+7v3H0Cm9p0jbGH5l3uoS8nyirnM3z
1CcNokB7iEWd1GYXmSexs9juIde4q6Mv4aYcrhd6F4Z2/0zpJGJPqePwkv0xWdnX6HlymKVYxfcE
fB7safV3I6uG6nsrq3mp70j+62I9QFYEvPeAiKcTp1dGgiGJe8QmUDHHqHg1CY7i7BCAROlwVwxc
ugrzDbKGbHK7l70ueiRrY1t7t79vVGI2OJU+ZV9q5w3qmZOGU6RCwSGzzzi/LRqPzwwm9XVx901w
XMIK/KVxd6IOmD+1Lq1AkVd/vQOiWY+ogFp4MBCG1vlzF0pNBArQAyfVXq6OS6BPxFZtLXCWamfZ
yxXp4e1UZv11rDt54x2ffdwPwty9dt49plGzF1yo/uqMv+3UkUMU2N100FQJNDstd+6yXceHdZLg
E/1yzSQzr5ocFTPYnWvDYzU1rdhhFpV4ijWQwzvMAOnoLys2gyTsvIcMQACGycVkfxi20543OWcp
faANcsuopSifYno0OEiJJfqtirHY/Thojbk3DbCCWop2IBFUSvQTzTCoudbHcm7tHtpbRLiks+9e
I3btYSnrieGp81R4XtfxGzq45YEFyDKD0U1dFxYdrOHH6R4Apf0lwv+qF/+UKJScw3tXqfQx75IL
K9s9S/nHs7XKnrQyw1spROV2ahahQVhDhI+kzJz128WYtb8nMCgBlwW9avJR1yvMdScHfHaCn521
O7on5bAU2aakTgciZvUiy69WYYSnQZAKxEJ2Pt1YY0KPe8zVtCXesTx1uROSP6b4SjDsVXZIQyHt
BoxoWaiqGLeaeaF7cNiuiwPyrxMraz5WUvYYyJkXornmr2vfENLZFtujiRPssEVSLqylgTzCcTdM
Q/LLAv9hqNNvrEC6iO3nYJlrUFmoMW6A7Jh1y3iGsS3f42eoOYz1OLNqnlYvDV2zJ81au0oP5p3B
l8amMJx/oemcCvaYF1JbklnwvNTT3VhVfvVsvlnNA8OzEMfe4W1NIwOnMDTZS9NKEEARVy1yFNhd
+JG5WuP/5jLxwR9w15FmHKjzwTtwymAfqjsKv6ql5Sun+y88XFExI6F6xzzbZLEAXjgtXdRwoIDv
veDm0f+TnIp4TdRJ89FNX08E2eQ2EfDAzD4PUkzMDeAi/1uljO6qjwL57NBWsiZWOrU81OUyuLhh
SJfFtiwtnrqX2wvHM3pOS5wpvgH42pV94jTCSaW3k6h3n7xskgaIU6QkG5y+9t9/7oCaFhu40Utz
zXCPigtdsZwM+TT9tTRfrsOjuztLIsAJyr+F0Dt5YEL3I9njC5iPKC4XZYSU+KVlLUTGD4mhmmhq
QRLsUJw3sBCTAJcuMan/Rm/zlKk3IivUdG8ePRyouj8WqiHzDCgGdyWtawBJv5Y05xUdGif1/38L
puYfc66UbzGDWL9dPIEo79kEKeCnn/OpdRsAr1oZV1WIctxsU5H9HB9hkmuAbYYV+zRon5UfT37b
k6EvrILoO4EUHUMC1XDlEqd4IMwXSCV4m7WD6x9zMA3NaBQebgK68x0j7UfpH+RBxkIWKmlnh9c+
3VVDu3lv3x3cYbrLmC/bOVKmkHcZnvEaHxg/UvxUFlop6uZtumfLyc/UCEexzMqU2Ljs/BFoKwPt
/33DQCpJGBw++vBo5EeS/Tqt3LHfDo7C33rr/aKGvfFH2/ynlZqhKnX5RdoEYBYpBFd05idOWBYD
XeoiEEX5VbdI8zAvJfvytZ9TNxngAk4LIvdZnwJ93AGl8EI11VaqlnfftgWuF01pu54m2kiy1RDu
CPsasbYs1Nm2xndZzpqkZTGq2zuXEvTKBlbtCC8kJg59TE27Frz1Uq68U27d15P9c0Aw97oqNZ36
m9PN214/OiE+sOx2XEBKuGR2+Kwoiycuvgi30guJhPBz+pjb3zpTYNoxrEEtDM4SIHOfhcULOoXf
TkpE5tf7xvdiOoULw3WSzguJpZfR0hrPZGWJUOXwhi8sQVynx4JTfV1z85og73gj0iXm+3pBWKoI
2fdf1fg4BgQFw7mndtmuHO6Ck9VUa+vXxSr5JNPRWF5LfaiuUSXfjrPT3zhvtZrymkMA21xrBhky
be0q+ewEOnu7rv9E85bEbvcmVv/cLNxZajcyOo7vkjDaH85zxPy0Z3yrrVag5Mm/JJGYbnrlSsbo
armTs5hpqOveYZMRMel8+cbCppjaA5joffxtqD87qioFLutXXvYSPWLXRhp+OPfYbSzuJjCbFOed
SOqqnOnqQOL3qzJgECQpidWuN3Nxq0Cc7ehNuoKOMKgRSWCICHSHAl9o55r9RAMvHSn2jmhN5HCQ
u6gHufN0wLjbxhO+LsG28/jmYbWkQcikf12sYXH8hv2OF8LBBQERp/InojRvBKkor/fFnZvA+ir5
5npk8IVwO0r/H6ygJy7kqHCoG7wlAKggciL53HaJ+jfnnjR/rsA3p9TYTkYSZQR5mYmsTBPzITIS
JBZ3qFVivSMeoeJa2q4gRPvUUg1z/8fDjTrIYhy6X9LJSv4he9/L7ORgTPSCuoQlfMEv1ORgDawo
FXp4Jec04xM5b4mqL0Ua5CJvNKmCm1NMEmhW1NGrE/hiZwD8bciPNo4OHn2vW7iAFf6hzh0NSmPd
PukwqBs3CJ0CCXQ82tKZNx5IOv419ub0w/lGGFXmqqqLrmIKg/rdjnVpnzoVPcCfopop9LpF96rj
nY22HNktTymZo3J45lrZyhzRQgwcSnCLfYVi8aYiUcVv505EcEpd7NUHGYTy7C25L3u4pFc6EAYV
FborZB1RI8Ym66NfQGeMwDXmMPaFAo5PcHJEV9ZOs6WFcbslxbEvcyBICEZEr6OFuv9zhtkGnhpy
6ul64ozzimYCwYa56F9iAqZ0LzPlCLRh1/a5/QwX378gM4iJTahga8bIEvP1O1Lz0ZBnIw81g4A1
21hH7LKhj08TOytW+fV38EjLhJyBYXNbJoKrHZDJSerFaWovFJW0qiYpMDVL5S4UJEADytnO/3CJ
RxieSSaJb3sC+AgqrSQUJu66aZhQAfHL1ECep05k+/53UO/P8V0l2aySHsxwUHu/jdcAW7ml244h
Hokab0xuIPrCGsFu+JhImUlcs7HDFVgswVoKiqVlApajAiuLFTwNyt8/9JhIj9rjYnJjt7uv+0bi
ArHuxfx9vETvjCAEJIVo7hnM5A9YDgJ9w8xB+PELa+GKgx0DBfFyUsvCeXFnC8a8oAidSbwZXlib
ht5EU63jd28LvnuL038InklwnJMU2ef/nMRHqmtK0xW/nigx8f1UaPtyW9Zd2q9EjnaW/uwJ75Xz
jjJqUmm3I2cSY/n5Ykoncfi0kM7yp5ZokBsgJovtfmJJHxjg92V7ybKicyTsKPV7/TaIMMU4M5J6
QHBTVCFuxQGI32Tn4FtngLKSS18f8I+aK+j1IberG5jlRA6vqiKP1TjETQK78TD3O6UPuCBV/37R
chU5283IdKu7ODIwXHwVvwtJTfsyQUs9RV30JfThOMVv+JVLwMDZZo3WH9TV3uar5TdJyBkCDYts
F8ktrxA879eT0ZdYMYFpHjb2cGo47qU217+t/LTZhbb1q3i9yxltG+0z4IiCf83S9xCceuo/cWTR
KJ65DcNH/CrJjr6X6AWjnHI0uuM/nwQW6SJetxdq063R4sSURyXrg0QzV9rKA6XLs2zN3EFIZWNO
2tEAahyQ9p0LWyZoSQ15/MO8AVmVW5+/O9fygM7dBlZFnr6fJvRuGgcPeshLH0p/SI3UaieClx63
RWGJvGDfwnAPnvkc7MTLjtFeBD1/OoOnk2vqDbgR684ov4IO8OLxpFJ9YneGibLrA940Dh4fRBtS
TvwyJGtVm48mnwtxM0jOtsz5xE8EvwEmk75SlMrHhgPz+RwYEm2qlCzvZJDK3RX0IfggJ+GRq7rB
dKnB8HXI0KNMdo1LG/pkIEzfeAfWfGP5HbtSDqZz4CLnxyBqzIDigEyYg00K4GlrbyIQa1lslfrz
cdVLjKDeodCBImkoVBwzO1FCX9BK+pogWRqmqfgEAZUu1GRU+tBeqN1TTThKb5+1HDCOy2G8Ggsn
DmnzMn+j0+k64zT4Ce2SCe4ML+r3yhgqvSyfOBq+yAY4DYgwEXJVcxOKc9RkD+xtgzGWSt3OlMvz
MIl2htqF3Au/r+jdTXv8+0N0S8JMyVA1M8SVfLvrKJu6B5gK+VCD6BtLUD2awEeEmHQmIAs0RWQt
q/3oTi/RYAb390hBUWBbzTrZc2LeeubG9yEuSygygdtcxaNZciThT5zfyqb3a2bHTrG2+8Q6LsOE
POcPIlrrHfcz6jL7VqyxW+3qVObncjv1AURyQEAziE4w0tJVPckoRWXR+bmYa63tioQZcOdceq8J
Z/0Y/o5L0BfaWGuxsSkXFq2LI12+K/BxkKQTBJo5Ykiv4b3p/Ets5N2vZsH8aqXkxfihclb0cDwt
x5cdCmXq/kE4CHi9YrwktagtQWA168GQPKgXmhNA53XCgSVLtBmHvU/lXcakGwWQ/DIU5M5Ng0Lp
WYiGTsnk7ECDGqRmOgpsEbhiy4/eOAdPuoODxs5NcA3a5GrJKorlSd0oOFrPqIdT0stmldV3qItt
9QfxEpbwpPzUzLN/EfvdUTbOmzxYFa2+xv4cUKUQwduKYonYzVgG1VxvlLqvgB2nROXHWdGmAFON
cPRCO++ad6aThL7/bw58ragVba8TewEsaqf1/C5DISLdYEoor9BUvgk27EzNUTChNnMnMGXZ6Rme
9x1eiRlsFBkWbsj3F9nUShZ0ENHE3xJkiiLfCgEBatjzTW7KTj94+DP7n21xNkzVb9DqGMQEYK1D
U64qW2RoUgOGC5POu2pcoQbQCzZF8jKX0raX9Nycj8qqH7xqHGTM+gYZSnAY7cX2LQNq5pzhM5S5
O6CHzlePKBCgZripT37GusrfQqKSsKx685EFM2zJs19A+cXnHFUbsCCCe3YM36VhXi6IjBg/v359
J+LhE6c02vrov0x2ZXE6M7DFgDEGXHBd7JAhS/LopNj+qloRl2EHokx0shtPB5qmWe4CSnSFHfFK
QJ2qughD0+2BsM9dTwfea62SGQSD9wRJAAIWRi8Sj1CiUUOMzsU021DvUG1q5FoT5TF4TlPFPlA8
e42rdKvwlRLBJc0ySqIVr296Saaq1sUEWXGTZLbIIARMSG0CUoBZyamiJ/+lxLcJ8NgStW8u+jqO
FvgkbQLzh5IGlGiNlDIjBsn0MFvysbpwrKyOzubCRFCuzt0Nbblifrb9z4vDLAuULyMRZXUprrO2
2WIOKk4XRCgOZDG8mT2xiwV+t7wJxore4nICtbdRc4Qc6DIOFwMVZ5oV4nxBzOyAJub5DcdBS/hs
LeA4LWbNxDXyVvE3KHSqR/okHUbioKyQ5LlqMAC5RGlVrKw6V9MzCKDVGjY1tgReXujTL8hoMubT
RyL6vE/e/kHz/aLgBp92naiOgQXYsYFyQGEAHvzpu2uXl6dkSpI+p7Wn28UswxQ9HmUdcP1CZMws
8KxN/T276tCuQY2m1qKFaMCJr4MtPj6gbEuJE4hrzC9I9aRaCg79Egxk9BiH44QrOKgsrie5JgIY
X4KZU8mwo8xkpCZdCkxQAdhB+30/6K1cxj6tMGjaG7s3gDYe1stW0FIr6uXiErjIab6rI4OnJZEN
0Eml0a7DUkDHbFX3VWcFrjusz/CBRGJNF5fJmlepdGRXf+eJYKXtzsNpgRQfhHaF04/a7RWvh0Fa
cSxJqSFbh1GGDrdRuB+1Z7yneStbGTWOxJm16UijqHecs3+xDFsXIxLX3RyPgj0o445s87DP2tgO
n0cr1dKoP8kgS6iJM00wKdPo0+ty1PkBiilgNdD3khMMiOf+t4su1FDQm/opo7ZCzT7xza+cyL6M
G2dWiADI8h/9bihC1G/bc+SMD/ue71oFB/lBmHK1Cts63dJK/fnRbyTw/WEj0c0hTsdzIKo62ILl
4Ncl+lkADpJApTCAmcL8M5krJ0B9uEhbNz2GDtgblT9PFYdxsgyay7c0Jw8v5Lt6FDZF8diVgrvO
lXlcMXupPt4jR5VExKgH6zqwC+v6J/3UxVP2PCo7HAJSOwK7DDYsjGfxfoCaS9lRIG9UG02ee1SQ
aFne4h8mSzsI1pR3Ar4yT5kgZLFeKfrDJJiMTy26Vu8AX8IPEqsH8kcHfeoXiVG4on745/ZrEqr/
oSpdBXY05wCf8IKs1pwf/59l9/Fj0eDWE+th+pAvHNGesuTfIehL1/9pwCfjy39oIHBWU506hXXg
OyRuthoIecRTAHFxrCqnHNdsb7u3YaonqGJ8Rb9721z7lgSla7ktcQS/Sk38ZpQKpyLvssBOiPY1
EAlgXcb5Rp7xbJtxA6mTs80RlUsh3MEi0mgTnsrIGFn3RKydJ2xHA0sdVYiI9ySpOx7aW7o/WAw3
7+0i12PYR6DLBlFYYlZNfKAaKrt7HVoOMJkFLDEI3yu7j+K72oNmzYbKjcqVHNwX6In8WcbRrebT
GOVRObEmkMc21N3p6SBsFoUSEsHvkQ8K9xTdXE7ciCAcP3zuz99AspFDQpU/zOAJKwCBYz55UEfz
Ck63EV9pjKMG7on8nqY/ISIpBnVJrdAHOl/MANhlV7rTMYzroAmzeNEL1AhPlrXFGDNTEfmYwis4
eB+QpDQVKwGBQfCV0s3g9Dcf/WBCPyoB35U1Hv2So5fI06e/eYyN5cvtKsH6kFGN/kDnm+EltMTr
3B6nNmQt+f3mnRY+XUdAXiEOIa0iwIOy9kh79LJAq/PpW+nibVN7bQDzk8dRz/sFHLL/A6OZCF7Z
EL+18TqPWmWUo7fo2qnozHnxVqtqSFIp8oGYLOg7Mg1nFACVKIzxZW6+kJMtFVbzBlMSPJuyaBYX
PJZDAini9iBTS8xZbjjQQApQV3NXDOWFWR6nlRS0npjoTS68XWqmTOXgEXd9SZ0D299bKQ0JYtC6
lSqiciQl52jB4rVTCb+MmnOl5VcMc36/SUR1O0wjIYKev37dW8+Mf/O3rjoLLDDbwL5jDC3HMOvv
QwdTM6mJE8eTUkEeJ5qLH+I/+/C5ifth2pmaAPe8adF0XRv78AlnJgKYsCTxrL03VSVEPr2jXfN+
NBbC8oSRmUWqu9Warue7j9ugJnsTuIvgWK3JZiM9m3mPJ19Y4OFK7f7CyUux+Jj8p1cyAz5fw7zV
gAaoUBQs+1bmVjydd87/ql82k0Y+eF4Q+LiU/zGLdZX9owzskMGKxOA/UqWVj51kO+PUy8gXpwlt
RMCcSqvhTEj7L1fRUkGBxFvTPOgLfGZ4MPSOeNLbvVx2s6n3EBttG4zire5azTvkXf9ZpoLWdlLn
y180QHJrkUQPBJGyOSCqh8N/Ulxm3WzLOvyNwRnjIEhJR8BcKTfR3VkiVf/wts8YTtzOrPQ0U49R
UBPcrTCQnwWtwqZNauW+JXeqbaYqxmGHmrHTgcP7Kusrntr1ztsx34q19+sGcseu0CC8T12rE8Mm
llUto2RiMYN7VezW/CSGSH8f6o8t5UOYECG4+UEDaHwYXLqcBW5XILbjqKgcZ1U230/8vYpDXdwB
DG/KdfJu+3KxOEUCg0ad9GEZJybWZWJyPiWsoUg2duIQl1Gou7YQtzDEsmwfpe4jNFqVHL2nX1GQ
ZdKoPmXlWrv8AJUFNFATWCNirCTPznEvo8k9ifOBtFWcntftTIsvHeI7hEJCh16i6cPFpx2JEes8
ff0GGboA4dJl/teUBbia36KYv2yW0DxaqNoP1eAMhHYVMvKxxGF2EQW3oAirs1nh2Mu1e2JlhYqX
6QeVXvUADRYd323aekjteAZ4TqyVhomAPDc+x42IZnYBx/gePjNpqyAOJOzjjP3fk7GMvT0JqVp4
HYB5waQ+OLRIiEDZCZhwkE61hild4simm5yRefCKOJmHMYIjCJ8u8alIiPdvKEMG/1hHSn/ls6kL
FXImcDv7C7y38L1uJpXfBEt3/O/CzfxOhGQnEow0nB+f6kbLJTGfDdnm+Q8fZRui4GOavR4pAuQn
R05s1AGRS06nsu7sN+2OLZKkTSXSUAYZ1TiQKaaJy1AvLwQbxgGMEWbBto+Ruvy+DliGwDhZWy5m
NmiPH32vXuDQdJhmaLkOrSNFOdJXHUHtUEYFkqeF7S2S8Dyzy8KM3zhLv2cUtQVmrDycG1D5dW6R
VG6T95miQHg3D+1W0gyyvcztPlOU9B0YGDtitwlGI94BxDD9fguqAbeYsleKB82vEs/xornxqKo9
TVw7fcxcaqj0BN/VZF9Lf8rQmblpUlQC6iacz9bgNjJ1ehwC/WyZTmijWe+LnjhIsviZjI8N4aI2
+JR4IeTmZKlktogKLPezMnsO38Kb5aB44HrOtyI9BcZsqDbpUc+jUoLi0LSsstRsDs+oM7OSLyCB
lDoiKWGiJ3nQ7DWWLxpJcx7E3FuJeqjI2pGJmw66NJKZ2W45Pznbt3WqvJvUOtyaPEYmYWD+o3Nb
XVobqmKaxBV5KoGmaGltGwyt7DKFXTt0vfjVrNOB14Uc7Bj4vWskb5GSO0PojhWiKRenU5Ej6E3+
32OQAzC8Q0AP+XGUTmDF25XIPZAvnYd8YDyMdy0VPH0UbicFE0oDvcAhYB09P5+k1hQFsFqAmZbH
S8G8D9JmdKqFlrczUE/76gmoMt+BaMLnEjzkOhiTHH6G7V2V3PreyfGcypGwsDjCkS456DyzN0Nu
Ti0hOH4rG/0NZLjZ5mXtwm640DCAuB0/wt4b3q471031Bi9GfW+uu6U+Mkpk40HXadAkQN3TKaVa
kcUn/+RTCD1PT/Jk31qtNuUXnai1N0ZRmuBTgHyt1GeC6f+Q572E2wnXApXK/i246cxuorI16F/H
zgvoH3DA6qfzvGxWoHG77Hn5Uo8xvc56QPb/uO7Gf7Kbb5rYYevAKNBZGWtAab2ZpT51A7Aycy6v
DS9k5lpRqvkpuWvOWGi7LG4rgE4dlrqJD85hNL8TmaXO8DSXc1JiS9eYgzcummU8rqZQo9glIJuo
J0Ucz0D8t2UmD4BDhye5JcPgHL+MRaJEniVYIUkalbqmSsLbqH613GxvcVKWMfxGyYV7c1PaPUcM
DDPvhAwLxw3juiHcSgyq+lNJSPxPxlIL8tJTmG9HWYUdghVVTwt3jsZf743cGftewAv3bGrIfoCz
T05YazWeIluJOWkgXL86TZ0UAkGnjS+dCYd9j5i1JTSpU3MAVm26mZZBAdI92dVSyBmZHUbaGYFL
h5GVaQbKUrH2uGvxMwvGISLZdy+CVEEIj2salVVcla7SBmTyTU4PaPPrz4Wk7DG2dTbJ70r5e6Fw
YxSuFpgr+1w/ScKpydzbXXCOkDN2u9i97VQnBpe4ZHMYCGf6x6AVFrreP56ODSFgKAA4ViMmUZCC
EmvhNjvJxMs089hv5ly82fj/RMVSedu7pIdADKKhWX5sKtqrbhEEiAsZ88cIajNAtK4mgWQUvb+z
ZU+B1/Ap/2EmIYr+NjpJUyFZRv4tnHq4F0iR/0ASLNDA/rRetI0iU4tght1ZU8xfDyi6Xx7wcDFE
qja1zQRehsG+b61CKq5tgYE+ZTZu8fpqCOgtS3eeP1fyF6C1VD8TeWVEr5wWaRzVMhcxXL1tj7PU
zEO/llMOasC+Q2rttQaVMO9Q/0a68cGfWcxAJ9SF+lLScXgs5bOpyLEw6p+HiDOmWxQMZPJAVWvw
ILhFiQXEIsZChDPwL+bg3LR+YJw+VErhisDNt5BXSQDRLIYJ/OTsnbg9Ee2TJoJKLmqjOjHCsSiI
XxiBWH91PFJAE0pzhaJT2d8VT5Rsy6CbhqaTIUE3LecH2oKPmBkePpT9HbhjB1xUwIHf91l7w52g
a3WPnUjQQSLGEOCXcXc718xPW3egvTXWWXW8BvuVRXdOTy1JZJNokYHrnvi+F3GUn0DS7aAkzzIu
GPMpyiEx2W42R99H9hc+f3nnoYGnUt0TRiB/BLCHnIB1AD1lnCVEA7PO/anZM61r+/PJalmQEcaE
UKByeNHKAhdgqlT0GPOkl1p0gyTkP1nI5r0CFSIo0nlS7he8ZQYqRNScp/eue0LcBFUreLoFClX8
6uH/oHcTKkO/JVLuvIpt9fwA3o6vjbKQJMEs3+cb9zLBu0Z2iZGZ3rxrtmL1F2+Fgt/hI73h5xw5
w977TVCEz1V3ugJeVBydC3/SeaDkxQ2+GpHGzE2hQ96rOzQhWr6MRG2ObJlrvvOD0U15k8jawLkX
7Fu4JUfGy7APgrAYliMVL8/ENW1xq0oRLfvoCanXthAa3eg3rRCIZ7GBfCbf5rxksjR9OeblYRkF
ttB+aiov1ajBW/WRJ5ORyfODi3TRdM1+iHk+C9K+xOJxrseDWsQ71jXvhYycaRfBSycVGZJPsBOC
Yd15pmsFAZlAqglFgAwUO8y8qoDMSF1kuAHM+2hVuuTTJyL1C/SLHh7NKTsHnTglOg9fE7stT1jZ
eONiHzHQxTcL05/H0Hwy5/hFWN7yeurGhr0V0iuVAuQE3f9uAtNmI5pbr2/yh3jRH6fDWBF1X1W3
1EJrSBs+wIf1/V4AalmfESqK5J/gjr8ao7hRTzNB0qkWs4xruO0ukGgk2qAm9XG3d6GBgU9Vhb6u
YTyAcwpbe32xC61yoVUBn7OPdlH18lDdFKd4JYEXIuIALFlAfIJmZWaH9HjRifIX2HB1T7ejHnER
PAkDGGAvIjAfMI4Q8ibbT74hxltmDjd0J1K+bLVsftHT+lWenK/tfjHdQtFhNyEECDlO/nqlcitg
ZtdxK4wK4Hywx+0l3jKit7gCkR9ajGQEnqql6ILH+KOvB4Z9bCMpYL/fiGbJvdE4O2imXj2wW2SH
eReCqj87arS0Yo1R8/l2VnpMqGYfgopglDbQR1uyKezvD0YgtsLLMiJrownpyeeAYsh07qabtTPL
vpebZapaQ04FTVURz3CjXhfSWnkj9IytAa5ySQZb0JhqmqQMF4FlApQELEU3DSmAokI5aglDuzar
YloUnTs3gGj+tiJt5ERslFi5p4ENq0NwR5CzAb8/fYEjfIsD4kzOPIilyQ9oOF1vH7d6hs85Pqdr
Bga2xHO/IEbzc2uZDyYhKUi1vmSbmzxgEdw0AAoW8qWAqYJkaJtub/Rb/Znf3CTaecS7KahMHYOp
0h2CHwgRISh41IyI4EdQXeTsgBhJmxWPGmD9aV7Sb7sKEOoIMokdbPUFMKnN72pJvwzAkWZQBLwK
0UK3pPZuPFAZIJ2W+7XxcCPMYrdFY0j2YIdxkdvDgrx9fg7FAjF7/NJEbfYkqa54xCj0b5lEc9tB
VOHAmWVlkF6qKCc/Tu+CalkAW4SHmnDbgxOejVv00As10Z5MgpiMlnbvnB3YXQTHv3dRIGsGmAoK
AzHcA5KgIa4Go6W2D62y5myUufIna9NfVaGBWlwdbJfmJUW1834R7NTgpLFu+3fs2Ft8jjgXyvE+
EnKKwLAwHOccqdGoJdxZO4c/g83qtH+oyem/l3AFNQ/ymgJmIYK08bUvVJWxP00lOgXjJezaEMDB
OQKAojXf7E81lJb48ct9JAnTprcIKS7Cu8KfrXfqmurJyPxVATXnpBoztPxrxqA2TxLJHoxETW22
xxUTdSSxJD3+0hX1fElORIXwyxTNjrw8eorTi76Uk49o4SP0jm/2tsfQqbtGLVJ9uGJSEYECFMf7
qTqWfcEfb7bqr0DnVhER7qa49PWZQGpLvvM/VW9wosrT3ovURynKRvO9plrUInusZyfM9cySQ2Ur
y6WvWnzrUbjB9PNX3/EDt/djx5SE7Q5G1BmYhYPlmAffp/e+zM0GTHzER8JLnJfV4ojJ29QCfbBt
nLWpUL5n9f7xL/QV5hjG/qzKKuKQ13m/qTcb5V5I7Sq2/vyxKt/XSnTis1KhnLDwfzKdTt8611Q+
dQNG3oQwM1yPVW5q2S1ehPtwRHHQiLjM3h4LOLpKQVrS+52pWpqUYt0/j6lEdoz4IYhSppR4Ob4P
dd3eBVnINlMAo6BGlN/dmSRN8Nv838Kvaa3XLgSuZxr0Tbm5yxWpVuGhuWwHPMd5uxbHsZyvEINC
90SVHRa9Nf7hyG+YGEq5YMoKx8O1Ftm9N8SV/WiGZCY3WL2w/S9f2Bqd/xt8yGoGKiTVw8kG6mIE
fW4G9dKZC/1i+yvXxIYo0v0BrkTgioFw8pJYzstGec0REjpZYG6Fo3+UOzmunCHS6UcXmZGN8OnJ
ytzyLKREnYYGPc1j5i4z/VW/ko5GPZwtCQHkMEXzIMZqd2lkfvqGxZdccZ3v9qpMx6yWhoa/ZWQl
tNDqTJjWDqAAAiGB97Avbabv5fxf3wy92Y+weypYgqXXBq54Hd6wTPNQxsYtH99MeFAkZqqci2hG
I3Nxg54QyuobfgxUSpR7IVND5MHu0zfhTgTk1j0/R1XSwZwCj99ipsOXk8FF8v5V4RTY6tubFZCD
jjs4kxCfY/Cb9gaDmTSDNmp95K9XuDA765o7Wnzvn0n3PcL4OWb34/sgiVCzs/F49DZ2hyXyp0t0
Nb8GGp93BJ0LlG7NSwcwgJITh//4iytdV4mQFxqxJNaoKiCt1lKlSeDwnxPy2d42xI3621QpDIFV
1O+hXoPK2Ieyyx2gL0hsoyPSnJO8006qWq4vol/6VWPBuZ8VdegVQW4/vgXrIPQwoxYg/dbQiNxP
CDFhgzeGuTI37+1me6xOAojRw8omlc++gr2ft3M986WzAxLgfIyYhiqAEEZAKzNMKE5cva9hzT2e
c4fvPXR0TI2iGSudLqK+BhnpHtflcT25n+b1Sw5s/EUS1QXjjR4MMb59ul8YxzrsUs0vpiGL43MR
k0K4GUq7lKLG7ATl8/d1/qAmUBUPKaYQqB/hiACEb5J3FBGnMZkuchCjVC3ZfqTXril8ML26gX/J
+QsrHXpHS3KM7SFJDPBiupdcilwspZuZn+jgJ2t7blm87kwCV91O8ndliNQidRK2Lzcu1Leh8KHj
ZfXEHJkqRgghgbbxgiGxxkiW0npM1wV2AZs6OQ/wv5VgCIZTWbdePVSxao2wR5n0ALoxO4YQn0m9
eMRlAJ8PS3phZZi8dOzH6rJlRg0rEZ8PTgevR3iDBzBr6PoGWVpjmeVW9ZdNW5lpAHVKwwh3YMGi
eLBEVORKBrslwpn7nYBIMDo1o5w35ZLN25nzKc2khgmDs9Tuvjv9bIuRRwG+Kybx4qjIunDBDGhq
uMVdgoGprsoyblbCShQeRFW+It9o5SXjr6xUnW24a+5Aq9iutT8CCr9nhf1qv9UdfhPL3CDjSVx7
GHdR3S7tnsXfBKbXh9P1NSZOah0mmDlPe2zkldkqbBiiqK1qcONmD2pms7D/ewIPJNeOzx7acEGw
9SkkG2SO1tiw4qEeveHnW4Ct0SKhh/hAPoO9itKEO6mWn37YWQxLUOrJBfYm+/3z5PIhJSar/Zan
2fKP0oRw2yMm/WXAabtwEL2WbewPj56OMxDaovvQUG0nrMbgkI3ab43b0nH5wtQ8tBx+jNlkuupQ
ODYl6RFyjgCUXt6CS0+3Wz6QVH+Ry55nTauxfysxpmYozL8TWwf/QVpGcQ+F2r9q21TWouzwLpbD
rk5PhtNqWYJqQy5IMAfKr1AX9pn+SG86l0w4pObGCpKzBVAkpwncxXjLqEJknc6HkCP0H0RBxOLi
7iHdDN6cDR3GDqd1cprMNMiu/ZHYrg3XjNsc421BZd26ae5+2Z5688LdzZfFWqGql84of9z2Jglx
BvlRVNI64f7JtwEJf8clyIPRA1lNTdxxIPKO+v+KDtKu757zjdj6Er69k9tMbpWA0LUMipVxFnCP
xg5gyXm+4KV14HRryWl8ODhA22LuyyTk/0dirkgv6SkcPdD4SlIEr2b9ZEWslBX0KTuhsd7vZlz9
DazT7HKzKJa/QokE2A6DErndCcxI9TeUbVqMdQksJATCsCfXhlmH/rNAuZ/HfaSnQY+7quaCntJs
9jb2LhUpy5j3Z7wG1abCrikqqAOfH5iLe/OlwABN697Q1X1UVlOlb3isLucoKcGK7X8dZ10w0o9y
6QKqGy4RE92FHabkK8Uq3DUDzxO//FpLrSfV/PSc8OrsvTTxFVchmxaNG+RBEW4dle2w22K/HAGV
oZmNA4mrvN1P4QHMwxNTqpXKfYaR+uwfQMuICaRxWMVEezE+TsL4v0WgmVwsutCCOKKA6ipNZR2T
bo/8ANam6Gj54AErcMBvuCpXI9cFYukLdNeTDb/LaWAshy3N/Q/hA/TDQZUDM+vTyDgCuNOlzvGW
hvL89bzh9H7vwx0tsr2nHvYz+HTiy9dsLLtcs6/U0RFR6KhXhFVKR8zZrmUwmXs5YXUACl6huHpc
gnHfMhCwQ1BKeGcTtVUt7Sceu5rGz478Jc68yzOYizOPCOu2I0OFVcoklmix7bazoK0mHNMTDvz7
LtlhEoHo/AeB8hA8qKHdxEPZsE8J7QrpGhU0NFvd22UhT0BElx5EoY0FllHrSJGlbF6AWkXtfVEc
8dnD81XMd24AcpTmi1LCwNkXf5aOSWywhMl3SATGLopwEDfX3amQFIg8uEZuI/NHtIRcAuoAHZVP
JiN3Cyhkt/d1nW13kWLs1Qj0pYp3AiCBMPuqQ3gRkv11Qq9GxN8o4sd/2jXIOApn2Peobt6lmiF8
BU9bfRvlOVoxL/oz4KUHlYXy3aWkFrTNJWYV4R+bM999L/De9dAZOYvfIAhToLDPXQ0jMw6es0Jv
tNDMH02a2YrxNnvScOe4oqMtpTpcksbWdjlJx5vTO+h34eInSm2fDyKm0CkYEVm84m9zwHvgrf+p
2fxJ+KKEP+fyOm5wrMrC+E+v5qOAM6yQq1DCRz7hJEjz8NaYeNkxN+IvywjlVrkp/hKwOG0qrCN5
SPZi5u9V5REy3ukVrkcqFJU7IdhHBE5DKtgurF0/N2N+VKw/eu7qATvEe3ZUAXVb+vAEaOO8QEAi
VYVGc2plHQBwV6U8u030TOLoUySAMdbx0wqyS3cQ5p5n3n4Q7NxzRBmxbLy9vQ3LTi/xsQ8MpIAl
QCrEmdgAkY5VvrTp+xQRuTqTjsKJ17bdIWV3h54s8s1Kk7MOLmqU+Th2QhRAbOSQwloKAVfzVAyG
zZ9rTCpSB6qS/k0b0V54SfhVjBie2izFMnPv8bkfc34Yj4B9aSrDfRJMAvmMXBYxP2akzMA9QurN
sMdzf+iDsdUzIWglkck/AHE/82XSjMVJPJalDuryZkpEMSoqr1F0aaTK3FZ9GvPG87Gh6iPMX9b5
067edQdMdWxtXphpCEoyG/uz2KYn4xX8OgPV3AOr+6oaKTEXP5G4qP4qWrxSR2Jo07lX3KqeVi+G
fC1p6OGY8Y+64N54gsSijZ1Z60xfm44nXc6NcQIiLMHDTkK3yxf5qQhfFsh6vtkUwJUU2BDnS1lo
u+noLRYYRsCIGV3Gqn3yMxwb0Mqp32ufqbmMIJDSGenMuM3as36lduTOeKS6spq1BOZT3f5Fe5KP
NBNeoEl5tSrR7AeQX+Di15n2Fq4TvL0P+bfcJk1wHB/uf1B9I8JKruHT8eM3zlAT1cJPSPyrxPt2
cVziXwBcAlm77UKolSABVFKBQX2Dd7RwMb5MYOoMv6wyl5LaG+EEmbCAvSls2eORpCdxGHsqEyNo
gUTAt0Xs6AnHH9+7y8GRAchFIr8rrjeqy/rekxhjNaJSljTE9gBsUQptDt1XamVLTur4fGlJTfcp
anWt7rnuKCN+qTTwTIuAwsumjgLvLN7Rd2O6fktWnir/xWZDA6IEW+ZsMxVSNhPsoI7HGmqODZ8d
34LA9W9WfEx9EvTyc6MR2AtI2r8TM1o3233PmGNKag7szqjCeg6QfOIgszfKkIXmrYMpfpOfzw8U
aoz2KDIO7FaCl1N+pANWdEjf9N2KFRiAoCziqsOGx5W35C/yiVh0pfheZiRi/1WVZHNxjz/PPrBk
+sFEtIDveTVtI0lmFsMUOvVelZl+MOjQUyftVVdqfyUPz5wuKjT0ijTYnRRQYuPqgeAr399rWly9
RBbpIM7r9Ab7TEZWV1kJMXx2xYJFYQhXN5JQpN9dq/nb8zV8ZVHag4xCadvQv7GnkAUMYiOpznC+
HjN8AG2sYlZ0lBhUp8o3+YPDSf2MykdGYJlY0WmQfgMEiACP7kbsJbjp3bgLvtSNpke5f0fU/MkT
51dAkkzvD+3tN/3fEjuU/YpvzlqN+9MR5Ogw4yreyDfbqFXUnjJD/m8/hmXwVe8+JMOgEOO4J6dM
JxsSdaCt5TFqko6JaAe6a5PoiSIX8yzN8IkBeuYHxpdkBcUA/JCJYSVRC+iphrTqeczRDnVQp9xM
hmRsztZiV4e7vraLy1Fh9AI0Su7ywNY/m5/uFHFyQTi9t3VmGfVJE4XQENC5EHiBwrWVsIFVH6Hu
IIUcYAx6nEuXduZL15nb1WLGWvnw778wJlAD+5uFyiPH/FlpSMjXQm0IjW/Hm9TU+dIunIID9u+i
dkl85JmLFz7+W9w6yXnPs1xOA+R9zE6qpA5uiBFVxn0oO+FEwfr21sFhMOEVRg8vpw/q6LtQw+yy
1YDmBqIvt5KPkOGzbcyAmfkcsRt0VC+icroOtuBNC6y6qJC0IaemRVcyJ1O2hKLYR0idBwv6qv5K
VPIDwmvgyaqULQg9yRxjkoRGAnlYNN9pbZvSmu8ZNojfic0fpIAiLVcdERRq7Sr1uDB+LHHSo71f
uTsXpFQh4YFqWRRXtPl2s9cmPP4EJ9pZNXCjDNAHMjQldMXa6HN0GUrm/+fcRWhbbOb9xcFC2fzv
74mzpDBn2XuMHSIw5vGB7q2ZRYboCAyEhZI8oHjTBwWYvDKOp6qTHYflkRUWVt46DIg3mCl7F/7I
yL8rCsq3BGeWw6oblwk04P1wavepNO7KYrNLGeVHbkQqlorV9bhxca9ve4qQAWGsyb4dOsAWv5gI
7rUK+dJV3bOnzAAb8Z39PIMpxElomWJSD+xyBK7G4qEizw4YE/2OxyYKGQM8UIEQi644Psv8yQ7v
1owSDGYUaqdIMMaEqbRNLjSBg0ZOBWMOCI6sVEDr8RjF+WDkl+pFu3wVNK4dZ3ksBp7k6l0AWcZM
ObgCfcXrDUJjYGNb/lhX3yKsWc3hpgIKrI1SANzBghI8FYf2NZQiad5CsgbRlsnN42np+m5v5VlG
YPMqim24bDBxbxcmMyWJ7zARq276s8dy6fBj2YWZ3ERLkbBBn/qdzsl6IMwrcejIv8RXRvVcjLKA
hCD4n4g0h5De3nmwDzIVBGnDDfIKuEMPuG1SjHe8OYjUZ9lfcOZvqQLEh+QjbjI2OxscOgoIJqTm
A9QtJUAzAt35BW+IlJynp+dbuM4Jc/td8K0GTwZYs7TFOEAGi3CbGIv/sR5kHfjbEA5gFanrvnfQ
7QL0jHqPuro0WdRKIiyyCbftF1YDmCDt2/4dKyoLeDWSZcuufTu6XiJYNTlMTE2TLCm0B/grp8iH
h9D+aX1z1vFJJaxryC9sH39SZiNOWbRxnY0pppMyFCk9vczAWLZRdw2630ubzqKyPydxUFWEwhAB
PrtVokcpeMbZCpnoocG/gTaiszwrF0mOuWXKWlG2RDkN/9cze3SH5Fdand4qPXQCRocFd2YZtbFX
1YKX7PsBZHIfqO70i0VtYpzoPKiboi4EXzdlsD3TGpydQBUcJC/y6Nm/dAqUCxzuDV+2qx9cbDkj
+2nE5XJI9eYL8P8RdFO1CHqwn9K1DXgfX3qIfH7yfa3hmvlJhCFDEXOPNCOG7Sf8hmjWQHzXTBJW
8iyp16qAM1V6ABF5CnI+FvzJvSnoc8DqUkPhRVgx6VSabxFRHEIbiy+7E7skG5BOGB/9aQWoYRmd
OB+dsXMBlZP3nikqmYyrhDkeAPkumwF3reh9T5sxir+SNPvLdzkh86nLIzSW4/dsalAKF5fbY5hc
lQllPmfvrRGsIFiKNCF5fmCHuX75zfWoxj6sCfrBVip9jhzneEWkhrnqpgOaWwls6PhCFO9vGTMe
Z1aEUjzrQgQo2FhZvaMjwjn8JXv9HD0cf9aUhoQIvFsiN0y5iY2c2L5lJP2/OuxI1JMbocoDH3C6
+G8AOuGsT4kXswGfF7mZcsKcKFhn3k7nTi8OQyEf3KDfo5gq9YznyQE2yXgJBCNQsexa8Iskhd69
VumIyZUcGYO5YL370eTg6mxwJEqYE9SCGMsy/lMGBrwT+Y9rHD3r6KDuvOY5wh60JjyLgxjHp+3t
UGl7Copv4uAPF3O8OfpVDQbtiAC+uYIg4RKP4DufKQpGIYJjk7q1G2lIbn0nGsLoU3c4B+V+ILLF
nx4hICye0eLMsUaZJRb+k5AHhAgNktj4tvNBW12vFsM21rfXedFo9jN+0jJx/7Mka6ERbZ7uertl
2Z/kaTyTmFKCT2AVhjqZXUsKPv9DHE5wL/nPvQn+TLcYwUOr7404tqkkiphOb2H+IqucYSmzJT+w
CE7LL1WtsVMByjyyC9skPI/R0iJWobRmPFYwau1QpcT/MMHM515kcP9khItWJwkNFDtqIcaRBvZt
H0Xq16kQCUWECOAuCE1BqgivkXPlHBpB7POdDfHFAwiRquqxdaMNgkmCguUkrxM1W3IwLLsZlF/7
2CrpeHhFtYEuaapcjIGCxJlw1SAverR9Jg0NTIVG9GCpB7fcuWDiysYWpSgGIgcsGHzWD6UxpvA9
flO2mkbVvl2Y/B8v6WNqmge5HTQYW45mFZrcdZ5LUNXqt2+Jms6F68uAGROVYBLASgAat0E7Seq9
kcknqEgxca/iEJZd4/3jnBcwPzZWYaiNn8CsIS5uY9fu9RQ/5f3q25CvPiFvsBhVjUsIWgmV5Zw0
zGHyk3aV4BkDvGimEsKQLn5Aw5IbvEJXs22MdWUJKvuAKoNCvZxvbeDDIRiinxAhkw0pIvC65gua
J1JLyvlXUU7w1odQL6M37oDsDFX9nesgbUiNDL4TYxNedQJTizCMr4iir7WfemLY9cDCisnuPORB
OdEiHc+Si+ABSUaGJrfaVkrvvjReC/3oqUN+PqNH+pFbMuVQhelacnLwYuPaZuf2tRpgQDy4DK4d
5WIk0Z6P/RpI2huNC2oYFAMc9gckwpxNf1KA/IzurHqAruqcjDhVIxzfqhEB14vjwZQ/juhjlcY/
/xTUHW71TQRZmZ3u2wp1yhp9pJBkyjUD1jqnEC+7sE0hdLOOvaFKZoyFFJzhwm5IEuAY4SNtN0Hu
FUGhaljtWXohhl8KyEUaBeEk+BRWg0qjjKqTYwe70m7tAWqxMiBSCpfuI4oTf1K34jZJjj/CC1zW
I7ij+7zMk/qbgsY/iiMJawl+KV5SZmfkPZC9A/NT2Jw4vbuS4zcN2tvr/vVfDgx48VRAcsQiARmt
ZOt0Fj4axjXUKbcdaQEmo43bPom0SnjzRBpPGR/Q447xUv4L50gaJa43uGOa9yBCidtvQuMg9bP+
bowxM9hNx8kBDU0VOk/1AWPjyjF9Tx1zc89b/oQ7082NSrqk9JsMg2gxAjVhQ2+o+TL/DZfShlD1
fMpmMZPdZjFsYjYMckB1RMDKm0qihqz4cNYS1s3OHFNqqpkM+6UUjSjjcaeLhU90BYSGI0jL863S
y/WTD4Pysz2sF5AZm6ujozixPPn+yfTlIVeWzxYt2dPWbA0GEB5lrpWrhaL7qx5DSf8eB7RkIzRL
vdeQ3vDLI7Hbi/TSIv4fCffRe/KJfDWWTfgvjF//i5RB0w8O7/Y+kfwEn/PH+dHu8UZJyHws3Gla
3mqg2esaeWCUKLGKyfm4atX0evpE3mxUs7JrMbmffbZ+ov49gR7hczzWXsHsQlPpumJeUtrNSBPL
M2mCQpcpfAHU1R1XTfvS7ubQM/3Y91aK/a+BHXAHMXkVegP2Ix8JSmLPFKIhNaTB5vdI8YCegJo2
KptjsF1TtNNV8z/kSmq8TJOE/yHF1kIFlrwyjLj5aOjKtJINa149ObeCCx0stLMgEOclCLv3Ji4Z
ap3lOimg/aFnaSPnpvxUkbNKQQ+Y3YDKw5Jf75gFH6qbHjPv5Mpkr1A5V6kfdGuBtJhSzvEmww0y
nrUsR4VZ2klV6WZp2CovegS/Q/ipDU4BSmCy3Vt2+pi4SHXf1cjiuzPmCqaQTbs1VW54xPnIQl3l
2eUOn82ctmDnKDys6NbE3501e6Y2ycs+C8KBLcdWkcxnB9L5mwGJ3+Ou57j1ukbEIkG+wMfjJL6Q
Pv7x0n+U3W8Av7AKC7gYmLUIqgt/YN6IoDK+bVV3XjEnG8rRUtOH27fpOpf5ht+bFaQOLtz3dj9b
JFoY4/t5zLZJeUd+gybOkxfl7cjIHohhBi4eD+4clsJkYGynWmWOBs9yE07/iDSBk7NIKdLxVVZ+
UO6dMd8u189Us0u4lE3BYHRORM2C8KvNTydgv36g4S+h2+Dtuez7OCEzoiVoh5515eZq3sXb4b27
yJMyQKKnUZT6mCYD1YI1u09JgFW9c6nFQcG3R0khdE+YPlhOfw347ZvQbOGF8gqdMWENUXQ5CrEQ
nEJjlcsUxHfuHBSj7hiFeHCBxdz7/zXjH5bm50wk6lZjOqg9dUiyihemVKwnuDtj+3iV4PA8T67f
Aspf0zlyGWy8pw8Ny+yjRbQQ1CdXgD4nTxbe61FGh0zoC6+clQ15sqxV3f7em7t1rHe3J3ducnNo
DwI5rgbQTQVSyeq8Bksd1ga3px+0pHy8v1yitIf60z1AfstTzs1AsQTOdz/Tp1RF21v9+Bh5+8iW
u1YNECybrsegXgBD7b9mm062PX+JA2b5WRtEFKatMLNLrsyCZzynjeXMlGjhAiPWWMDVsd+ln3uw
WfvFMen2iONN73tBAhLZhvc1lElXr9Fgadl9Dj3jbFb8mPLlqkUW8Pc7qrU5L4tMB6uelcpVXc1y
z/u1FVtEFWXTptqCczwqrxAcMAXYN5zSQhdrRiWGnsy+ZAcd0Y2vcQ1KSeTXK6qpA6tCrj3TR0BK
LtdOAUUyRGuhOoCE9lc+uZBZpHKn+1afdQRkmi6anKFdTQxAelSzaeRnDFMwMPG8PyPIGSjqAD+Z
aMbrzQTCfsPw9bq2ue/oS9JBwGUkVlNXd126B+bNLGfvMl5UJSfccE6OX0VHvE0FMuvTIUzypYhW
mITthfHVJj9W6jgstuJrI/eK4U7UGuuvsnQO3kvVxvHdfd0cS1pjjA6qXPjzkDnsXYk/t7lpjygW
QNiJSKoBottntyQVyhbaP8A2qPA5GImGlVSJj9ih9nuswlAirDBTE7ZlygdtkTpt9Q07vmzkbVP5
vHNhewKsxXViZwJ6+8pyX/j24tBRLUj+ioEHLD3RAxkLwhH2qcH+Wr8fjVfYwEkCXdMIr3ji+zvO
YArXGIMw220Vcwr+steCx3vCZPCv2fxI1llvysI9VLh/Gq5pzjSUPkngbSGrnsuaobiya1Przrbv
pJ33dMCOgHm/I7A1unvgIhfTK/gThqITNnRDkZwYUwzdUaUjmJwC9q2RpFZyhiAF24lfT+fSkQET
eBuafpewA3IiUy6n9BZ56At8y445IuKHLI+mjsmqy7m8zBJCWCuDfGBzdkRRhQNBMFeJjJRYe5eO
h/NH7VKrJnghJoAatvQSO7nW5KNdo+g8568eZpCG7yYMsHSzTPwEtw1zm6ySbo6l4UTA2AEwQwCv
sozvknEsWm183b4oodUwzYNWjGMCn6RmMwEQTKJY21hed8Lu7J8QBdDIQUbYi3ClwsYkT+FO+5+c
ovluvLT45bj5eKRLvpN2WHu3vINGwout9h+gps78ICQ3ziT+jUfGXUpB8VoK++JoGMeg4WB1sacQ
8RzSIjhLedLqxPXepicK/WI40FWYphaCgyjkqs8sGuRe+r6E6mF7XzqA/Gr+CxhfuArWpCNJsWfG
fs+nAwnUG4sZzp3vvc8NzR5niKi+ZrKeJ1Hh8o0ArPzDMIIb3ZXPHTCPOerNlgoQPdK+cab4yy0A
Mlb6ZN/Afa7csSiIFrhZHTTQyguefcw8+iqLSOTsCCP9yCuo9ktg5kzze952fOaOEjgVwVYVvewE
XgnGUEU3elzjiz7h0oc4Pw+vMW4ofJUCoeXumaE3kcNvoPZpNdG59NtY/mw3BNyg4gxNNZjrXXM4
2oS3Vf/P98q7cLX+DtK+cvkJUlzk5QkDiG5ZrXvbEw3gaBNrjo8EiuapHLKrTpmx9KHpjgmLrbA2
UwF2ja6oSNApZzoOnZNksh9q0/oLcWaFVJc8ML3Kj8C9CigO+U/e6bE4DDcYOYWBjX3rf+v3gwLP
lmNME6Zdaje53qCOvk9HgnXJynp3yk/Xi6/QSlfKvFUM40+c/BuAP1EUUmgSOpBB/+S47slUEbM+
VqVB9IkjjVQ3osWHV18tAWrhX42lZ8So9R1DgdAYX7441adsMEPhwysYGhEY4Ulzc8M23vWxvYfg
OQl0QeiYmHG3LaPULCu3n/q0JqRhMmwFZNzUvXV/qJerVuQQM6QmwIsk/w01C5jY1rwPrOKVpZfh
h0LP0S+238oCTwOds+zfipl3UoHlHeAjJdmrUkLeGyLO25JP00sQ7JD28Lq0rCmSs02JgAsyhB0P
wyzzVK/RsuyXgWzt+0pbRGOhXtCjss//FlPMBejGkEJVG19KCsd4PFpEVoagSvK1Q5Py9fT2afgK
6wXkBaYpU7FeEVDFlPx9py/pNQ7lVqelNa2o5GX5aXyLwt77tgg96g38VGiG7E0LJ5DpieTgIRQJ
IPhWsRY1OtbDRBqyAQ4PHX/yWQr7CiZLUZWJHzDRs0kymtSz+/w1j5ZKMzbcmcoPO1YNp3sDoThw
NkDcXs3/YPKIrvKMx58Lq1IFwdMBaBUZbj53LvqLGwERVEgQ//BahJRsM33m40BI5zw0zc0g1PZy
GVEfCnaWhdlIsmIQA/G3e1rLlxlUmR30JOH9A2zt05d1kLahLKFlaiWnfcxPJ5v9tutOy/vKH90+
vsJZGc72VwUnsjYkT7SIlVIUc8SIssIxiyvR+P/q78bMWXHtBJlScmUG4UEWJRvquR7F0vgEOy0S
65di6F+DoKZgXX1fDTKUbDpahk68m5hA0KdWMHPlrVwdVo1l5icxtXlaXbBS2J1ydc9GMPLEMVdY
GrYsnrtyNMfBDE2++NCSh2zMMlBCRNT2XpYF2J72pVhxJED+6W5+W1xc3K1eWoPQmteTL+qtXKL5
IGCUoIplU1xaDi2eCZUKUSa3NkaR93n9p2Mjx1t75Z8oNtt1EBxkhrDK3d/jhITadrzB1EK4zz/M
ElSSE7Fvx8og0Rnn7ztLmIOSKy0kvnhZLN1HeD5ehtXmX4UVjSdH+49NW23P4HwRwQ3BDWFgtW8e
wHOCjoJ5tknHqjqwQ5xfkqrDdCAFCy0GOchVanohiK2zr9tDsMa6Pzesm9eD/dw5wu2l8+x2vWme
6mYS97wDZpeOY22QL2JDtH4LZL0o668ZxxylG5Kzzr4kT5I08ueB1QBqxel1cCuqEn8xOyqjjvWK
Hq2ZFKepLphP49loz8OjyolzDVyB4CmUu7wuQ+P9cK8wwBUxt+7k1ynrCJedTUSEIVGFtdk14tEC
Zj+0h9e346BW1AOeHeFOFU5/qHwCb5PJKsP79zHyfqD2pEVLd9sLh3HT5omPm6vzAgMXSYt5CEEF
FkQlfMlILsKoaMxEQNIJsVjL/p7bXu5aReAEBySADh4YrKmeY628Tj8VjNXOuJg+c9gCQ9KEx4MQ
dhMYyItlyKb6cNvCG4jfGtOJ1uQjf+Qu34iaRjjqTMmIMFxOjKbR1I10mBKHy8KTEMM0hILFIm2Z
R6jcBJeUJ5SFYASPW0q/63ZawvOrfp4tv26B9etqOyB8wX8x8cKsQtaeCf08DxuidBcFGF7Wg+Jn
VJ4nhQEH5m6BAxr/4Xu1WIKn7PMKsUy7kwQGKK1GQx1/g6/yIiHMLxlPaO+2DzHja1nc9aSWUjmm
YMh3M+sOle921hBKQCRshtpA4LOsYA+oMti7FWB/7GqQQkX2Y/S22AieC48oHR5aT53LBjW13XN3
GXwrbUdtCRx/xM7nYkN1IeiqjMhDtzHvQk90Avaf/4sTlgoAJw38uq/eXp3K7bz7tY5llrEmOp82
cL4DYFcjrK69chnWY/vbrMyRp3NlbQX9KUXlqhK5kRjysIHikq5FUtszm7lN6SBInMiiO4wamKOn
JD1fq55bgawhd3PL2Qt32a84IpGBS+odgEjDk6uNrVmthaTpBhH2++Z2LV0aADuYKnOnKCHB50Ko
GarVr41VSwGdXoS6mCd3T+OQ+GG+6dGSIqGwgCytB59uj0hmBBS0MqAClnM8HQXGCS0cPgWr8FIv
IH/hdrFN0Acu2+XkijIyY7GL/YL3xO4qYtphxSa+dYyleQUw+4neR3Kb3kPpcpdOXJF0NydCoogc
yHw5o+SYfRSLNrlsDaYqM0BfLIbftsdNn0KOyD8unfKWruB0XV6YpuockIv66scrzmQCfwhu9FQJ
kmq+eLHNtZyia1+Xr2i2ec5UX+NwaHObdoqw8Cj82IeulTZcn2UK+2/CYYb3+RW1YeMSI0cWhKmn
OrgwZmOD1pMQlyd4+uGMTH4sSU7vq7fyzwLSwV37wLwkWmdH6dQnYg4uqA8MUtRQpmQyqAnl3vyw
VTSps2KehyG31nO92Bz7UISQPyslbSc0wyw9dJoFC7IBYy72vLEQ7twAEH9mkhfvGeDtT/BgfXJ8
42oCPybor2jHpDGgPSK8tKPhZSGgvUySpa6aVD30iMlpBIrSNnj5bilrYTYRMnx6DfpVHl2Xkjel
U8m6MezYvaZUY9Q9MvhmXo3j5xe8gZPVHE420LXw79tHlwAXwjt1j105XSS1Ve9YCIBWdZVQaKQb
+Cs5Kqe1fJhsTnq3O1I8rTttl+LA75o/vsBnL0dBoPM1fQiGpDy4aLTHLFeR7lB5Ea8qYGbFfCW3
beBmJrbBZy48dNrfkY/se7h2WUIZ8qVvcuTx0F/SVU8xKAG2kmH4Xi5mAyYkM6lBgUu6tiYcydhj
J5CfIc3qUXEjNRm7rYM/j09u/5oAkQtyqRrEO/crzU9aHtslABBqF2ICoJq9YWjeEhoBUoQOHSXk
BSnNKJ6o9rnIeYPx9OZ9rW+lu+BEQUEgDjXToe6OTbOVAmDdFgh8wE7lWJU5eP71B1G+6Qkpj7D5
3kQt2e7FU6kVVaVDgVheQv59/c97nxPgNiK7VW3B3IXepAZrrDwlCrmlvOPuaPlTnoX/pZgk4qUd
4ZmJopyGkDoNWcwOUUXiJVJMeTbie7ftz/g2ma78RWQGom+TjGzLd1/JB+DeCa8hong94pFUsBxE
6hA31bWapDYfWheam48qtknq2qc14Pth4R+LfQX9ty+EuV7okI9FgS/KTK82AZ9U3XSN8R9i9mhP
bp1WcFYIcTO4pqH26GjY4eGRuvk+FYPCq6ZiW/HZdXhFML2gDw0m+0OoIK5A6geGNBZ/ZbGf7/je
nwL+Ol4k/RU1uN1XD4qY/aD6WCvHuncvlknDr7CtP4tb7IzLBDQ8O3xWAe4DlugfeM/bIx1lAp3K
g6T22T5mMVIpoyhdlAadlox/NGnOD3C+SHPCHNLAjU7ohKwrOpqCY0J5xsD6dIOFh3Rh8qMyklfi
kr0GtbBAEN1bRlsTju9GyprdAJ8nZdfeu9MZsfo7N1yoJGpYyu9TX2Z6ds6LNufr5IkUcw4thToF
TcTBlGKUK2hOWD/OQl8f9S+yZ050oe/KGjw3x6xFsLL1i2zbItHjS3hPsPBTzBN4LGnFLEoewpxz
8qvoI8rT25Xx1CyAUReIPKYiWoMTfx9f/SxztId4Fc3OEu63fPvUZ1ogdJteQ1VQwWEMxr84J3xw
vZq4Qx980lsbOXi762qeMRmQXwYlGp603Jg7N9pS83bEgqqXS2iLck9V368vyjYoH54xpLN29HNy
RhkxTOK8Xo2Ve3/1ekXk3VNsCEU3GStkf4u3Fu9pJJsDV5K0744P8Lsz7C7qN5JqcuOumwunnz7S
37EOv6SVHJGnJc9JMxErp2tsPDUHul6X/Q916PoHLvSazkM3jTa66TEIaQVCsd/ZE1pQeMp7kC66
94tLqG1xozfG7DkFKCmDTVc3TUa306YlU9ovMkPsWYhTe9eC1J8dR1MMAtbrSThkSzB+Y6b69hax
1aT7Q9vlm8zzRCBpyQcmcd+dp7JO+6W8X3T2yAS/geDiInqfkMhmGuT808FLkQI77SvQO+kfGfn/
r0XFazSwh6SB9+jQMo/JHaMtqE+ynpa7hM7PQhBxeUCwv9xvmaA8EZLL+RcoOZVONXXdciLuKE/b
bCZ6UvIPl1xfoBAsR9jcchgihtku2oV8Gn1vP/z5EU/F7Vg7t40+R0EtXWM9UokTW+wwWbYApgAU
r+p7TuRB89eMixrRWBLBRI91fBB+kLdeP54f9QBGxzFn43WCEqjF5B9QtE8BGJjb9a0o3fwna6zR
fI6k+WAEvaUqVDFsSBo9uM85tYtYlWyr7ZA5Dj3Z5rjB4sh26RBXCgMfgv09iR+W9t9NuEoYEvCX
I/0fWoC7EDuwU3E/3/tNls5dVtwVgzijkwY+0EGBa6v4/x8XSTXa5+DOK7jyt62cSsfzmfKpn7il
54FJXRAviWWL5fhOHIad7mUalFVhIwusckrrn3m9YahCTGlztzLq9WkxD3aRVH79+KS7bA6fQT0a
2X8+60ACPS8qX3Loq9yzGONo6iq9+m5daSko9LaX4Oe2d/kOU2QH39PDhqNMC62NoPqj2/X+5Mkj
ZC/wsESN7CwQIiGYkMG6cs1vQ+p6gINQiI8mTDj4ZvTt/OZoG4G6IXnZN/HIyjKz7vLfbHvnp1Ca
RXewbEjzAD9aO6klb0QSYKOxrSeL5QtG8TowyFdgW2pRTdXPI3SRLs/6XWMkQg2oON9iJYnIMXGH
iV3bI9Q6SgGrIXI4Ph4LW52qiFgnPwodDrxMIGxRJHrUENBIj1XkPeGSbH7doFht1v/yn8z080TN
/AhI1wNNPQ8Goo3PgvF0KMHnNNzd5AmCP5bgQd51fjpNitthvytPAKpU3sH0GRt0nr6QwhJeyxPQ
l90r+d/qZ9nyIgvHfPEIr4ZSJkoLqlmhEzbhUZdZBnyhPK5Tv31dl7XHxpR/4kKUpcvhYxK7i1hq
SCAPDghKGpnE1/iBn6BDvNIhUOfnVwBBmKzS1M4z3PiT4q8slkjJdpBMifgN9C8msFW0xHWQYM0q
AhFQkO7uWadBrdAe29Y3/tsx0EkFSIAtjCG6pNV/j7ZHPBo70wjYTaia33jAEzJpMkiT3WpuGONY
v74FIJqbfvJNUnTV7oYZ5j0xS4uSXNBsct5XJmNr7N0qvuYwFBcbsoPFr6QyUAy/np2AtsUWUb8F
zFzigepJ5DZG9AxlDDqLoY9AAe4ejNvd0SYF3722GVhy+yeQ6khCs2FNJCPdvuPRlJa47LQ8xQZu
e1wHaMpPOjhdQ/CBi52dPBXVY+Zd+GNT+nGz3xzeTZsqOSh0Tq9MXObPewFKt+8f3XrzTuVyCmFH
YqeWLHM6U9Dj2dK8PP3d00LFOWTSEWTmzuHxPWzCIOrq4ASRpeNzGh49bF06m4aUl4sOHSmebm4b
vpaT2qSHfd1qEtg5oPbIhqTdSeEEf1hqm0QA073hAtxME6Y9JRHoIZSVA9gYsF0sbB+LKTO4h3j1
oUY64wdprJclUWxyaTdbF5mLpy7zvg+kwPqNXgy9dkr9zFf8v7cikAAK5o/4b7wiKU/roe/s2ImI
ehMejcF59fIKfgqqVEa6AFLZwv8m8Bp4iBgucIMrq/zqG7hZ0YWiaBYNaXNDMzXuV21+qzeKwUrS
iI0dswpmJ1dgYYtBKqXYjXySfnOEOw176MbS5Ny/kRridXNsBaaB6fhYAeQIfon5m0xcUuY0dCMT
C0L9tSgQRa1SUXul8aHTZ9+z9KNM3hf/wEL3DUVkD0j/C9WvByf/maD5HuVwa5l03QU6RxnXn5vO
wzXMrIvLECyIDiri1yTEbt/X0FJEFXkALweHJFZyql0ipYRuOaSbP3cQZWW02q8F7hrzoI6ZSmi7
gLOIV3kUq7zcbOQH07xoK3QsKdozEXFKS8wAx0sSxRUTQcjjlUwB74PagjF4FsTp1iWDWwkSuhXx
pSZwYW8YTW83LvQx3fCMawJ/R934IHEF6vOsmNtbmtko8Vm288aeqBpI8eyc3Q7Pqb/QolpZjyPj
rXzqRCb6Zy6Y1gYBAm0k4kgkIQPsq3OquoUE00lbct+nAHcNvr7nq+wGdRubZtO8sUgQjghAeIoS
+N2Xoe14q+7nDjmx9L8cQgw/wIw6H8lOg1+jlrFmiqqsraqb3fsUNSfVP95zd990BgcO1pYECnWY
ESkg/sNMvfMsoSKIAgJeJuFfa3kG9xvlB0ksIXtRgvIkuCT07ReeLsv+kqK6gkJQxJzysocxGu0d
lWj2ryBkfAFM2B5azR2G1zQxIfw+tmLJSIUDJryIJeNofHzqmMXSwPQ9jh83z3IaTU9BIl9YiDxS
sii0Jrs8cVQCGmxgHiw+Gc7cHcfQdjoUGNkSoUqrIKo0tkAtyl7qbSs004avkQ82YXhiBLZOlW+3
soxBIpWDFcq9IFnut1PvxVqPONeayGuKHv9L6VOewPGgNikP8ZTsF2mHcdfl+9ckHimYzQwQeREk
i3g//QFn4ZAimT3Mj8I7XPtFB94N306NhbuDhrNypnjUN7M6Ec0otRCqmDzIzG0RoaNajArfaJQj
3nhkSn+nbCklcGnbjwJDEBmy1idASrSonaL6onuliMzMjdjqOcl1OCcahQEDU7yQTUJ4ndVEjU52
T4s2mMm0chaaa0QBPspxWIXRUMTFIBExWz23YeM/wnE9RzOsGxuIbrkFPImNCI0fxDUvX7X6S/gi
F0HM9fsGE9sKhg+sVl+PPzV7w/06EXzbLdVUiQZSesLOZCjfH1zaX/asoPp9xwGhZJLAFs/i3t7a
UPmUFNUdoF/xi0PkIHWdbKtfS29nn2iTRzY3X0cUhHmeHnHqr+jNzZWvBxG8jAGrwXutb5ZBlMmG
sr+OCMs5GTyNd7F+/qrSa29o4y2SoQfWhyaBGIJsDVMxwdBFKbZVs951MwaypNTcRwYXgfDSvCl8
aeW82wu0toEPcVSjPkltJY5ljnF24fa0Vu9Whn8vGNliyUBp7cLkiDHYK8y1VPGnp8MWraUPr7sH
zMlDaA0X4JStlAhXzI5vhFYaGhZlTc+M9g5qaWfCt5Bv3uUB5ZNgVWm4ulWcmOzU3yzMRLatSiEC
asOyBLMBaBQKtjeIYpJmVcZTTTT+o3b3NccNPWfgIBqwFgFwQoStdoA4V6x+3EPAH80+YUJYJ9QE
RMQ62o75vZTsdqR5iZEwhHUAdRO9wBLcrKLaK7TGZWTnAeOhYmu4y4BLjrkjkkTMnfK3pKoFY0Rg
mcSzZZgPCzMdJ3G07m+Ejq5hxxYMai6akO61mdMb2eGImAcHVWtP8LBuY0upZDcaNCsQvArd3/bf
H5UZ3a5EMyuS9hzXnvYPKPUDz4/Jxjzevp57bWhICXHZS78+vby5FGP7oycIPOMbncfumwn0BDRj
xGkVeDoDehGLqOqjKE/d8dnU0QdvxEzglwZVv+SL9R+ifZyPP5Iter9JBGk0LLzGWIGCIQklwrFe
NKOmJrPfpW8dYEM/9x0Khh2EHet4ZWVHD4qwSBGgigFZ4HAilTcta374kl6LxF8J7hKZ/F3cD/yn
xwfPRqkQr/T+9V+P5Li6XnAAtnl1SibrWndLxa93o4fYwO0h5J1pb6QRU9fhc0hLAq66b++4pXMf
5kjlapqrfNy20vHUhzbBRVkDBo/mSGVDGU7cjxND0fbOH+mK+967WUMGUSbLHsZPyxXHHLsQ3Oec
RxYXglm95P3PLLdBWgYcllJMpz8WUnHz34tpiRtjGjwUJkUkPCFl2ZSHQYhwPfcWEAFXL3Hw5Uq5
TPhn1C5V/nHevx5JsvTuYl7nxi+VJElBil0wejH6PqDkATcfp8FyuPP3OH2ErfGtTFJSYmp6Z25p
fk6RpvHXHUAGGnZe/x9SaqKPMFOlzozp0ffXu/RmI7Ox/gqGRrFo844vug1u6SxvpX7a1a7uPz7/
a9WVxmGwBTQ5ghfS8WhjlWpoNTUCoTJuqR+/27r+u+dzrDV+CdQovPu5p8M9t3T68q5TLvY1Wr+J
IUqVCtcBmls1F97lg5yJWFkflED2sjMCsGrDXe+tVoMrB2lBBF42fJNChrEpKto4gjyrjGQXJ/T4
xkvMdNMpp0XmPqlD5YqNfaQ2nyw6VGxnPCIhwRPC4efNbb+HHlimat3CB4jPP4MN3oH5p+AbH46t
vIAZQipEoXNsxMBSI0uMP8R0I9W3yvVQrBt+XxyZj1ML2ZtGTowpy4dIaC1eJalRCqEp4zctXPLc
+G5q6WNGCNrYMY4hMJKYSFXtWHR62lX/xlLRU/B+unGaTEnKVJpOmWkDYKatTZ7F02H1OuWQSQ65
4gKypmyRiS+3is7CBuxq067dC08LzDfpyEazlg/3fMf4s9GMZh0nmUXlaa1dvDiHdYNL1Oqh2oQr
oeY57f/izGmZLhoWZxLLMKq/gIVBkMCpvPRwbL9tRxzzgAYDXDG8E+g9dosMm8/uG2n+sjtZgCws
qF45HDuWlMYskm21MIuBsVSau9i96wYemNITlO3Uzi8VBQsJuYv+ileO8/wVT6ZL6kLXByAFz9kW
zNJwLSjeqm/QLd8s+TMTgvlkir9BxQT8BP8RP5+Xu8B7od8H0o6aOK3ZIQIxPxFv0AscxfuoPhrW
QOD42GN0vkR700mxJbWZ9xM7GUp1Ft5ECZfV2Gd0xQ26GKG9LrDhicy7/sQKFIUTLzRrmWjEc7ZL
Ycx9fc+1dignnlsXo2ymjnwU507cdOTTdQFv4j6qEhJWaUPSO6h71WPFuun4Dfwwx1ObV9YT1TyN
5P25tp3XE7zGsZlLGakbsEbJ4dHeQO9/PyuBKsKlmnMMfsXC7VF2b8Y3B7NDwTeKjR/92VkPYuaX
hRn3pKkfY+5+vq7+zgSGt7N2+N7FV8n8tGWJ2j9/L8z2EkysX9DnNy7qKoSA9wu5lCrb43CRLzU5
oOi+9q195XvZ9HL43pkwv+qm6dAirpvIGsDwpJe8/eGNb/Xz+MFuRHZ26sP10zWhvGovcohmL/Ni
tLN51XmvUqD0HwNnSKQzmpoEwg9T+WBzBKMlUFUqNLb6DZkvYykmFHe+bvO+Yp0GownXtAF38wG9
kGgpuLQsG8sGFvwFmzFlwCsK1Z9O6AHr3lKyJ8Dt052Xd0CVZGuWgpAutfUtxjmRrPbi4f86oOtj
e6hkTanL4AsB/xKBolj0drxs7c3FYV795jh5mnxbGkAuN5/9/LJO+aBKfhdv93KPAP0g+H0xdicY
OdGquKPm0Yd0S491Py1qB2oxiJjpQdKUfqkpqNiDDMLTuE33NY3ZQWwFWY/cwRujDuA3f1t9osEP
h9xv0LmnG4dlObL0QnAwaYCGsPjlk3aOFugIXkbxU0k3plo/qyGuit37HyAwz37rtAy/r9bIO7jv
VHDyFOFjTHvJWtStFEgED43vHLyh9iHzm0M/ghqR4vgILL4Fhx48S6S60nXzfpEZfSzXJBstFDEB
jSOfS8lmYKRFGBhF4yotNYIFmx7ppnco6jivdKK8LuDwu1fJ3fOcYZw05VKI7aAVIpF50p06QZnk
Hv9RUG6NMgzYyLzL19u+sBpFShgs7UL4nkiUNWt6TjrEkm4J6ryUaY/HhZhqwAP5ism5nDEQQ8vr
2/5y1ozhmNOqjKsfthJOyVK3jxI1ioB3V8FRj8G/rKmsRn5fYaED7dbOtqPjF60Y1AS1o91kdFcu
Vbz0eheMzRIzYQga00cOlwWbGmCF7YyFZTJ9rsQPq68Jc/uuUjRZIT5qdW09vP2Dncy5OiCy6YAZ
I5rP6YHbEbOqgA4GYSfyDH9mO9luDY7c1yqKPpVRy6eW0n5iSWBl7Qb0w4ZJQc1WQv80V/LBV3dS
DdKSCdbT6d7ddBt1mPO8ZwRDkyp9NtlRMrHCnOWkmue0JNfBtdDCHNf8wjH7kPaoyTwf3esc6cNB
qr8OTj/lV4HtbZCFLSgOy+OXyIFvuI8lPZ9HoGdB0YV45GX6wo2/0oHaCYEhwM1o2+dIwfQ9E73M
ZDtikNBwJ3n/NtPZ2dhG7O6cogPKCAnjsDhjWBJbTUT6yBVrfd6NdeodLz7u8fQODuT8zBX+JUsi
O3KYYRs3kUmR2GMaYgTR2ZvRyVM1JMefQBc3X/wLiNyXUE6FpWzjI6JuYM9mASTR2VToHw1s4IOO
qJEcqwaQ0YfINH2fQEPXMW1r2ZB7x7F/ZyisQwyIpFjmqmGOPEsmPxErKLcgT5b9OsyxEmnXEYTX
HOdlvIZ4rtrFZ1oDHnTBbDgu+LsVExAS+SsUsEjX3Gc46+aBbEcTQbpVtmMOG8Jby9mmu7YjbxH2
Ukbimil2utTJAczz1T4k6Qc1jH+xyHrdEhUFd4euFOx7/k0mqcPljaZitS7IP4wVJ8CxwtkYb3pb
WmLTbGshJrmvYlyBMQLGcY8rP9ZTJkdB4wqZNaJDawYE1AmQV4hLuvUWKISeTpVUXb9fJ9AsjNwk
0+ibhQ1rIZdFS+TsuVBw3BfL/dlbfI50xiE4JrMgQh54SVMQZ1XtIk8cPrrAZSU7XlqCAJFRZbu1
y1+LOqTvO6fh64+kRUYa0rKTHBkmR2R/YR3YU0nappKqBUroYkbgDABmiMfnaFZGPwQ2pdzr0jnv
I9NlRa5cFMRfZz3UICTgsdbZbKD2x+RGVo4ZsY3f6fiZ1vPPKHC4VvKbULiCg3ViWgkI/E0hCm/X
N+LMLkGxW3ORNnnqdQMDqxSYVx2Ew8R93YwOZ/oULA586JgSFz0lSrEbJZmbUjrd854pADrsR8vZ
slEjqNsK8YgNVMclrhpgRIjTycoJyUP0M5WvlDQI5F7n5xcI6X4ivOwUqfBiE7iECkTi8EiEC/vd
/BUn3Qu9NwYSlOMMoc0YT16mVBepNplnedR5McdxwdKUDflLhJjdLWPODVdzkPt7JGV+9zrbHLw/
IYG3rLjCO7ZqVGPbfVzWBSDZfA+jM5Y9a9KRZHZMy96C8g0rhuV/Dmq87XS/sK9dpKVJhlEJahvo
lkbmjoTEgpAvPd5w8vEE2TIGpueV5uIxlKJfOaRkYTH/6cG0jtY32aqr2glwchu4UhSiBruJH5UQ
+hRRMvEBt/xiQR5GRdBPNU057SHTUnXCK8Soa7z/cs3vU5oJtYz+AVetAD09zB6HCCZEu1q8+cLN
t64Gb4pElMuB/s6wtjFHbzR5yssoossi3qjc1PtvexYM1hszLCdK5wzuwgSILXSQdGxtcZV/AK0o
yUYEflOw1R8DjJyT/MomMIker2HBhjx/Mzpb9Unboc3BPc0cJ6tFIyyhVwk+xnJnSAJeV5zxccc8
gCS+tE8HqOzt6do9/CJH9OB9xLG/Nj0WLnJLgTbcByci7MCR/h0SOjt/gxpZEOG0h9fw68BgbgFK
0My6WK5DDqEtZoxgkYMw8S8OL0MhCK3VkWAU9OTPU9cLuyu2a305uZLNCEM9/SFQLIC2NhwS91kh
1vQTfGISFUuRbBpUmzf+5kFvq0hj/CygFJzUuwc8Ht0hxvrb4v3ZxPSbflvyufrb3NsZempxDJaF
IL7+fzYUCUVwwHK4jdgd7cjyCYj+YtfzyA5qR3bt5qQzWD2c4D2EmDwwy2CjL19tYQHfLIQMoN8+
aPGH6Y2gQloDUmqr3/KBNMiZgoWGz5lBN5dYrhN8KYmwM9gp3geIdMNQgXsSHyU636nsTRmGBOJn
356F5uMQHQNMoif9x0x8s55o9FmTzmxwlGre3/SzaVGTHbDPJP9UK3HlBxIxJ4qTxcCtVVB1TjTe
zKvjOp0SwRUPYJRbR0R7ZEJuA4AgSEwbuTNWj/UuzcVD9sgnunGMpCEeUzeqIafXEjf9bOrWJXDM
npd40wpwsmiRYiOXP/uXFIgJ0h7wql7eEmBpmSO/mR85HChBxWxLUIewuNP/hUURm0JGbGRhf6W3
ecCg3fXcJ7HSXmDZSSrvad9/HduwSJNyxospiqmqwwrrkROGd4HsN0w2NNqWUO90h3TNYAwsgA/M
anhWzsLMPf9PyAXQMkP2jQngV7Tt87bkfJ1gj1ZtSIZr4gSd+6TZL+32aLtPv6B896b0wy/ZdR0o
79W31j6crRyUzA5sDFsKZBdz8DPzKk43efE5+jkE4Hs26VAu2Ihs/W2U1YsZW+F6bpLZIxJe6mHj
hwr2UbXiwp8EMMJNCr8wcQsF4pNtsk1SYDFJoK3mJzbGCDISw1uWfbLRc4wx9CYYg9F/uxN5YVBi
KTHN2nq/ZixzC9ASEY+CtcPuQJdTpjI4ZAfRA5tHxnvP5e+IDGivUOABQif1tQMYps8lKdbrz9so
1bHQiEHIrWbq60FCWtVacN+B5frOQ2RPg7DJZX8LXobFKk4KQ1psPQ5kKrjT+wlfrucRui12/aTi
/5SfLgtnWbc8MnLzlc2WRW9BL7RnWBFmesivNFg3Az9sKGTOBOS+w6RPVTjDJLF8euhGr9Gt2bcp
59B0DeTVcgzbNmBsBBF7C20UfAAiu95QAkBBPFf9/CbH/PuMM084r8tSCX3qfYry42FfADr7ZTXV
LovNLlbcDMe37eUI03Ci+BkGS077LvHrfDJIWsCUqGDx2NYsgruAXtGDbzkvuqln9Uf8I51rM4WI
DDDEs1kDvoTifRQUFjU8wwb/dCqkvgwLRAx4VyiP/0cTQc7GcKET3sdkm043qgEprhjnj71mOsY7
raT6euoq7ig1+X0/5UKZoGulLByeBo2yi5crGz7/WCQqU8NBk/eZblKc3hoz64HXK6oUe1gvCpqI
4Rjy9nEdeO8BlhObdZKTW6C/fA+2U6uy3ePcXmWxKI+tcAAOlp8H0iF0V8nwEpxALW7PBCWME693
Is9oUWBjExgL6nJ1K6fh0UYgCri9hj/9uaozlqVv1m/LYL/yNzb5TW8hEVp+sU4h4mVd0sX/k5B7
G738mG1UMGaOddh7FCB+6eXwbsQcGJV6SBcVBsmwFAjOXTgpjaSfv+qMYqHv2j/dF0cG1W0Ifss3
uRp+OvPfJVgWBZhT8N/7ctPXhvgLofJ24/RixLwTqROtxAd6BM2LjtKzmW5Y6wIC45UZ7sLHsAE4
dWXTCAIj+1ZuVbP6NA8ozq758Kj1md7vk3lM6UP2AqNGR8ojYNVygTsOARYAZA64gcOTaDOrJ14y
Xz1X3CINEBwKDczgbwF5hqE5QH7LweM71J5lkhs8ulH57/M+X42/c+DwQN2+FJg1M46Q3Xf8MDWL
V4u1OTMm8/V4bqWuv78wSbn87Z0j/sEBBeirGGWXNlr5U9dF2h2i6sTR3OCnstq15FI8nKmoY4jY
RkwZHmjMk0YE2/o+D/5W1LB0kCOdloX77LrBQC+KS3RcY4s9C8A3oMwpMeLafHgNZyjkaEXxLspP
D/WWRLXWP+sDjAwZrLNIfwCslcCfMCOdGP2eq+u57zQuksrssxbq1MXnHWa2Teihuu7vJdzXkPXB
41CUENO/hH010XddfzOLPid1pzles+xbpUOXWCvlwZpsNuxORFcMMR0fiGIfIWexUuXB9acSXIRR
ewVLUHr4v4h/0CUfAuSXB+H2S2eVVKbFRmTs6WWWl5CL0ft7mrnO1zjtZ+UTxyhuKWJIVbDlidjS
Yi+Sso2Uv9zcP4tAIkDoi8v3nWJNYRtCWXI9Qelb9FcvpAtxFydpakkrDkq7ooNuyuX77uYnTEj+
HlYk0HJSskjByLGG7nkBGUi+WTCQK3waDBDkfz7jccPkvdE1HLkvI1LGkLou3QKJCDgQ3nwS68WL
gvHiXLbSDTSAWpyRLUDKy1C6nN5KeB09+NIwp5Cot/j/y9HqxDAreWKonVOH8T7DP/oCC34Z2Zxe
FCPuw1qGzHjRXjHkqSv+3ZwUEmh32TQbxRvyK+9xSGUheOX4ctfxTm9GFebJidmyxocNnOwJwBoH
dpVqnLzW99+7COyoNHC62wuKUoRNrOOrWfAvlVUlgMPCNMds5VVMmatBWcM4I3yJYYlNrCUO9M8h
9MczTv/ea3qwQHTcNQ33xr6xYvLieopuItC6l6+hDAdA5DqPSePqS7nnkevL2N23YentwLelQHDp
NRv0RlZsR3Awe4lCSfcI9nSLovZVcscgKM4/EtRSLb72/vw3leRR2Ix44ap7Nx9eoz5OH+Jkc01T
VfmmYjz/yExRpNMoLrFmsAjrOoqthmsYeOD9l8p/jgcBY/G+uBQfXnXi5usE06TU7+KJrnD3JB3i
pw4QOeqoxxo7yY2BZII+Sg5jKsHN/XIRQW7UW942wMmqaep7M2sZPYcrsg/fRW95OQsbu1X5uW3v
hcjX4qTh46KUyzZ0b89L68scFNwV9sdRT6iiP6RpGhaK6mSFRTSBBwYYXHa8A9ZUbICsC0Rx+aim
SlwGccwoDJUXceOTQ1KnvShHB4SpwIt1DtgnVVWSTqN0d6zYsyjQhqavubaJpG+h+KE/qW1LecsB
h/dmKAafdQD/WrkWFNvyX3RT2OiniK0yjT06BTaZMkk17IFgX1HGYaiPTLQ+5UvATSrK7Ku5+tmi
5t85quqo5gDM8+DZDjFAt+0PxpMeZSkKI/uddZ6bMiDie36xvhRfzVjKJ55wMhM8Bmisl8tXAN6d
VUEtCBXyAywtE9vxKCTR/MDkLxqQ8jfuCdMsmsh1bwT8I6TLybsZFEWjoXuHjmD9FScne4IjsGtz
2tbvbklRVkdWHvf/bLswF/Oa/Ov6kroZuIP7yNyhk+NKWaT/4MD7QO+FDhxWysdv6yNbSB+EB/rH
n7oU9Wf4MKtG/un79EtDHpe73xokBHOGSSr6A71yRYXY7djjTDosWsKcsMsLwJegP8HmO2tIisme
u6wrawa0EOgPcdqTb3NabYF+zsY7OEphe2w1ZE/ITrS/SE9r4Zz6ic+vP6R6mOOiZqTdhvhmvNMs
B3EbuSbKtsfdpn4BBMsoi3Vdgsvbc7yUsD0DztBwAVVjE82ov7HS07OAq8tEfb+o+jvks2uJXbEV
uZKrDf6byvA7tETs2KupvVUKYiaTJ5r/DaOuUmD6VMoSrSLCn0vsh3tU6KzXxNIH+BkqOm4/wWXt
PUIYiezcoCvWc/QllPLcc0SwuwuG71zT7mwT0+VbXii6BtBh0XtvMRbrXIfRqjAVF0hWi6B4B+wP
xkqoxA3XENfrhC2576R8zyVgldA6PBwyvgzOXnYyZ548AjG1WI0AVK1/KgClt0ho6n/lz8Yqs4Rj
qr+HSwPZj3Gs5g7dOrBh4dAT224w066MpSI9ySc1X8GT4HYrD1uuEaW7tzUbg7Qr20oXtl3AodaN
qpFVH6/Je8iml20uXQGFo5d71KTuT2c+C2YGmcY6rwIib8e9rNTLaI560u+3jn+ND9DKKucVbBfS
92srFZTZYSF7FbrtjBXUIt4d0J6PNMoW+aH/OgZ/FiQAPTSl9B51GQ6fcbNu1Yo2jkJvOVAA02cE
JTK0EXvaIRhDX21zEIF/M582Z7RdhkosCFkYb0nF/Fhg46MbO/i0wmtIY6G4MNTZBQyKF8AzdjQC
w4nAoJyCOCBXJwkMlf2Gj68UZbl6P11expanBXv8x8cf+4ATkiitqaVfKkrkA0+oWta8uLjBbeeO
N8HjcUw9aKcgjzRjQf0niE6Vpr4lzIaHrA/kiX5lStGNKYWMouUybUB7RJVpL1S55Btgvixymu/l
bLxhyEy+LYRxavIBYqtrw0aDyFmVk+dk7BbGiqGQqczAkwm39fMuHMWPFcBCRbxiVfa1cM1MN44d
BY4P8J0SP4NjOeCQen4p4gLw4Mv6/u7pxexQr4/l8XK5XxCaK5bw7BkPXo6rOrg+h9xB1zNB8RzE
yYalMFHqpDd7vSmvFfkE9iVIa/RJ3CQd9EqFHdXReP6OMcrQ9oSL3VI689XRibdFtZEuZu0bbyhK
KmX43OtHNDyDE7VqHJTlimwVTLILG29xod4j3xeEcLbUlU6LKrMZHSjavfjC1chX038CK06h7kbR
k00U6qwi6THF2/Dro7aBly1t6i7U3sIRZQQPQJnsbZzwKCJQybEMDwhu19CL8sD0NTrxqGEV/JMO
bgf8+aicinj50CW3Vn+yuJ/rL9ElTOypHw8ZJRBISsou0GiVh2To/hIPKnOa5wePddkgKbeqh87e
Wr18tV6rWA6Iu6jGG49+CGxs6hBbi9JhmWRODaIEZc+HyO+tkdscOCCUhMELTwPnJLsnXZ4t5PF6
i/cRM34KsvAv5ZQkop5QTKKyS9MoFnN0q1WmAXxSlrjMToE5x2jh1NK0n7yfnTpeRmXT2SaCkdWo
OVxr+1f1X3zTf2lEkWbDwDBpRduRtRca9fwpMpXhww/mx7/NJ6EkK3fcTxdgfPbzjv9tijAeXsLx
Egz51tJEYs0EAUWM0cospbeElomBLBdeK0eKXc5c2yPUjXKFQAmKisfEhogNjQHWXIdiJPSdE3HE
5tq1SwfujayBm0diZtnv0BDpu1UbFpdry63JTvDtxvAokuNG1+Z+ptsxs467yzSPCpfZGJAcZ8av
28gBNC9RH4yq23UcUWL5b8bKeNhsjeWyARolihZL6nV7upnHsq1ypbhkrCmLDXP/ci1rS/zgyt+s
+oF061IOVljb2OB6B1kVgZFUFyrfnhfdwhKuZtwkaOvO4X+gqQ58aguJ7fRuqnMFtPuO1DX/xqD9
tE1GhYXTnmE3xNHTw/0v4W14f16854jvFCpykTLPqoKf/j8T2flvWtiwng762AGFyGa6Sa4cQRUg
dItgJKYbej4lpSsmv3brdA1uSaNYscjcTgtcRK1tGbX7TR8IvulsWYn/SKnj7rWIkcLWMX+GoTQ7
AgEI81HHisfNXUgsk9sf7GH9TSpAaFlUPKSUwJd5+RChlEI2LZYZN4J+qjaB3GIpWXoGieMUgCsj
cdlHQD8yyMF505iG9iZNcGWIoGsw+CeYVzAt4Uv4RHvw6ktemvQtBlSg4g5J63Jl2hibKvVd4wUP
iT/rgbeMXsBjWNsKWp3wDnTFjIfDd5+EA14em+0Tl4yM9TDhtiTzCTd88sdhn/37SSxwfuXP/fuF
DsiW1JFY7dW46rGbyVZ4ol16ENqaHcWrxh5rNeqoc/Z4zwpZxyX7b7APMV+bG+HrCP5UEHvWJaFR
I7HtXUJ7lr+UoHax1l8UL5/lePm+9XmWuQlJNP4GZNosXXiCRyi4NAzw0DweFn6u0A6PvhvUqc7T
vjLFwxI7TbuiZ8Mn3xio3Qlaxn+KaxTrrwCf1jATo3AJKBhdMiGCj5qpK1zwX9TGfiEAofLWcImB
NRqwJzuR1wJsFnQKmmTijZlAKXSkdg1zBp1Q/YrQmS1OgQ80du3UWUTi+JuKVUcQH1A7La2KQjwl
tM3CxmqYCvFNbjtavQmv/eUsuX5w232OBQ+/9dCGI0Rdp+HCb/eY/X/vPpYMWDhtlq3OX1I5Ryc/
pwd5V+6qd5RaT5M3zyOobMg7wFfdgo0Wq66bWBO4XFGEijTVFzLxr5PyNMvaucdaGlBEIn9kY+ns
sNGa2QVOpzjy45JL4Za98GOTZAFCLnYNgXocr1P/h1IrBbk6LRL/x+42VchvTsmLw9qhpbTDBCkN
BHDXL0RZgKJ6LCjim6ttW3vvK/WLgBL6T6yg3shB7lj371QlEOBovFKAnh89POCE/GSC0LhQqodH
V3IpFVF0RZA+w7H6s1cA52ytcNWdXGmadHTqP0qrM7t8T/rAfpkU2XpJ79iCsg36mKztLtKPbPih
P/XHum9zJgie+iJYov2DJWVyuQlFty9I24YVoK5E/TeHqGpcNxGu4RoKk9AfvR+1mKGeR26VnI/k
xYp8KRpfLc2j1J3/ltx+BasWhdfv+4bH0sp9W97sGz+K41df3Hs3gxUVxnt1oKceWVyZo749vpPu
QS4ZHA1fwJ88vUyufuZluESZIgHcqEr+5VluobUJa87QPm1NtIbqbG0MZNKdfg1J8oMdycgIhLVs
16baAcNAdOaPeXi1sor2+2yT5dwehYtd2BuRa5DnWWnV68JESk/a2kZMVt9CEmVNC4bS68zy5/9Y
yeObVsDj50iAmPZQEWKksFdpXzzX9EIH7Nf7sxbRc3Ro9Y5ju8D6UXuvTC+82H9vzdnQ0Cr1N+hg
ZhHVLiVNm7POfobNkzbQq0/O4isleaHn9mMsVx0Eeff7RLLhTWOLNxut5muEw3xmQhoxYwa2b0oc
qW36Ir2pn/qFBHehZBSXA+u4Y8tQzFkLCf1bONtSGBqcijJ44dAoLtqSEzHprME1nAP07wNkeHXv
PcG339dREvNZPkoxhXNtLtIp5l0fJvZQAJq+yRvEXDURhOfeAC4xC+EEo1GN1khIJm2QF73PuPX3
ANXDsZLS3fYOlVzjo55IrKcLqgtw3qlqV7NoUPRqzLw/S65Z9AHmhtw0T4Dr8eLJBzqdfRAr9INt
c7xp3gCsKE3Bf3BZka1fAcNh3a66rRTp9aqxq0fDyn0jjlITMSRDXVZdZ6FTb8wc8WZQSK7N2BRA
oc5T3W2Ij//HW/wLarFemV0BwZKtaQSYP/vM/m9NuyMewJi7dCeyQRmnJsAIwLmf7SAEvMRk9Zun
me3ak6ABb3RjqkERVV2Hol/3Stqg9hd2EMCcs4/eqOe2OqyZVf8spc+cxA9+tqo4S12umAekwNiI
My2o7jgrz5xcr2jla5ObUJv0XybEMeVLvGoi8t3pyeNZfSjFB8QBqALhPKCiNzIP48ruMnww+Iyq
gnU2gNT2KDjyo+k4m6Cuv/GzguA0NwfnccxBwGTZdVENnV04h8yCBDxHabFJdHa5l2/3XRlARfav
yOcTe3vpQdqWliR1Hq4bgfvkweuq6RUTX1TOPuysvUpSaB9hGXEzVh2k5duGV7MqKmqJKh19qyDI
UE5o324+TaxDRcFN8Op3LEBmGNkpoeJ6K2xa4RFKj1YYsh/gFUNMuNggDRZoOQJ2tR5wsQm4MSBr
zV1mSpafoTul2Smpf6Ns0gGurw7msKuIwcuhPQoFQbjjoHEwhG95GoQWizrqe/+n/dCt06dnVkOu
lFjkAdbhCV5r2H7lwnrmNy04PxRNWjK/X+PwdVyPTNvSbJA1tvQyiboGOVYg7JdzGLs7SUCVe72w
guVhRmY3R7HSfhpE3KVJLWkKG8MIgfjfZYDyvlBrxVPW72d2kMURNfxZ+RZCL728EQBczoN86ahG
ZZrQsJuaUlbZ4eZ1GKWqeC4FmB8375pl0V4iDVPKJG9uxJPjRE/sdEdO3cC/Jd/YdprMPXdHWZTx
0BysOc9jnU+yOsTF4ETisPNm2jtZLXMxrOY3v1NhhSUKsZ1HliQtxw9zAUmhxo+/Qzcs4gSgrdqL
idasyptbARRhRb0gVe3rEA/sAqTMV6N9900GdXrvtL0hC/5azUst5u/qMo21Y7EWUZr/HQMICAN3
+Nw8YlOsPrHI3zjygt+zcdUbvurXaSO/9arXQ8DMFpQdohNgzA/ZNl3GbmtvwIc6y6pQXLRZFxDJ
0Oj6klsh8p4C2Q1q8kbhzWGS6jgbvgHkLmXUG8ha8TJ5ZJPu7P155UsydJYW+Hu4fEoF8FGbhFza
vT6kg/XUGTiVZzFLDCq/nXYj35I2a1QjcXZKbDRI0qmL1r8PfOUchc8kr73OD0Kg+xTvEe7ASa/G
iIe3oTnzFi79bumcD2JL/w52lYehoAsd8E9wYbZeUHqFy6mIIvD58pi3CCegAAKMV0lWWoIxMD0/
tQtgJJUb0CDnGRAF5FYIFJffx+0izYybMIGBTD/KMRPmBy4XjwQW9OBc71pnT8uaJuWBiAnj/6cl
7Ej4Lg7IDaXz73kevw8u7g7z/xtA1Uv6SEsXE/UD+vQz0Liplxid769pzJbWjkkw6mKYY/hw11AX
Vg8sKJBNCTTKdPWaSnLRDRv5RXTuugD5Udk5aNuv35YzJamTocFo9Cu+bIYT7O/kk7u+TTKDaDuW
siOFgLBSGkBRs0cr2FZqdbVtm6KAxc6MRTflHn0inS/34P+v4jzsoGoMULj/igih1TuQvXxLWDEv
G0651uIEzGy1csE1RKUOYoIiNJTnEVOlMH9VGezN978TEaayygfh+ViuwuORxIqHeVlhVFf4Wu1J
wr/aS3pfZ3a/1+1Pwl5s/g+B2T2Ko0CeHQ5fFN4FD7HtOtYJ6RvSbVDAsrFgOvFN5cMlrEFsW5aG
S714vsV8dzIXw+LOlkLvUV5hx+6bytKYCLjo+A16EvxhPc9sgq6V6wUOsn4KiW3Po4zjx9b9e2cq
fBZH1nBoUb9EBwaYEYMvpFsc9F8fjo94cLzisOk2zaLT8p0tD7A2w4wKT126rCofNVCSDUyjFtT5
H052T6xvrJpuaYCEjp5YMf7d5MKaQVYzwGX4D79EVx8pScT292a6peI91v/8ep/15RVftO+HGPRE
F0r5f680RHKwbP9HKiIyVjFfdY2N3ioF6whQs+c8rUkLP6MwE1sGmJwlHepdnfIA62iyxarZw6sh
d3j/5INKX7wFDWUo2b0MQlaaKOsMm9lvODXaeVbqf6O6Rh9iYQ7weub16CQlY/HP0HzAGgLNMCpZ
nV7P+DGFWMw0wafpWZUdY+zz1iXR40JpAtVWGMRHdIwEm1X7bWadQkgyLPXsKWqLooFJojy1jaTn
7wb91H5d9t4whOxTOI8Cy9abgVEuliMP98xnx3xmD0zubrpgYys+BV7tiQqucVfVxv3cJ11I9Wr1
/A6Dwyedx+q7xjuXv5COp+JpGnISTRwZLuHgssl4Vfk1Um+L6lEXXmiHex6DVDsE/lroVV4HGF14
j1XYV9kOMa54E+snCjG82/wAM/oB5KRrwoZLWMJNQT7hMQyLp/hvh2QJGTVe2z99AViP950+1mNa
LOrkCDIv9KPzVWpFp3kgldIJiwHtH5P+BfFblzeK72Sl/mDrlyTpJ9EzYOU7mAzKlzuBqv4zoB+z
uFLRrviE2JS9VREhK61MfTqObsQawVJDt7TOuhTvanBz1yf21Ne+oUruw54cv5f+HOfq2ELGVuDz
xULCXalvl404D7e6T+9KGtReeNcdTK+ke3XFqavMkruPouowozV7wds1S9GrD98d3BPSPuSEPWgf
sF2owFZSMtOV3WvikCb3c+hws7yWaN2GGeA/N4rUV5hZLv4xVsFB4Q9XgBZEKWhkTjDRlnIPlnBU
SSqLv+jt9eZ7ncv6iEGJnDW4D9BbBjIKxjDVtOVl6BDWcyLUFk6BDT6gbxs194pAB2CPfBdN+sRX
c+S1vPA3w5f/rJHyIFLB80frWdiUxV2X3i2xincBKsECLpati+itTwonGuIKOu24p6XB4F1LESeI
0dqGhMTpm9b25G+vM7xhEPnaIJ6PwxjrDdpHaFg4RORjXzXRk5FbYKIzzsK2MhJjZOvhklFkKoxP
cT8EuHhszGiGLXGoNwLVzNrvfC/MPBc1CBBbzJtxLpPEnTgVs1dUqqwNkc8BgjY+dDtxby5f4fur
SwzzE5IMmZSFcxmRlzyPCwBdXQEBe9k5PXJ2zyM9xESzx0UhU32bs8D0Sw6Z4XGvV9mtLUYZnXoB
zo7bDzOS+64uWwaEQe6Rr8NI3RWw2wn0ZDRv3fRcB++U/qCaJrTW+VhZMYHmaHDGFyvmx7aZB1fM
3QXi5c7xdW/7hqm01MYAFQahRx8JADUKimkwFs+kXBQFLXUPPgQnpLodfCxn60+vW2ByXIbL5LM+
Iv95rYD8mMcA3wv8UkH6cNQyqQ4CNf1b6t/eTIGs562W5fkrq2kqrLdIxOOvSMd9uWXBFFqzeb8H
4GJZaLGl5h5Nc8lWfuUnOJYvR+ybFYfUTT5o3pMjEdS94XUr5zlf58YBuMKmFpeCp2fG/Z2Yrfsl
QiMMg5YT/OXyxuvAngJJZFRmnh3kZOBZpOMdysOgvumcAVr6t10rfUmqXS7qx8z/rR3KjszC8ILA
mPwoTghuDUaIVdLNZUoUfyVsXEEDjbaIRkOF+nJpitCuMrb6VrZYF+g/zbz5Y4CzO1ieSRkdmlkn
CVqIJSIfnkAtBLSoBtagRdtnZZ2HyTdjxiDMRgMcteWAA8tBSP/CA1AaeZxr3qEsYJPxJOOvngQA
AseCbZrRTSKZ8vywxeOxJV7NBEUKKoYHlMRyY0V549KvoUTRjCB/7s2hV4I16+y6Co8B5O3tRU9E
qqsxDtcTDvwRs6lzlhIw2S00i5x9x5lNGHsVTU2gLtopJ6fu12Jk+nGqneLreGwTaNy0/eq/EJn5
c6kNKf681ExAh4Es5ccYGm8b99nwUl/0v/kuH0iqQCoUmM8HnnnbHW8/BXMyLQNgAyAcMvZ3RGUU
GrKV8siK57KemB/jb1frQcGVtr2tW8iWIbZRuFTJJdnL6ssUebymjG38xmr4UXNeL5QZBJD274+P
buOcJmkc065OmYtLh2DoA1Xp5iyFx+3CJhEuHs5ELFFLQBvlqp35+glVOgcc4v/RMYE9byoApR9T
AURq1egJ6qjPn0KNEFXuCWfvY+6yplSx1wjj1FF7orzxMMdYQlSwidEj7QibY/wibtejTtyALBmn
S5NzbxukzBnaj5QgjpmKxS8+rLF3FlPMC3myggLG0m9fh4mM0BFgMxqdfCWbkDLy3V7DvunNLOpb
9I9q+sKtrXsAMPbvZO39A+P/LT1FtvhoGEjlpPzlv+x31WoL2uQFCEwSh5dKqKlR+jK+XWa8Hkce
p5b5S90dowpDvDAOUHHBsxrDgSz3x6WatojJdVre3jqHbnwe5stqQkt8UL6ZzHIk5B1NNB6Y502j
g4Trtt2em7dwjERjbRLp/tEghuwRkUCKghy5O/LVH8BqGM8p/zpWn2TJlrHnOPeglHsc8Dsr1Ttx
P2TSeXfvwmZlyxMB3ZKKx8yheHqddUwF7XPI8/bGe4hW4XwlY+ZwC3nfOYi6JkT4DU72RlpQdI72
0GuHPXaI2u6wHYA/kig+qABPS/x4lArq2F5kXTwfZLTHSi+e9iiMXJKxiWkY26ZSCAApIeQLpz4a
H1n0ckOk0AUyLHgHrGG3OD1sPk0zjawp+UMxbZSMIngk7FzFLoNmplLQg9rMSnMDLCaevny80JDX
g1TemBjJn6bVhCDCoPYk8p1S2r9RfkC0GeU3CGfj86s1a7szj5o0eaZbT2O26PYW/k6Rz1O4d1zV
tvWXOwdd0lFdHJ6YmOtNaVcOoNJCn9Pg9NsuovK+ELBOEuk65efk8bh6vezz5g31Ua5xGYu+O/3F
k1uw/3lS/pXqE4oMitQQ+TQyRtQ00L3z+804lnhEX+Yqh0DUyiO7YDjHotiugKoy7hNApaM/BrMB
09fKjaURruYhFQG52KAXmCY2/dOg07OX96XY293N1HpD0+EZBOqcnWWHQ4EDeXlMK/lCvPuTq02f
N6FCsUq8ILF0ZSjJJl+mzMM+YaS5zgnOs3NmI2U4eq1uc6yXPHaBVZa75vjH8Suk7GihZOMskn0r
sr01vA4Fe3hg8/d2RBt3Ike8bC4RoQHSC1m6F/wUNurEx2a5lWVQX1nCIm92GpbDqahiaiwL9tec
M+mnB0Q8OkITzfN3J7eKyl+T/x1vH/7gTzi06MjubK7E6VXeAbLrM5us0oXHQC87jYbSGGQ7OzLv
1CymXkdoFjEth5wS/gGHCZrISwYm2MvGcIAnzFYbckvb5Nu7DGJ2024b+VxGIsBuNee9sCIN0om4
tKUo0uDtL74+RwiKmIdCBiwX3Fmn0ATDRJqh8GTqOmLzS2QZVhF9CPQapFtzdvTVNRcQFp8iSGDY
dYuVWO14wNJK0YD7zrNhIo3qvhI2qbuHQEhoTCX28dIXTKd6AzzBTHYHnwUnFHFOo3lwWo8iqAKc
aECrWZt9ZywcDjteP8nMEK4hR4rSXceLfAKzFFne8tnvQgvJqavOiFzBJU89CWuOh0mt24MBVtUs
U4MQto+AdRnxbkAEhY/iS9Vzg3YAKnRamVcEqBLUVeuFhIMHcSwtoZC/hSBz1fOnkfRNBL7Do9Ai
SSwxpTwiRhjSlo6pQb2cwEKmLGLEM3Jyhr0g4J53u1yGseEf2rsqvL4R8DgEx2oTBEa3Yj44HXMq
J5u9GiF1W+4oL4jvtWAT3lMYhppfk8xWSW/dKhuYNebNsZdCsYvvQmJ9P9pJJKEP7h6rkDXltCCa
6CrcsBHFq5xDjsFLpJ9ogMhdpeW68GcEOVeXBcD0Vv9Ti2hIll757rxNxPO7YM4mZ12TyLtNNxNT
WuI2TEZsOtx3oxNr0hg4urfWZ/XNRim5M5w7KM6zDZsAfVgkIjnJFxYaJn1NkelvQVI8Nop+BPmd
s7SVd/YbXjG1chj1fbv5r+zDT1Ke9AqSVAFglIvnpGwuMpVryLLRvdPP66arPQ6NVbZmK3NfjtEt
KnQbKU7o3HtOzQ05yfb3la5O17W0CTxmPst4HFZSV4VW7iOCSjpI2xkOO9UP/xcoyTDyWF6XZjB3
aDZU/B9jJr9IFrTqT1f7dr0jLHiy0gawhzSfetcIBa1Wb6KnZyCQsVznXD+d7Dd2OzPCxhlZAG1W
qSBrh8ct/B1vVEXgdluQGe5rVRwMUF146Z4N5xDBKzH0GvOBaqrZsvWmfGHWnEK2gFZSkPwwgnCY
9DuGDb+lXbhsN12B/22VUtL0sP/lhZ3rvGr6GsSbxGJKFFHqNR2jUgipVGol/IV8F+bZnCulWHet
IT9gwRLa2rUfzPtwgxqcb4LwU7VJnOSptGxuRNPEEFbogW6khfd3+1Lr/jYpHZI+Gy/yYHqbYMWd
OAicnuHtPKSnn/JbfcHx+soW3tMtghuHYc74MldW96vZEkRNpsPYi3MX58h0MBj6DWE3rCr2Dh5I
BVejh8wiVDF57o95fcOEBndEo9OQ/WuK47yJhb+0EZIt1P53CKQ3Fo3CnT6PJsulUqZjmZMPr6js
a9bqNjbXDrEAwu69SYumFDQRFbPx7daTPhccIG9MB86ivI0qAN2iRcFTKlr0Dn4VfVgliWtZfU9m
3KOmn91DX2sJerILbBT4eXMRV9ZTiLt37q+Gf2LOU0x1OTRxaMJIhROe4l1ssiNp3BkPTnCZL8em
0pgztioJjkN54gsVl3PaE7BH8fYVbBVecvretG7fii3jKa79L5KT7t1fvcmiEydJNSgfllr48Kl5
OzU3+mUViBp3ohFrYJWjkNpWwAWs3P6+jwks5IBOe9508qDzA1hwNXOCXkWClnvfgHSX7PnghPSB
XQlsRD8b0uXwf1wnm//DiQwi93cZ+d3CxbZC5wpFV67D7XcLWPskHbWb78wDMkm29SmqKTF17eaR
5DRqCHFi4auXTfay7QKpn5WXcQmSFloCZkG5OawUrZCojJInyuIrY4ArGQgmIVkja4lIAe6GpFw0
YcNFvSrRkzwFHhjyc5U7mRpfuYsyREu/5w8NpApDtdoyqtSkMtuctQdE585wQJRTSVxklLKcdNUE
7xjafz79bEGvgenJEI5bQBsYJwLn9qhfDbq4O6cwAILy9tnpx+8tAmP9PatUWQy4uWyrWApL77Em
PNSbLeyVg1RNc7czT5q9rYp4lskJuWGHEgWw0VDRVGPQ526THHdgvK1e5gIFOqSLvrmLvwJq0zeY
UCA1ZnVK7NaogE62Ge4aQa/HxnI+dldUjquBHfoahEVufkuvD/md/YjFT/jfaam/IevEw/0dDxFy
PnDOAQb4YePuyIrYIk9VfKzV4ZBiQOuoj8Zcjxn+YgZoFH4t8zK89wAHMMU3rwb1iLe2WEc2Cv3E
jgW2X5HgsxX52MkinnE15ezYLtJ6vcvcelcG56ZNMeVu4o71bzmltLSRAS3oIVIjyBCgs9CWgasw
D7OucI3mFZlNUY3fLgRZAjiNFiGvy6a1yGThY8PAtO2hIzjxOPPk2udqGaF+LMJXaUvzIEqRDZJ3
vhmh38RJH2CABomsRubqAfoLWGeg8QpTGTcvQZxKg/GnkxJkJQLy3LJJP/wmEanTDjxA2XE1GWXj
bljodzct5rZ2gNxwOX34CFn0bavAB9hMkhAj8o7onHZ8XH5tJ1n8z8EiNrrukjaeQNKoi57wFnPs
4cFBNN2N8vAVLIGWn2u/+zJU5sc++l2hqsrNlp5vzb/+5w36Q5TOZfo4FRB1j9e7zEDoV5Zh5HER
jUcT62j6P7/p0+LDXt5gJvIdEZgO3gjdNFlp5QbT7iodW2Qz+Dri9PpPxe2gsy3n3dM3flQoUkJw
mKYKJgDkN5AQ0JUVPRWGB7NRXa4T195E8+p5RzuhPSJyownptJOFbwrhseTphcludx1BUHqCCr0Y
PGduvnQTTKU+D38F83MjiTPFzJXGrk2QZt5ozQ6fZ+iAO8bepdoOpTs9vM3lrGrme0SjvaRYRQsv
TXQ08+ROvyljnm3APZit0ockTOoB01P3FEAXh/NeRz5Uz75mx8C9ssBu8zqfszRcqi5KAz9iudl2
C/44HHaP/dvdAyu4X9EbLpHU3u0gx0xgGZu4foFKFe70XJDXsJY0a3+H18q8n9z1ixMylk3zgtZQ
BTxIyrchLE6vly9sQVUcml6wgxudmiebWzjbYmiLBHeBf4QOsCh0bR31m8apTSOQ/Qkg4SKduycH
Fb4Sl4dlF8N8KrygZGOf4b1C1l7/o9A6DCAmRTBIhlPMKJN1qR22i9/l5Rv/69qcIP55dYTRaZ3C
PMikVeJUAdIWwNy9PwSVI4ttjnKdPz+CB4yBYro/0DUIahe6INtxFM1qBzyYBHrlDO1cgrSkqL5M
EduJQ6A3sJyrdoAThZMHAy8qZWccNMzmV9KC5iedGnDFdU1VgOOu2vf1e4SWFDnQBZ/iljwutb6N
ngLrMB8IJ4MmWunrvg6cUzpiTvDoznj5rvBlrfVGGtX5d0x3Q9Qltwe7G5N14TYFo0TKEf5613oY
O8/BNQ3Y8wLjwyOwKTiP16vyMw2nWa3t++dKTT0ZL3bHy3kjG81ibeLowlmsJ7mpbtNSycsrXD8N
iFhqIMKW5apaVgOBitdkIv79V2sbJkjLLJ/I8rU7FrDq9Ov20cVAdQhTCPZIcFYOqu0uBgShRyMB
9G+P51cFei27PDIuTIqFBS3SdovENDrS14qjMkMn0s5X0itk3dJcelizdfsZXaPUrfSbj1iFBspN
i6Lbj+PRQvIl0Ejz3Ohxji6z46LHuCXklWE9gAqj9CKAyyGj2vh/UG1wGjxkiWMJe5DNIRtEnwv9
Zp4nNBbfcL+WA8YGxGWlhb2EJJ2iS8ZKW6iHi202x58GmGIgacc5B+Xqbne9Fg/v7lfmhMNaqDJH
6d9ttjJv9ecmCXynWyckU0b8sab44e+HfIu/E1M1+HbssTXGa9CHA0OssW1P5lxdqOdOgPlSc17V
rjhGhdoSbxl/uxh486HwHF+cDkJDu/Ocnyy0MCAVBCzwP72ZqyPJsI60bfWF7+7wrwfWRiw0iNbK
Zzgvs0BF2cD0EVtNwl6iSUtwHe2cBh7+/l3AGs7afHMqXHGFEK1s2KMBrWx9nVO8W1h3ZyrOkscu
BDnQeBCmnhi3vNDsNpyHLaJyZGs9NKDpq7Rm5sbprkrVWnzdriUJlqzMzacd7heZBknVglqS2yUn
Xl5zEk4/KRtJJSF8PHGsKZEGDQewryA/y9+4SRHumKwyjU79vzyd6dnF430GFsROcjMuu3LjKkVw
BWAvP5ElNuJVMXMhwd23/aydbkfKc1oy7Rni59/w8w/XQwuYX63QZu6eTQjPfwKhMOVFyj3I0tBY
EP5fMvOEtaYRe7g+MMKD3XJxWI13uBrQG8hX415aZcl3MK2GukuznBDixas16IEesF5vqCgxZl2S
tuR6ndGA/d/j5avwZv8BIrK/OUdZO/C3pd6KzWtBpq+s4RnjXi296XB304xoZWPpXa/Un/UKTPOF
UdWpG6xDLeIxqgG02F9XGwUa7R//AbvUlfFiwrIWT3K6NL7aR+QHf7IF34oDeS7DW4YbRywEjnIy
k7IzIKUMgtUa03XVOli6m4xDIFR1u+poOZeQ73KA7QKkcF0t26rrbqYvIRHtKJlJ6EejjG5TJj90
mFzpO5tnAtdNgZudNRP8T7sMyXwSgXdZpX8LcrnwRhIX/j3eYa0qaoNE0FBGT4qqorQF33jviJt9
QK/YZQM7ToKy9VVF8TeAVsLGN137VYjZrvAE95K2SbdAm+Br+TNYApaia+OEAeNsc3m9tNMKNz18
TbdPQ2CSyF9857zdbYOLgGtV8ZKpNccRYzemt2DodKbfOFSUFOwwfobilx2lbs3RGrR1W+eYYaeG
5knTlNYhFJktK6Y1DvsKuar3MzGRStDQA16cD66c+wYprlGltRIMpMSBeVLFpO7prtYvwP7tUHuo
jjm+3pWQAT6VBfZESfGl63mOrzRaRYTXR7FM61jooXcvLAInZeBy4yjXuvckMlaveMBcbuWXoe9G
EuVfSX7erW84FcoKmtLuVL5jAZj9K8nAuB03LfyHt1+Rz+WmkFCpTD0Xnu+1N/VfR+YNchpgyzIs
6KfD4D5kGezhx/i7xZsj3xnH12m0+uHuoQGvwIrG1nC5YH00L0oOcbTIxwHfEkbH62RHyfdGaU9A
G1ltDkGBPwQYXc81jPnZzq+xx47HBDlBhGid9/tN51D7/Z+ErbmPcvC1hMN05Ivy0YuYLwPkBhya
Wqi8oWH0mAGj/jhuxwLPzAg0ky9PbY7OQg4+3d829HJjxM91mCnJGCYuPTTuGeMGSc2uoo5Ziprx
fnaZxg6EYELj/Fl8L1elzFD6XtBbwJtfUO8BsIvgTyFljT/Q7MQkkRARdwU/Aspuo9vE/7pXxy0X
KFwED/VVOfVLaviISb5bZ0IQZGTIWDHV3qRZJNa5Wz7IDM9oQTACzCZuWoEtmAvLUR62BtPQ5bu8
jrPRscZGGVUoV77jA38yO2PQaSH9yo2kO6gRsAjvwWfLHDBHFgCrfD0eb1vP0vi63bzLS0jgt0d2
yu0NSuZVmTZcpg/PImxLN6KxzD5OSsYBs5qYGzcXLYkEbDIy9f2mJFHaKeT1fRxadcEFHM/f/m3s
2lCqhcAvYc+njBcY/qI5stAF/I/9u94jqTxPU9o3vY5msTlqYheTXNuY28kmoRcY5I//WOG6p2Sd
Gr2f852Wx+jiJLqeuAqviCFQtIchILrQZb5S55024v3/1PoUNXO7ZmK/XzfWbrinvTlze9L0OLJ+
TN/ybTKT6bKYr+uLPh0884mWLOF/dsob5Afx6KgM0wa7Zex55hapaOkU/uqxFRHZ3ZUHiX5gMG1/
rw0OsDxGTfKd38+uKv8lrDGsifrdjN/DrhdfpE/SeOA0C+bXlXPe2Th9Dw285Jj/IdH4lhyjx+Rk
4coH/7EwyvyRk2La5GrCnlx+jKPGkMIBNgkFdd4jQbmsjF41L4VzjZwzo/r9ZUrmsGhEaTHJ8far
o7xJHbMeUhdBe39OvlQe/oe8sNQN6loQEc1R8XDx41JQPUZTVQ+aMq0RqQ/ImPQYBaSo1A76KTZk
vk5V1lJ6mhpzfRdExHwcVZI5BNmehGApJHVCH8VYfDyUEipobE+b2WIePhPf14OAA8ALQdGqCYD0
0CyF029JsUU4UyD1sa+mrVBSO8zKoexPcSIQJ8JGPM/sON+3zunOUAr0VEyOLGEf0lPba2ZfZKu2
wuOK2bPRcBtpAIT8fo7oaJYtXa50OX5+aGKwqX0/rKxzc3MTZnFupaCYV8CW43usBt0T7hI44mgj
/R19edWc6ebdqZ84mrXg9hgCVuMOPzvdeH82GptAxs9tUvC80RALf+gmacW7QiCyPeeRamnnwTc1
4HoxQdb1wridOG75C9/u8sncRD6AECr1HwuDwhbUeS3y8/C5mcuJkLo96AiVgmcoTz2iHBP1oQdS
ly7piBqV1d8/SjL/3keNHye7GuiQLxj9xPezZWdqx9x2melFC2Rw0CdLpdhgretuwr8Xjg28wfTP
71GWuJniv+KznGQzsntTQbTMv6g4SMPPrLToqoXzoHDEwN4LneE+FTTqZvUIxn6Voz2eDX4o1WF6
zrmjVBl14V/U/rZ08Ru8LuFlnT2hPcIERhRPjouYqoDz65sqNcgXWnu6yCgWOck/n1PvZPzcB9BN
FBdr/m3A4sn0kmJt4g9VZvSahxaZDtD9CPXV9boTJbxioxnc6mq0Bw6KcRrPXzZR5WlEKoK1QqWh
gi+r+gdp+pNb6FsvWxndwm6DcixdYGGWvGRLizsMuUaMwmmxQ8Fj0eZtYDCMbPlfBAbWN7pADrAZ
SGm1ykCEVk6PYZb9nxHd2eaVoSpHjdicmPC6Xqb7Z+lHwVsUvoNz0Krtqbp4TFKIWvBJluGra/JQ
J8a+bWAlpkNgzow805muZ0UNxjPnIcYgeLMwO6hijfmiVmCKsqNj1RbV+WqgEKYpSrv5C2rUcx8E
e6gVIf7XLSSKxEXXqPnDQ3Au6VDWCbLmLMjieL9Q5gmVWJ6DD7gv6JLF00p3KxmgpX00zcVCAVnG
4ulVpj1Tj670Y2NUAKmfYb3ncFH3YA3ksOaXGmu1Giq/jFbz6Q31k16PNqeU0b2LTKD5UvhqS2aK
w9wAa1TK0hYd/hYP/AvQ9Kr6yZYqQY1xZ+ArYbkvzgVHk8v4uFlWvYHwzenS7RYxgBMHkDCbFZ1P
j9HSgmflYwovb50t4k3oR+acBUSKwb+ch1moaedVea0aMLur2sTdIEnYT9gPxwroDtXux1kzBEVN
mTab/JnimcGFiZNSMidxdXgOa6AeYq+0FIJzJ0olVDj/Ddqt6kPMaH1RdXaOMQQqbr0/B7h2siaU
x6EasjLmiaQTSLgEnXJexmMHflBkniiwQmDNgeMGcrNH+KpQgv0dfX1AkmsXT08UCiBZC0LT9HPQ
YegWjZlyr0iQquPmzUji07hO9En1zEXj4nfH2w9BRg2/DhGRHw4l2SUVL5uxDNqenkTKL2/pmx6j
9g80wDvPGH1dzTWcp30TvguF+bu9v1fdjaBX8vljq/ujGNEJB4ivOyVcmsZzd8h5+O/RdhhnhjjE
hS4RdjvBlo2rTohhJ4QHpfdJoO1m3a0yAXoJXkf9ccbtE0zGw5gq55JufKfymnuWzEaU7BRI6htZ
9l9wUIwcWSRyF8NPx6Pl75/KaERuuoW7hMCif76eUvUofUMdjlwA6N+SIjfTCzgZsve3otawP0GN
bwDJY1gf446LBI4OTMDapH/ya0rAIOS10giMXiYZfwVU3Mo0onr+nhu56Yi7MbQ01QRB5TOUaS8w
VRz+FbMCrrtldvKmLrDDTVSGjrZaht9Qt177YIJBknNqveeddOonYKF9xnyklv5TIUJMPAxZLmGF
tc52g1c5O9RGudDRr4VRWK8in6RxNLZJttNf70qnoVbZyKUZVJnnjHjKqdIZ8gpwERmCLhZrqVmg
GdWBkeRMxHaGc1jzxJ6qfE09mNFWzYbNXwR4eFy+5G1IOnuo9ch+SR583Y3wfTOhc7jyXtuw3gJo
wHeZ8rAL16KiDBcTIlsE0hgztMj0iMBeFNieyuO3vdUt7UcO+UEPN0a058sZz13wCRpcCapjDXSG
WmeMNfyVmf4QA9Osygkjvskkf9ps8CkJBGt/wYyMMxX2bp+6Z/1qgi2qgs3MPwN4pjWMgawS+UW5
m4eLd6E1dOTp2Scx7ZsyJBQkOEdLt/2NMu3dOcmdNvn5Pn6SVRh39wkblRNUd7LYIUrRbqqKrNfM
Atw0IehQHy+u4pk0GaVCQTJsys0e8Z10b6VPbwCxqqY2tiCf2Q+n+d1VjJQT2I1fIX+Us/p6lD57
FdYkjJjx0qcpa40VjeVgW2/oMhVsQIOPYNhz3rpqPHuIijTJFr5SMbtBUbcbiEoBjAAbuy1UBlsM
i5s3uC70e5a32kbIty5QVODbXPAO4Vz8nOgSIr8131QAbeTHuzSVhnQF/2LWzSKIePT7Xar9J2Jj
ExbdBsgizPEzLVCyoSZtv+BaPX3NhtPTRZwrxJjFhijl2k9/lA/lnb/g4Vh4E1tpShMIll7yxd7k
b9ZB78TUidrOligEcPB6Vyd/2g79xECfgChVa+x/tSOeXzV7dpO7NSK4ZyRqQQW+HVUDWmf6dv5w
4D8F/OLd9Vfl/AmLtBYNaypV2WEPS2JcjGimUaR1sJWi7dWIPnvoTneH4GHQz/7U/pjgolKc7OzE
WRhirX5vdNTG/nYodZdeIN7/O7lx0n4S6Ydh5FyGfK+M4ylCIpf3Kc3DIn4LUG/QAyIuBHykr8M6
wosNkw0jDtf3kGGKUI6+rQ3vUb3mCqvwTMA64i/q4VXzEeHeooaKdqAlohe/hgkoBfu4hOo8O8/j
THuOvz1jVl6GPFWpN29iK1EEqZZNBki9N5JJfMIxcQilFmpHZ9UkaUjvuwlS2NvWPMtzThVy4+xT
h9XJHqsA4Fab9WYE6+7OpXM+/g4Q1/LIN21ipsOjqd8ITbhNSU6fH5SNuXqbrc9yEHwjWmuL4XFo
PJFD4KMkQ4vTerNyAH0MWOZmwXUahKkCYCqN3SDq6BdjH5Qi/vpDFLuI740dN6LYXcqcAK+f4Gjv
Iwckb2N9D64AuJDqsB9c4BXV+JphxAIb06SinR1T1KNXYmG/p2lGu0vjBEgVj7unw0phjWhDl/Vp
fYz9XIY57tiZ/U2DcrrDLET841nGXqE9xDnheetHUSCqW+xict1/7VUY1604Xo8NEGoTTcZELvbW
mbvpwP+jIPGcH+TT85WOEWBrzE2U1VHJBGBnC+V9yHnEou7on4bJHbo0gEcpq2+3XDonkUVWJrgX
axFbMrs/Uef4TgbWxCULY3cKWfmKWsoO38r30S26WIOq4q55T8o1SLm6ZLNE3DtDQH23LsY2/ma5
a8Zlx+dCaaWG8K1MYe+V8SopvNyOvOt0e9hikFfCToHHaV8FG2EcNnFUhMCjaQEolYxlqRwgfEn1
Ud/5QTMlkEBK+N58Dn7z8OU2AP0sa7YxGPxHg5Ik1hXheCiempg7pSX/Utx8B66xCuhv6u2rze36
gL35nJi5hc9nGwR07OjRLSHz5NM4McIRULmP97kVpC68rjpdcK9rl92ldlm4frM15LkJ5vNrPBXr
0xEKkycyHIYl4URXhNXVC2QXvpjdZ9u6FD5/H3FG2o/nARq+KvGEYn2pNhL5dTRY0IWhG8fwA4fn
QzEjDiHqOfeAW/ivFjBCMW1nrQh2HqiftiATO83hURrT5VATUkDtWKHDHnREPkfWV0i01vmE242f
uTPrV2uVUF6ZqQdyxrvLoupZRzyZR0c2wUIqH+Ldkq25jsoKjnCPf2atj/Z+RNr3PHUpuJRhggl5
HmJnoR+AM0Hp6LIIrCGZR+IVQ8KFxyK1bmegBABP0yL7shBbEc29wgB+9D0WQIbTXIUnHgS2bh/K
N1lJd+3HZFTyJiksxj/0PqTqiLyH9U2qnT5NWmh9OXExQXf6GUph4sQNOp07OWovxR7P/FYUfYsO
2L4pnxGqd21sFKUZkPW0exfC5Js6Xn9Ibv1wIQTgUCzKdz5V8R81/+Src6thWy6NDI9f0D7PI5aZ
KrgDJnajaTv54+mLun7Sw7rPwt4ozLSEooZ+uXiV2I9e5BQRMji57i7z+Zgt6ssot6MdtmkaFXE1
xQLY0aTLzU3tGX78dNm0CwOHLg/cms/kdd5SxZ6xBjjH6hLExNgVWV4N3HszGOlZG9LqPQkRa1GC
quzxeC2johXF6gPWI1EIavvXPKEqCSoOtNQxBfDd/NxKSXmbPPgHjwshQzfIaapHNzMi52BqMmLb
3iUijzQz0WuP79rvypYFo4zGHKHadJ50c8+dnZwb3iTaggF8f9UxrYHVGjLxT/YmnvabFoVouA0m
1AbwwIkFGfSIvhkOC4Ud5dwnxvj9TMzDaXy+oOV/o3n3hxEC810Kfbuj0KTe10A/mb9NkFgF2u/l
76Xkxun0M13HgO2nbKeNb0Y/N4YzmnB1Xv6qRp7F68ww2pO7yToaQnreuc0Ph68e4/y0dpOpNppg
W55+4v1NYC2NTsckC8ivaC9VXo9xPo1cPnRy7G7k3TMJY/fHQmJflk60DowTcd+fjsjq/eSWVK1s
OxGjeYe4pTfQ1i5ZUZNO7p+pMR1uc9iAphqHTEMoytiJYgrj/YumNko4A97Fk0Cy+iGSiyMuQ49B
op8jh5AJT6e80KchfyrsQDh8yN1XgJhaO5fSdjigEK4npuRF+sTVAAG32+B9gDpY+CIrnqo75xM3
tjrV4sr/FpItbinhJvLGtFyC13mF0uwhVW+nE689d/Cr/XBLYjjR/OXGDc8oV+00XPqOhAPcYwq7
1S5WQs5fNlpsl4qSSCqmy+OAAlc8DYEHrS+ijhFZdRYbHCiwV3+QEVpEeIUasZ5E4dUuG6uWiIL2
Mx32SgvZVfzx6BuN7LRrSArj4cYeXusoBD9pgb2ndTJaEU2na4yDx71OlPDaPVoTBM0Be4/VDSJk
Uq0uYyUYy752rv9e3Bt1k19Zq1QQNVkLgEgdcbtt2y0G1SsSwW5T1gVuPjptTRquqbjfao+DhML1
YuaNYFB30AtfIX4KJDilrsBMgi9wqhToByTwhvTPAJudYVY1lTd05WTcBbw+JcWn5QaT4akoSO8A
L6b1psKE0qvZEWe+RicbjXCTbmOhZx8oU3GmMvDdlHxpXJlAlIlbjQBAoO752kJu/fOUWt4cCMNa
Tm/sC9w2ob2vBs3q6T35UheqHS+iXlI+7PpgvCV/AjTyqQTW75xN1rgxTJcn0iLFt9GHFZSLmOUy
wmqDrP5LEbjvFFRU1gU4gKeapYKhxrvsi0aWJfrNP8AemMKbm3pBVwBlMHHYDpefxZn7OFrkRXBL
7dr+d9JkxswQVkubALxK1Rgmn3g2ozsffwIo+vz3Nvc2Wovm6IQn8ihNSfAk44Oop8mjW6kCGJV7
wv2YpnM69/EFO6aahfD034xWi+zNhqQ4gDQnfuYm9I6jCWXM8I9I3bSnze/JAlvPihuUCfpYSxfE
dbBWgjR6mWqELfIj9gMmFjJXCg/b1TLbzsCAH3373vUqJqj1jajZBtwpv85q90d02ACvEBbrvKiD
v6tk80qeqsbNOxk69XSsYTLt+AzFQrgsM1YUKvkRRv1ZJiraqiu4IICR0AUV1+yWPUpvKNjQtZMD
4SWXTNN16YsR26g6SKgWi45jThZ6mEaalfidxx+5djT2pQgZmV/AxXf5K1UWerCgclu0e82zyKw4
4Ux8NLRNe8DKXu+sN5mu5RJrnQRNnz7L9wCrxH9YVcCD73XixihFhIJUsgdcsq19wV9hIQ9jtkJA
KcdLJ0DXBdqFkJT/VgtII9LP88LGbMlrGjW7XJ9WidmpAWZ7HXLmEXvzT+K4IU35UuTNjawdpWut
yH74cIIAQOnf/LlHwJfoMc6+R0cTicNQzYMoj9qsrC7GDX3uOA1qJkPGuWfMcUc7CMGimKqp/b/D
OrgHjqpJ9zHV+/zbyyGvQtopgFUnjlxSyCuKMAwKHbxB2vbzqdjZBIv5TrjUYX0VH/+v4ojQoVS5
lorKyqQSmyH3WIPjTB0lreEzN0ofoHUzw/eKCNWJ+aAlu1CnAkhCzYZCayUCscnYoIGhMwdxBjsv
3gkafq7j5izqwsSS+C1tog6wjpEGh7YMtjsLPszQzDyBcwginxuCjBZRTEsCfWT3cSFWTGo5JYvJ
Mrwg0FBAiB2qAzEQsfVM3qRyDM2tV19Kj6Em/t+YV2aTh9nb8hJ6yO3hbp3EoB+rRpHDh6ME1nE8
g+4MMyBeNIrvj+2ddPo6dk2FKrVYWHrJNPYs8lp+R3iyX00197Myw4cMYbJiI7FAuFkLZVt0LrEy
7wU2wL0YTPf4AIsc9/hZpttwDT/EZBegQis26lOMlj8U//+3+COi5eB93f+6iMB8BhhDArWcDsWw
CaEy1pQG6NChzdVbijBwAajQyQLHZL33t/gpSwCN1l9N74AZdjQ0fdTRH4rf998FlcnRfG1zJmc5
MRfrp1SURqCxiu3+FTxhto3l1NPr8nDodss4vcOxTO+Em8fcehln8GwFvHrf/eHUktVKtu63Uq6p
sPX1Eic+rjlvXwYrmitKzS/syl2awEysmLK8W3tMp3wtSyR+t8sUyZ/xk51Sb01NWo7U5wwqDK1Y
rmPGwJ2AHiBCS9zwi0V/4durj1Yp0AEUIaGKaxPLzditnhUuHdPPy4bNUMMlzO7hHYY+O43L83sB
GfEgb5ITAX4BWxN3uueec2DfPUznGUTGg3ozaDNBQU5YasEpaMRlHewZuO+qXPb3zkFe6h7EM8af
xfkm+VceKCZ7qyOn6FAdWH9+Ws6DHFJvNeJ+oQHH9bvhlSd6djqt4vBLrVLkDj1kT+xBiUSsFdUk
2jjcjwrnKt6soNeSJJMYOYMeqUq5T7pzYmdvnlwETJCP6rHktD9YGDDiby0zmxdX7quSsxUBZaO1
9QrqvErcD8TV61noXqxK7LihtDB4Mb+iVaRHnP7WE4KRWEitux0Eh3rZaNHqAndaMB9eXGAf6xau
YXUZK/zbOjeLfoz3nGU0HCBqVP/op0yW0fW5A1l9oTQKwZv8h9gBhWeWLscdwpQWTKDrFANL6hdG
ZLIgQ+0daksTVblU28+N8z3hmyWxzlFs/b6DX3vuJdeOhdWckby/R8P/WGSWpYnKxwVFErEGSPHK
h3kGAC/3bhBqY5tRq3PZCMIbwT4+q0/Dka4cfBVQGIzhwqCwh+S/QBG8pd8vShN3VkVzeXi+yFda
eWTK1DZc+iNwT9aBq/n2fhu6ccSCOzIdlaenLlLHaHGTqkzKRlA8JE9nFvdYmC3bAlXJ2szy0Bla
cQ+1NnmlQKkp08V//1gqZLy0lJ2ZIujE9SoxPW2LKlBegOvOel1z93fwn6bnq5NDzVYkvJoUXA6O
Hp+DOwKizENjgiAdaW2xJYwOqEieUCHNsiqvzRjGejL7p9ULp19edetLqsCql49zSNa+by8BveiI
xZj69iSU7bU9/IufSamYWfu2XfrMFRUDVblhOS66TwGxcJJZ1m4r0cVUaDntKa7+JD9Dr/UWkq9d
/ebHjTk5kgQ0+IM8+cOKomBy5gUTPzy3tfHUIt1c2vHiczDiISR9/OJIzVOvn0hRGBZebF6Eje6O
bC62nmjPLVNmfB5fXoNqueoCOt282lH7F1lPye9nRuI4n7+LdnJ9Pn9vCdOrXgUPRcmkXb9WzG3r
RRbNqaPhySdTIzEDAhNKADW0jxYbOWFcd9KPUn+PMytUZ7KGMnCAxnkd960z1rQFY2895ikI91FT
7QVlqHyUk/tXUf7Rf5+0qk6mnZtllL9oPWIrfiiZaS5vbELiR77QRnq0qBF9JykrP6pIsAI1W760
+raUENNIRkKj76sCi3vCpm4QxHLHviwtwtB7CHatOCmUDwbU1I+7ec3dwhtANix7E0K68wuBCYse
357Mw5Od0PyQXMir3iQhIgKTjPyqOwlIHw3NxTVaRYP5pbbYFyJTwX7q3yyhYiy26XAUkBup6PV5
kkTiXDDkw80eWkEtLGFkYwJHCBkwWG7X5GtVQMWKjys58967cckevItKWZmtGB1voknNy2fVa/Nf
3byaJAuAanqHeS6ZTsCnsX+/OTUp3RZ7cTF0RA/u/H68HHQk36FRa0xe8OStPuSrjGbfAXM5oDY8
WMMqIFDQNjFs66XEdZdyvgkLAA1QVHHOuvh/SvTJSsSg+/nOtiCQCeXiHOb0/WMmi3pJPulmtz/t
bsjIJI8k38U6zX5huaP/BOSI/E2AhpEohCN3wauVI1ToaO1MBMwWW/tD9QnASys3BQBPL14C2Qt9
rnMe63aatcpzPOoTegedO6ECCPxLMKZyrF8FOb5kBEjldRqhB7r2toRHQlk0CcWmDalJRyfTFZvy
v9z69udRbDpjW3vFGdYesVEYEWrDXU4FlYQjrYGz2FNEsAMFeSKVStvUfOz1uWvjreCDANZlLesj
WK4vHHdNOrO4xLmKQn2kVuMXWWU4IbsoBmVZPBV5IUWMvGF6V/3jgsr24XbZRHuj1NKsBTjzkyKv
HzJW+X4pyo7i34ggTpR+cewgfyygwXFtgeP5QR0qZYXUWJ/SBTev87VpYJz3U70jywU8ycciMk3J
On0mnbT3kS3WzB/vuvXPR0bFZlolO+URY19e0I4XZeKq10oLw6ZZg/HByLIeZp91w/g6Pt8X9KLE
vJdaxs12ZLrq0eYPoxS6xmip0QBVX0MajeDTBmXVARmh8GTAbyD+gCsolwVoBxWjxymwiwdA67YB
ooebThrqwe6gRfiadkuxXVplpN9nJ4YDk/SpD86ems63cb/Yg0JtmYxX8M2RrMieCMyyWUtbGW9h
4HSsGml9aN5svU1t6W9IlmAT6BPu5Lk1/sFRTfU/mOs6F48R0SPFwcy82R0iT6MMRJk77/AdZTVK
Jm+bOm4WRfF2TIISrip0h88eyAQ9Mz0lj6yhVCukYTBIP3OzqbZJvQR5r0TVD6p1PqELCCCYbVmk
ZCowIlKYBbUwMYwVI7XVgbepH/1TYlldV5Kx47FXz88bbvzGXHyj/EHxeblVBBy+y7U4OfpYklR8
YYHbzVAd3SmdW7bQoS5RltDFomEeG5x05JkgaZGmi5XORvwaTbu3+slqq+3wyc3B7fYiq5U90kQr
Lt9hQ/OEkco8MIcUun8aIDISNNnhuXxgZCZUWkkVaAHtwsPDrWHjYaWJVEkzqDJR3aFBnPgOCilI
ZbSccvJkQP5rGmzYFU6XCDVfOl0j7bjI/RmdJga6uXQYzrtAk340awxKYYv4aLg2VemtsztQKkrU
N5TOhOQnxwC4fXcu2re46O0bI6UnX9Gtw1eRk5tFXv6t6FX7Spy39/KOznCiRak2rE6NIA3dsQ61
MRb0DZ+44WJaHRbS48u+3125jQoPwePFWQN1EFJxZI64VVMnT4K3BV4jaZVaPTZ3zqqoqBIfGL+V
uycHNwGNIgsgaAPddGk6i13Bq9RXtpHC+hSkQDHtH1ychBfU4034hnv192rr1yrhrqKyfC9k9E+g
f7EDLtPSM9uRSYKnUOz7XQQ4H1fhODA9tLYu8/HKYFTDOHoypckG9aQevSeRjE7lkbJLjASYT7U5
rHw4Ccedm2kbe9pgD2t0QSKAj1feftK56aaSbO5/dJ8bqndfX750Wki6MLsySPjHt0LnCNvMiIMl
STI2FledR7IkDhCqXuaFHS9w8mvp5anTBHYK3j/UF4HkexGhoW0t6MU8WP7XPTlaQdGIRPllu2yR
w/K7GLEWZJHdMiuKvMdrbd4kEIla93fGjJSTQwR2cfqF9zsZtjCtpTVukbHCaQ28K7ShXAmtFG2X
64Cty3FyjdNNESDBCwbDt/qUUFTD8X5HdgWaCdfdNDOIPhIr/bbcdQOYW3hEJjJaBZg64JB4Pxpk
HhU01s5ziXiH1yX98W7WamhaTGANuYDuGqOm0juMGT/+uc1ZDwQzay8Mq86ZKlxZ2rQZT/3J5nw+
/A/Q/05TUha223eV9yfqyGZ5VmacrdxmJ9zLTjXkc6CbHKIlATw1AVe5nuJdPdJ0bBHuOg60lR2w
irUdlNxuXFctu8BvzzD4zP4FmLQfjUcSIJXB2m/Ehcy6ANui648/Z1j5vgjgvrplQiicG+kk8dMA
zVk/ZmYb0z9ZJUTvt5LxSy/R83Ed2Rx+jeEPAKWqVLSJkrE2z1TLcI6zrygCU76y9aklYQRfevKN
HxT1hnk4U7vLyjAWAg/+8XZsV/nGwO4DatHpdcy5ruj8ybCp0VGMV3ZgUp8MH0tdaA98Q0O9HnNu
+CswmNJydOCuqsq1XUQb33Ta6kDzqmfXR9eOLBCG2RjWXaTJ9/BiAVjS8I/J/OXmEZUxCZeQCQKr
VCNtrUqXAg/mNzfTjWeFtEPEZRH/JT7Q0yP5h5BqfqVomkDWW3+u4HF8EZDFkK2+tQMlID9oHJlx
VIwKh6NyI/slcIMuTTpFOPogLQdZBB3Pny/soJJrQFuXcVimWJ/1/qfqBK+h/t1mgCWRROmoKxiI
T2bNnx7ndONpeUljTLOmVfJ1u+vXV8EK4ALpM04Q4smAp6Mo1bIvpem+Ok8f9Gy2S8pqzm1EE3AS
ULlKl3CNScSTv5SLQv6XUIrvWE8IGgSKRc7m76eSXOy/RPWntkx6YigQPD+XYWrZ9rhev/3LS2gP
Oyxtbc8yl8Az+cFd66NKbrimczTvL0mM1ZAhc9gkyJblxL08TIofWaTdwEmRgTAiWkzOip33s7Gu
AsDpkg00gYgL3pp2QB4su5hB+qqzk7uKQkuXhLVkh35u4V2bPQoka/FVQFrh9vQjeqSoP+4T+RVz
x1c441IsJGyykRBXaxnhVLmotAPLoXk29Qt4JMiZN0rXTyuz8HwfPqI0DxsGJmf1j+MRam/LNkIs
N8HK3stKA9h7uFIHSPYBqdinPmzJK+qU4/7tgsEeBruNVyjTAzRzGiZrgB+X0JJ9uPFL2tSHf7EU
/Yf0huROSI6LHRlVVa6ukgp9IaG/gFRWujsR0jQ0tHsGZtJwN2SaI+Ni2jsZNLU5KFaeOcoQjbRA
TchSt2BG8lslk4uxy5ixsP095d3ne9aB3DeVP0e+QWYgEdZjamajUZe/Pi6hdGxdsyamvd8wUp5R
bAyG543ffAMkDaKUm5XZAIsMpKNBaZGZe3at2y1rljVgJGHnzflPb2mTonr+Nn0H+g1BGz+zbZBo
qbYDd0TM7rFnjcpWvtNdiKyzyGPZfBj0QKaK6BCD3I9t6W4MV1RlL/sRcFwofeEX3hr2EtO6J7CV
NFtt0i2xD0IaU3byrA6XaooRMKja3/4SKXONM/WIJce2miRMGhcrLm/iRiSNvF4YTBCSqHZCS4xv
ju+QJAJtYYh4v9kEQVHks7bmAbgWTuuZ5UAzNn4LTxbgnHdoplOkLR5sJmlE9VrPGYFCG0ltPZ8H
4LHFg6AB80m3jmAYos153aQL2qX2pLp+R2Baz51NPe+wNerI8LIAGrn3FgeSCvF+wRc+MP7qBdpf
KkPp4mKfuoXf+MwlnMN8/CYtV9KBGnRkLtGBY6s6IC80CLmg+MeGTKXTu6Me5mlpw96eiLG87J/J
WcfjMzUsclLmq7hV6iyyqoOOpXbvgUSEoVoI9pxL1roAweAOjQesLpaH+c2zYTFgVAOyBICjLumD
zHZM1C4upuev5KABXwHtllcHie8T3aivbmjuTEkloppcmiz83ZPP6HLK+xeLXlDKsIFFRCn0g34A
h6O927bxFn+OkfRZGlZ9PDK1JJI9l2wS/jxFEgqOIF6bUIwGiiNhnt6roqz8XWOBfHDOp+Usgt/b
85cR4pQnv01VyTl5jqlQmLjmBVEp/iqB+GSF7iyLpeE8B1aqzg2UkKf/pYOC+kF6UkBeDHdd9gYJ
EasuKXCZJOsLA8KntGAS4rRVuEvh4n+uMBujhN5UROJtnGyjPgj9TdhPRSUUn216gpoxdDskCnyy
eBvO8FNHbkCfICoezaCGG61T6WspAKA5gOfNsYU/cPXhOuKMnoXq9fGpLx3yHKU2Z+qkc1tgLIWD
dWSp1HJOG52cYJfO8AdsetuyUN4350v1ls97Xj37dm01GokeslSignMj7tv31knvr31N0/ZJ8odI
ushOQUrCKELP4O9WOSXW5IJjdKEGGdQdT29J5zoauOFSs8a0mWUUDKOYHkxDK6MXicMMbXCS3nm2
nBZj9M9dTzNfUO4I41e5a4OhkupwWJFYwWBbi/E6+kt7cpzYPQmySFo4mSK6z8To3sRO4b4XfAHh
zSuLh0TK5jRaE6suoF7Q8R6Q7KHwTwxkLu4i7kJFyW65D9n37F4xwbkoD0DKi4hLRLto8wCPq9JU
eyong8d/K700qy8d3cXd4KJiOh50sncC7aVDrZc0W3HPIIcg9l5mQN8js4dT5nCsEEkTtD3R5yRh
mZkhP6vH4YGcrjJsDh3WCWIQrZOfXdEIFIjdC0Cj6sXcnaa0+dwecP4k/9ycb5DpInVfb8rtcL3N
LbOuJuZgRabRq5XwVk8rtZMPEd67svCfy/PqolArRmB0wTqHrYUHZm6rBPUZHIJKLV0e0LMsSkF7
7X6JD3kx63uO7+lo2jeU3cUqhybeVg8s88Mul5t/QiUfuzxxvFp2wt1wSYvYpheIt04rVRy6/BN3
wxF6dny00NN+m/23Cqto3BAyVVHfl2kRsmIORxVYfRlMo/u1bCqI1qmVGXgQykLr0/w1GO4lCFPN
ODX1UcHaA8ZWVx66e/xs604ENTqOccrWYMpqjF4gmStY/wqgEDAuQMF9fzB4OnLT3f9FzmZPY8aP
wozTAMFHsZa1FaLHHARmLKwnBTefiteyyj+dufXjBN5ZkCuDMTYoN1aGRC9D/Y2uxhNVpy/uBwGj
Ab51U4uhnUa7G5qCP3y91iIQJiuZhMvPZJcn8lERQSkYx1UIuJNxk/viI+BBDyy14Hw996JdLBh7
KFI1vny8jzMPqn/QpefhcVocg6Zbof9MaXp7SAnwFhegcxgv78T+cJfDMBUloEW0XfkHew826/Ov
W4ZL+CEWRzReEprCWzNBY/+2uRBv510O1cLbD7tNCk1/jvOcrhPqOzTN9J+HOG/kD5uzfb6QFvlN
MKXahllnI+GtQf8zaTy6qWc8LToZwhCTkN/Gf0ED25woAEo5cO8H/2QuNBpdfNj5oecUGptFRCLz
z6K885b/ygf7Isxgyge9mMCXVYZP8UiLdnZrTImz0yUqQ4UfCr4/XalcwVqPSlVtNYixZI3Z8ja8
MQBwu1mp07STwq8GNDDDeVueUotkVrrsnEwFWFKPPG0OJMdl4s/9DoKqKHf297aPchMlu+7bj7Kw
6WS5HqBIo1C5nFe0HtU8dFXxD7kSzdgPG8gwcRXjGxu+OSU8R9wbTPCNCWm3xZVJE+Sb1dJpscvM
fT5MMC0sXMnU9LTJ2/9szJNYKX29+mouZa445nfRlJBc9Xg1cS0Zsrtusl0yRZKhZIk58Y3ylwyc
jphy0AjUMY4lgVWP/oCh3KKnMNQOZLbcfzfx6D/C/4eHil1a/yL08DSyNz7W+JJirlWjalmfAp1T
PsE2F4QCBbLfFr6vv4NXMb4MOJ5MCIh2LKGqAm5ekQIMqPClEOwKTGDkwZefRdaPhjCo8YXCcZr3
h/ExP6+VPSnX++xIYkI57+gTpO2T68heboPtFcE3+aFLA8uyvXcubaj64mfo+0Hb5R0x080oKqlT
wo6aaoxh/X6Ts9vtqjd1cikgFHVvQ7NQS99QEeG6VMXcER42ER9LYKpGDys8Ttox/Bt73ZBVyYWZ
593J35MlT2H8jroNtiuaM0sJIf3uxzd1rZ3lZFLCzcpDCKFH8ClF66rM9rrI2yyq5jeK7K/eyxaq
oiPH4Y+q0TPI9OUTtbTF7OCm3iXKBFE/b65PZcdsH1EDJKzdtzNdVFRys1siZJjLrusViV9v/89l
+Jzv4d8dRbJ+dhLgzPRhrTnot8FZDYk0phJqetH3mQ7VUCCJYAJkdxspOb/6WZ0IAkLaY1J1z86p
o6Fu9qbQBdy/jP/DBNvVPL0GT7y7hZbqrpKZsBpLY3mnw3lEWetWRKONtja9SwgWjTxzX/+oSmNe
xvbZRAXIHyHCYOget2OHOA4pCk2zcg8aafahrxck1Ho7hB8NlqmNt665FC2SJGcdpccSufPqRu9i
+eLyM6pSgiLiIPpEdaC+6RLpZdME0fXnBpiQk3nFWNhZ/fP/ihQnutWBkRpAOhA/l72ANoPsMpyQ
rEsxfyNJiUPAUqcCNnkruyyEqaQRdURco1Q4mBlaaklSS8DQksoEjt0aseHZosApHUW7d3PjLcZk
yaBJgrovxT5ayuAY1B9yMVf2SIAWyCxC8mZrQwqgims9bw5nxWCjkKnfWXJys+KJ/KkF1j0zJ5hG
ZEp7BUxUelZvWKyZFVuqeet6i9GqpSJadhWWNqtWMJslzn08h7Ys/TEEotDo9Fo9+qA+JnrDrTMA
znbE65XMF4c+tBzc/gjbbrsjSQlc995HLOnD0nEbOJkC84YDT+VcH+QRq1+q7N8BwOtXjswqzPWG
YTKV3lQKrp3D4TK8HZdZ4b5bKutwyw/h/a4jXTLCc9YqlQWAX7wKUC9AB72qPAazAju4M2l4umjR
qTSZyxr8W6Cw3JRRl3Guyq968TlFk8Uq1QO7wpcT7ATNTHO51dZ41H9s37YYZ/EfZeNM98NfJQJF
CVgCKslnxGy4jlZo23wEehWZPnfmMtj+YrQTIIdB5rkqaNA+6kYa7eNyZKx1LjAFN5G75dckFhou
mQjhQ1IuRxaKGtvIyIJsS2LKyztq2Vcy33x+bjaCJgRYZ+C1vj+p09XHwBRqbA4q/HBpd6kNEn6X
jvJpdBw21ZtF7YkDMutlPeeo8lT38FczkU5Q5bGWo29wLk0HmaQhSlCXBOhNRm6Y+AmT2bwprAdJ
Mb5nL6/5zN9H3YqUSzxAnMsOTDIprKwCCEwWIWFqtS6mst7UUOuYVqDlv7CxS4fzdLBAWbJrpU6J
FbYy9EOZA6CLZmY3wJKm5xyC5LJMbLVjLfQVP9WmeqtDJ9Oa3lA83TKMOPdaz0g7T7pBeRTqYTnE
Ik/MRo8Ku01vK7U8gZxeOBcS6iyMNgPBWNMAMp4JQmTvf95VV5wPAEZ/bGPPi6ih9R9TQvkmSEzU
zyj+J5K7kpKrkkMZlOBvvxO5lu5s1NxrP5rVzMSITKVAVjCuv3Mx210dnVvmOiPAqhjfowrKOJc8
qrBruS7fTckWeZnKfz9wByLHyuo2ovKsnuqRVsXrsFzvwLEUv60d3sIYdIF6yph3rvZlc8NmE+yU
qyVrcdAQgkLr1zHFaFW7hhOpE/RjRmz9Pdk92LUHHxh/gDIlCPJhz/zL6h2UD+LV2a5ErZ+nHPpM
HDBOiu/MLkHWFN2frtzS3XGOO7UElT896dN6+OLc+eHigDVkSht+4x/Cpz7UvLTCZTgef7GoksTq
KIZ9F34up5SrswGKQkiSS+2E8L+FjnecKN+2EehCGAdQegAMkQzLfD29U+1B4tiYgz3JYqSvbVpX
+W6TcvmYklwx1/6gtvJrGr7V/mfNJ8zfnl+EAh5RI9C+ZPirxHmydmVNyssy/TrX59ByDf7pt1hq
+rvaUsRHv+AvW97Bfs8ZgUIk9rpVW8onx549Q4HR5Rh8vp+KaVWoyHuI27q5hpKg/Qtz8ohQyjw7
+c0OV8yN5wcQdaIsRcMLXqs4xY/Qr/cRMkSmh877n4eM27gu3boJDt95HuMnmcOGJvgPiEiYhYlN
PHcqMZuZA3AkfxFnVjjPwwu9C9clhMWp4FrqSpI75kUAkjjmMRnKIpKUJqCKqOIeZiBxDOup5i9d
LEpLOiIbsyrmBwJ4ilnEMzkDxJJ29N0MYECnlYWQGVuk+bcLR7cLcwGRgSOsnxVvJ1IE8WIdXdDa
HJSOC6J0R7hNQgxQalEbkj5Wtl9tqIFjhmio88+VLUppxVAzJIx/QM+O/CXT9k4rqnLaeE5wRAQu
2E6g4DE+IZYvg9JelgSUiV3F4B8sW1iBsIj/kU0+qol1SFh8AJ6LCHpHwVfpZ02lojyrhxmDtgtg
XiKLjHNclMryiCuOAk1LsscijtQa7j7KCNMsj0ioVzDnzf4XE+1juSt6x7A9p9/Mlw4zmGmxJp0H
h5xvRtLEuJPO/Bw/n/IjDDRN6grY1AHpkzoYC3jUYPuFI0FkA4X6CPVtsVO5Dn8QMtXl1N5lXaNG
aLDqyTQR39dFLGUCl6xnEn5qUbYSHfTev8YhsL1aI2GMIjhf7bcfobPiaIcgukviJuemQQ6TSpbi
5IkjIH1VwKr3w/NtVURRPW+mlUjSSSuDZ6R2OxpFhy8URKwxPrU50FOQ4+aFJ/riWob8K8uPRH/m
RNCh7EWmZH/2Cnw6ZNqmm81ZAOhgTP3MJoXZFwH6yCaKHCdif9xx4pR8Zsak6hU6Mk9MlJeV7+6a
VDcH0rVz9GToZrX66ll1db/6DpsfpmkYofwnAl4WLjEq+uEmN9qgSTRXpTE7w016E35GPGKyo/N+
vtyD3Oojco99YfgUhU3rOUZUKELelaZV5WobNh+/ie/ki9Ezznz4G0vck+gpoiy//pQ5BE4WOjuG
L+jA+DMiLaILt0ZP1mASJOXgTljS4Dyxn4ELuuW5kbDdLxlHs9I0IXXae/YIJSik7HWoS2w0hvu/
qRk8kkgtI+GgaZHscwC5+eabXJDivLypAw6FJhL2WA8q3SIfL9XN+2JokcRa5YFDi9FNczkM6Fl5
cmpjS2GaSg1b4+CwBdg1IClRsj8PIWRePZg/75tMogm3ObhVLmn0za9LpDTFK5LUQmiAVK6Z0esy
pq6NuXG9oXcTjqBhf2uH47fa1gax6I/WijFsSre3wFKNVg6ipx22VB5ByWObq3wa6g8HOp4VKR9K
6yLd8zgfb2dNXwTjwJ28CF1noiu7fjDy6JUlGsxjFXB4AsaELxGTV+Ef4HdF/7hy5nvHgpKSSUs2
dCqZNqZ//cvRAy45Cfs8s0aHhlbl28Hqxe8DUcHK2iX0fh0I86PHxXH7NGzsnyPYXoD9AhbxcLmz
S5eSmmqxuMQAm0IF4L32NHfO7qlxMQ0EdFk2VsCP9bAbOHBP6LD488+BtDEj/zIsU09y05Iqy9bQ
KwCGOx+T+0prhJJv4valiySKCw0HzCTTykTT7Phkc5SiX8gG/FSkrDr2pzpCaaRUqwVdJSG3AE96
h/rs9iJjpI0I5lE87QLL2cGtL6iprSOvtQAcEMkPQ4Z0hSjgEw3/f76bw23hr9dkItMNBe1qVjVV
gfVIhVtnQrM/7Ro8JzPIBIGmbiHw3/lBCRy4vzO1dLYWZcsYFCgnyeQ4F+N2PFgY3nHaeQGg+MAN
uJUqvYktrUZ+ELxjGeqOo/9seIamTIo8EWtxf9v18cl2nFcdSCJ977cpfclk0glchXCRQo6Stzqf
tOuHtoYN/WhCndQliS8KfQpOHf82YlgTFekoILIPMH8ZV5irj7skBRECnZu3EGcMZL+dbO6jb4/a
bVxauKvwB+ZdIXnFlY3AIM04+bld9ekxsWI0osbG/ruNE2nLWNcnL/pDodd2Xz2GqbejwkiP/W+i
Z9jN+/jBfcy2fZNXEyAc+p0clss64cy20hkedNX4k+YAjk2/FoFemmJO4+2MotrKVfdqctUni2eO
5JnBLbMQxWlGfMJsS8rN2TVV9G+37T7bEIaYGRHvRUjEKQMW6SS6BDIv7aBdtSn8PQjq0uNywyC7
e65e7Amhz0sSQiPyYmakP81lEUeq/s+rjieHQuAJIba812yBAoIcLrGTfuuG8+iS9LWrygqRSvyh
8KkHt32eEtAk1FEGfWLL63SEocAA/J4aTWyp0D+BYkbLwfmCvO4g1EWLFdZbbYEiXZJ01K54MTmt
um8rsoJ2upV+T5rT0mfVwIPlo12+WNIKsO0R6tmGgX97VTf9flK+F++GkJ9J9IBl/4BS7ySRA1a+
XVwHUcg8c6+tj1RMOnsKDjbpwGAl+Nl5+fGy6P8uJkeeaXKY0ZkiUHRlVN09RKcluNmf6PEHMQPF
2SwH6qj634w7BifSaJGcD23PhooKizECAHWnMsqvIT+gXbR8RvGxKYpDi1XK8XojrEEIuzqGI7BU
G+RbhJNaqD1zBdE8uXaJsQQ+Y9Y7VG2mxZ68MEOm4ByEjPww2XgTZO02Bswm4aNhOhtGQk9AslLL
2LyI3j+UY7FimyOmw++zXNvCHOQxSj3hxLYXOtEmAh+2dQ6ICTnZ0nFr4j1wVSR4/k4a9lLWQcaA
eYj8a8w4TELP0BU/LTjg4t9puos37Dni7gySxwaCw+j30/QzKdyFx8CetgBcv+GvxTTmD/lTwBEf
8Em3zpZbDer7gS7GKJ8FgI1R4JDyK4ND5ivjhd9vdzL6mN+Ok8S+pagBBQXeyVmqLrDDnbIUHxbw
lXk1wNgFN7/3uS5fhr9sivqlLapRCtXr5dkgLn7af65hDVM0bpio9r6rfcZRcySpaRLiD4PTfwVF
YmJJWWGpxDAU0RJt8SakTghRuaW0UjvV/k0nijxtNgxoEpB5Ci1JDBMb4mB8IPQRx49lNVb791YR
BF5caMzlOKKdReZk/Uey3zDVoBkybrZJGOUK/zF+bY9OKFyzgZaG0mh0A/32CZxfzyO8XeiiJL7O
cziadWDSZvUnET3qTEPfXvvBQ3VbKQBKloro+0iot4GbGpPir/nWyENl8FkYtLDNB3W6gHKzFFMW
RRUFA4V4ITPdI0ecIyzGsjPW74nZ7RDvfCG5HVTy+XkGzoqk27oJIbgjrDMa8xbW53VAiJfytRhu
pkRQBWSAFQvIiXSNCp3RyZ9O0hByL8Qkz5I9OYJzhaIawYIoKPgENas9kvUj0oQ5EwTGNix7J4m6
4w+MZNRGKjiB9pMrZlTv2A1Y2qdV3lRpXvG8ZTh/QIJsyykDFS34EOMwtv9YgE3Rbm8zHK6oyYhJ
6M3BuEBhfC+Axf2tBaQNccg/7nJsDAGWa/IpdD3q38IUXr8LZ/bfowRcNzxuAmh7Or7ITrKG2bWz
ZJJodZ48BHDwJxuvQf9N/TsEPURrHsaiFbGCr2cn4LN2cEFkXG+AjFH1tyBmKh3sLeGH5GBtPHXK
W18RkDQrcqMewlxZ+7d0ynPyapDxXcfT93UGXbJhK0iF6PAc9sVBGofubwKjabtOsX7zZj7EwAvm
k2s4jMIm2bXVXQVIGYNB/Q4Y70Uz1yjbPnRaiGbrz+NnclLxeayeJT4O8SmUIVna2/4NLjb8ZdzA
u+sFAiZh9S/xXz/+Ky6OT7SzxepUuECFhDtTMukOIgHpnACjIdBlMKqXD4ZAxODLK21cQ2Y6Qtau
hGqErhrNRiPVCOQiWBhBgFRy+bfCkPzqNP1I6do0aHflJg35y+ajavnWeZ6Q12vsUaLWCmV/tLYW
Ye/n9BbgN/fNRhgkp9v0ggv+wn+xDAvuPXLJQtPpkC3E2nmrIpRwKrSYivVFMv5T36fkGMb2tSqC
a7pI2R5Jygr9pWU0yplBYeIl0AY9m5G/DsximtXmPJS6YkFSybD/dvzuiB7R49zc59EgevyOdooY
mW9q2fKbEsGZ+DHGyKj9fXuR+rfebfua33JyCSvt98XebC4GsF9jE08+yx9qm9ey8Cqs+VB8Obyg
kawBR9y3m/LCs/5ZrCakIp6B3M9CdvYi0BEMC7ZJIFmPmfA2wqZMTgszKuvDjaiF76RTeZ8y/j+B
A8qkoEa7FhnCqQQ459vZBeLfO5lACQlu8lKhnx07QmiEuoHVYsxD5vrN4FpCGIo0FiurC1L5zU5E
TIeiONYw957TtN4DFFV69ZPsfPjTD1iVStAaMXKnBY1qJPv9/eeAqJ2oNLSywM8JRu6qH5aXEWZr
8iRH279l2Q8syIxgdis9xrD/YVXk9lxsLniT5e0F98JSl6mSczMjDuv/9FMO1XrMc0o19sT/rDE2
hYZjiu/SJDLcUTY7rF9vGW/3ioGE9mi6lMKbP3pISPI9M0bPqeTygvLvrXqkCJi2/muqnSd4jF0w
bVtVgaiGgwIQOJ0Fo0+LUEmEDJVfnCqMzNWtj+9ea4BJUjfQc74KPqs/9eu07v9gOV0oOIlrvux2
Kdv/tMy8zPsd3nRJ0Op6mz/1ADdPNhj7QhMSOXo8tXaPB2ioPUvBvq9vQx1K1HwXZcuDJHkqu+K0
tnA/R2+1PNMRe3AEBX4bqdjoE6dkf36C7Yv5MhKzV2BNFDDr87pzy0L2v6XFNfh8Fo5KmBu4QJLP
4GIaTdHsnlIpNh91JBYOWo7uVNRyVgctiyHQUcSP0CHJtyuCTdjWQd5Ge6xfhUZ44vci+1CWZDun
C5+tpHylhI2Qzb/7BtscVb9NbzQ5HjwYtQHTJcy1REW+tyE/r4wFbpiWSeAb3UL95hEGuMS0d9ZI
ddRNtl3cfe1L8FHlu6eSTUP7Z9FDvmyP/ZEQ9BSDdAOpdbXMqAVigbsRSRZ2QZCdWXjuFipGzmud
LEad+sYniz5v/kc2jKDcWAksGZMerHqaasa0kyr9At6MyfT2880pWs4NAM1SLj9jrBDnvvhv5w6x
ZZPZDf31utx6ZgFIx/61v86QRAU+D0bnSo3ODRQ6ORIJz5xbXHPGE7rmEyIOsXvGfAUUfGZ1QFl/
+gDa94gvB2+YSbA4cZfEMLgxCsvl4YLr9gmmHAuV9yEM4PDtYypR8+K6r65jFpYqO+Tosp1oNucX
iuI9lfQ9zDrC9btIptj3p8gOVQmiRUisrq1ql95xibdfS04a2Gb7rMNaa3nGPvW7T28hGknotRNk
qRotA0AePug1VRf1HgH4t0/msHXOEbGaOCNmrCNFfIZw0QnD47lsCEQXTsOWbT9Oe4mq7zLpeSyG
zje8egHkoEb1eH2HWLIaNVJ/zfUd6g2VWl8LrVM01E1ToBgp9LAu25tPZeD1l9xz/mD7/K4XBkdO
3VTkvnXCy8SBMPOdPn1eaALFg2/mLmCOPj4XIlH1yNjEL1bcrDOc7NQgZWSQVLvap1LvdwXRK8P5
93i04am1/qTFIkhALYOfmyfLzo/wMgHJxWJrrSJ/PzSrVS3ib7FMSd92iv/xAgVhafkv35Yhk3de
Vi5titmkXE0vc2Ph9dqC9qOnVn/711VD8J+6iSJZ0thC03noZ6wYGtHl4qcMMLdBSo0/omZFVOli
XCbm/cxbHk3X3KYPRhXBlU8Z+z80jDxDYLLfAzf2jrvGuWImEV99FGNpYhjiKTAJvTR+l9z97RpG
2wxppiWuOCrIXyzaAe1SZhI5nHAATdDr5TPpcWlpe8DGZEB7YeHELDixucM8NKeqaGKE0aBmfFTI
dWYPFDyGdYlc6pcZm6nU3d38oWnQz+mYqC20Dne7BlAfokz9LVdeCk4voDbngsCRPXPmaarmEy/k
kAyuSh4m3b5wvZhCae6oR2Wrv7ANRaO5J/A9XsovmO5G9gWomn+TqoSjV4gWKJbok55gTWHRM47o
d7X4osb43Luxmr36noPrHuwX5U4jRfP4k7ivpXcwq58z+9/PCPYFwloV3tkJYB3NVrhLbqENyF91
4CsoLkoIgesr8Lh41aGHIWOQZoKsZa47ScHnAhmdXAteq7cann9uZutXKxveDiNLlN+ug+l1Dn8F
6JHdttAwk8xu6tqBMGxaoQS0X5Ag7NHdZX0UOyC6xCxMCKMOt+KO8h6XWkpT8CNwGeoHgm/4R5Ep
7eO3gK2M6AA2yty7zU1wHFNAXGzxC3lNw6vBZ07JdL0jMU4nBgcT5rDHFI6HxW71B+WwYp+1MHJl
lW+bt8TASTzG8fVCp0fe5oBoOlXQB0K7EpQk41fsOaRfKSajrmhMKDZ/NhnRjDrApEcovaIzFvpb
6dIKjoZcz1ndPXGGTrLEy4yzdyN8EajxPqk7dpouQ1/JGUaRgQjLC+FHSb6nowG24ICVSdEHv++U
2UQscaH82lBbvNcHx9SnjLQshui2+8Nq2DHFeZ7LgxjMWz3PCSq0s5SBZcOxDzUZ+4vnIeaJIkdf
ZBqhE5Yxk1TaFz9mPXmofIrVrBptOZbjRYzSWvxnGHIcUs/zd502OugkmJappEXjxpszL5Hc2cbA
is5wepb1sZTCYD7qt9//XI/JAZ5NhDYfaw2VNupEpvJhTU5+qWYxTBTxpg5kI7mZAZ8GO6g64Llo
nbRrWl6ZNg2xacsbwSEMOGy3SoXiaBFMGuk75p1IHcex1RWsrf5nurhmUr+fn88ZyvIpge5Xt3wN
f8FSeMtN0APHiGVqoWxZtGBNmGpBdakAErl3jA0aGEa9hif4D1gHhr6KADJgpDvaP8vRrZVOy88m
OaVvwkN22lk9ouUQdhgPMJ+wX4dI/TRo+1csA37QeCYtz/L74zIkW4RiqsvL5E3xsreCuzpwWJSO
H6j7Ujq6YSB1JzjwC9GqUfVDc7VpCcjM9rOXIr1a9m/ccInR711uJqVJeCV9SJOrh7cVEvz96DEV
y5S6jPInFk4IDDRn7By6LSOgQWBvzUYZfwoX1/EwI1O0W8z6NO4jMlCzmizdhZF1/xFJ7jINiOcH
To2ku7k+drG8zNMAVlglQAJ7naqJXaTBaaP/pEt+9qEhVTVjgneqHvJ5msrG1+G7Zwo6tGfT9lVB
HujzC5BXra0Bw5gDfP/e3KEYtSZl5eDzqS9qp6pAyJg8PC6zJNO09xyxkmvnUptu9r2xd40s5jkT
E0R18RkmlncfBwrpn2JQF4cR/zsNzJgtpsUBJZmtGw0SR71u81Hj3CNjhh9dKq5K1M3jhy1B8Rsy
XaCTM6jt91eRAjDFRN0MEAAHyRrKQFnWrdo4sdhJO9X1PNZX1+wRU0FPy3rtgG5TLnCrRuzzq4sI
08E6FXjHpYRwdfJuPJD0pxWSyntxp8ks6ormPeeAkgeGbNW/rselPk61Qq3PMz7CLJb6yCBOlQ/W
j03axLMOIVWV4GAfdgGGsOW2RbIYFFsQVMqPsV76l78FxVOFIEJgKQ7Q+OwUe3RXHpX+UhGZac09
BWhL2+tUKUrMj/bo7HFRHwGZpqD/FqIrb6WwBv4ff0NgHVbRPfx/5Zs/PdiuO1NboCeD1bNBcY5X
0D8EWJH6nEAc87S7iYwMD5TNA+ComwPQiuhZM7pbXZOrJgPlZBoSfbZDrOEoX3b6FakmA1teLd6g
WjZxoXpCW4e1CDLsG4wMEy77sgC0Yt4XYR0UjeE862CDGxY0LuLqwFFL+vWBOMYUnAmaUmyqikEN
G4+TaJfsYjmn3BULv2F9eBoNSxfDCMuPTSlnfRey7JBsmNMrmeLC9faIJYXWMT7pe7lY7MFg9azA
SgfJp7gpmrRPJkUpWy2h+JhxG4fxdjgkmpRGYhrrFhWJBQ2VoHtXADONPry9GECS+JQgp4Ctfs8T
DkegK72ZJmAwCP26B0BxVSWJGTT7yeDiv5NRzj1rzWKQD3ZGlLUmWeXleIbgGw2kgAMIDORDNnVa
yDGKFVwDb2pJ38noodyZl8/2ZtNzciVXPJefDrHjeOJlIuwNgjYxRdzKaDUr0uFWRblTJHnqY8pJ
4ZvENOhADjJYFTDqMBvjKo8P43cJFVDlmcY+y9Yf6jjZt4EqZdSDuAvegcSYhepI3FkCEVFdc2NN
MkrtCcONNrk4YUf8jTWRm1s/s/g24ecf1QqEB3MMPAwD4B1LMTZLeCCiRqHR60t8A7TzyUpbU5j0
VMsUZnjRvOciXO31I2r3m/UWUAyUUs2sN/DQ405NK5M/Eh9CLECyO1BSvjb+RB6Y1F3lWMTR98JP
GVC4pET+AY9BmelqS473aD0ZoZBMuDHgFSe0KFgKO4JUIXIzk6s8f91cqpL5oTbVhhgg+SE9YTJy
mak5hxgi5pP2Ft9g4g+Cm5UC+/9AYnMyQ6cTV0DyL8Fi0rSdrl/T5k4wToImgqQJjOqwfLRQMLQU
fWm5Ajvh6xTk+49Fj482Pgcqn2v/8rh8rrESNgW58/0qYTFcoy6r63xE9ATX14kC/3+XT4/jRdD2
FeKuJW5GucyDoAv7if3CKXN2sN/c1fMmaEUAnnAcFQbf3pBV02PxqzMuPjmRA2x+zA0i7qclbhg6
z8FUTEF3w0unN25L+1dv/EfWIkvrXOd/0lT7i8u0S90UyxmVw1VdTXakuk5P2Kx3o6KwdpVZ1fa0
Hnhca51mCw8eF11P5O73yMV92hVpIYy12ao9oHjoEik7xZaCvzavrECVCH5v2dzH2+hzofAhhx2P
nm9wn9eaACtJNKva52D3p0GLf2sH5YRYdRzreRUM+D/5SyskQtqnD6IruDuxs2pBNy6LDIrh0su+
SUO+P+RFWU0jDBi/OSUvF+9V4je232OAmOR5gE4bMr0nYHtJtu22l/dtWeMZfItxOt3iGNesV9TK
o8T3BZoagVA8uH4U1OmGxqfQwRxAqLCQNzPAO7s/bh9bfiClaHAMcvfkgiCvAWeKxO6nu7FIUR+R
rDe8RYhSPyZJ7nsCgMO5lAGWc/zR4imdjddMrw1V76/d7p1gbmuS3zudOI8dVMBppv6pzmsBuHOl
ZDrFqy22NZ+RtmYZJbAzsZqsbLaQqE5vnkHBQswA1zncd7TcLdfqlwiK9ado9K8J8/n2wCKdBCuG
xOT7+K0ea0JmY9+1cKv0jQv1vgGgfUDJs0m1tbtSs1gjSgkFNT+8s02FSvaH+aaIGwDK+IGhbNIv
g7B3h5+wYF0qrT8QZnSX+sjWV8AY+hp1VLNn3CWR5RRb5+lBqLlhBs0goIjtj/IAuhS9HzMBtlvZ
+gYE22uKPMlwQ7oSQ0VY10Vn3hsCYufpetm/7rqGJEE/c3a3T328WXOtcQ5S5Y9QaS0xr+mAtESK
/XEnszo6lUxByQTYGr9vAAx36omoOv5h2kdrn7YY7rUTQVEm4bPHFy5MmvRQkNfz//9ggjXaI+hh
b8pzLOe8jm6Bn5tDXCWYPX2ZMRJ/flvbvhKiSAHhHfFhWWcobwKzqnhbXRtYceuM7QUqSgXxiUMw
L6xiGVrqNTSxFQAyJFLVEKeAT3pC4JMeJEVWyj4QsOW9uOD5l9cZR8TUpPH3ahTwVjoqKoG6NDrH
k5S+mFNwF1FkMviMapApXqZiV8s0pcHFhbsDO/x5/bjnr+1+9CxO7+xeEM3nh3Nk7OdCVVkkdTHp
HkMtXk817adY253VLCFuAReaOfDmY1z+Ps1rs9ojKeFOPm35C1+vxqqiR3cH0TihRhlrbucjEBix
ILiSZT21gxxzEBgDJrSiOn1KWIt3zg9n2Tsmliyz+zM3cIblGmhLQviet47m3quFNpdbPp70ITUu
KL/9mM2mO+CVQgHvs5jUxBE61WVVt2gc6P+XEXneRCXuuileV5XMnaVIutPZwOE9IuSiKm8OVM7r
AXOQSfoG+N7cZE4vdE9Slj4626UiCjxej/F2qB1fMhwkbw3GRGyS0J5oOwQHBmImlT7beY7WXh7I
MxHXwr2UWk+6llPYLghI8YAtfSRSjJcqubkEqX70Pl1zL2Rh8TRZWIW8ut0Z9U8A5GvHzX5YWGOB
tU5WHUxIZk29QjXX+IbFJ2bcTzcu0I1cOKZv6fF3e4Aa0YSzxFQiblL043QvMwdxJkpqCR5917Wx
GMS1Ud2UX72SotB/Nj5H6XeFwjqz385Jx1xtJmYpMWVW3POJZTWQowadkgL15a8GeWFL9VNH4Hjt
BemUTiGKZ8H0Z7n2Yq8+GlO7mdUi0d3UxRty0RxILyAyB6ikNxaH2gJFfe2cpyiI+w7P4rkFjMao
iJpB1lMA57JZhgEIySaog1kMaDibSJljuGIehxU9pdlzj2jQ9vhGEKE7yQqPd4hRxMrH0k7gHasI
uJq63toI9Pp19FKuHd3TQYVk9nlLWIQKxPoKpEfWysomxbZ+8R0y42WfSA/7gt7C0kytgFNKwMXM
6XoLam71QdEgVAdbunbWdSjdBKcCntosfz+Cv7VFA36E8gv659PLY8Ej9psSPcx1m6fzhIxC0ayt
Pb+zJBYHEX6nfWEG0ZCAkLywUuWZwRsm9ip5WXyWHQiuZuJTRmr048m+meuRFrA6LUyAatHa6qbB
DQnP5c582vWoe3eXWnOGzH7BbRKvfyhD6ic2R0HuJGCA+iuQGEOtmpv61C+KlwdrZDDjBk/xlZn3
Q9CQcU7m7tFYQq4pS03Lc+B2YEDlTPqRnhw8py8Y2gfV/aoC9uW010J3zBOwVmbX83RamPBbTn9h
C3a639pNBJ2dKnbNHqqYlJxXEVrOLMQ6ZsKlTmmOVyhddPoekr1DVSNWWp+F8jFSaQDaj1sGjuhz
u0rzo+arrYGjdDPPuylkZe19ewu82T9vuMyVoDo/iyEelUody9muF2GcCmQAAFmd7vE8IZn7p9Re
WrNPZQKm8gIZO7tzrwluz90JieItcAqMot5redUCPjwXuuovcJ5n494bX31z5TZYWV6V/HrWHzYs
E5d9nl/BauoG4ssCvr8GE9TEV3GhEhUaBzSn8EyD41+rd2B9dOGGITCrcnpAVEShPXXidJUAs5/H
nh8pBMMVu2HNB1le1v8mrbksYa+wzXEOr4yeHjyEvqcljW6n5DFN5rmX9Q79GA3QNJpVq84zuvjc
svBvtA50l/enrFFBhtKCzUtyE+TrTVW5MWzF7N2R9WF3GetpX/3jGHy6LrgUJvvOE5YeS1LmDpgo
F1GFMB3CKI1cuu7fEXSGQwE/J2q9eTrbp28a6cwQMLZ0f1wuW4apNovvGhaWH/KvTQrqwH6174gq
0ggqMDlglezssnhpybjpQDQVmNrj4YWTtzkQCvyid1B76aUNLT1jY2i9/GGEGEtjCGp0rPjAjwIb
+W3bFzze97XoBovFAkdz1yql8lkhoHMCvYyi5PFlqmY9OgyB9XBu1PtLrBfzVZMcLvZc5wkxT1aS
98vwFA+goIwdUdpMYwPiZVPfjgG2dbZDjXa5vYxXaduwG7b7KD2pbzBKN8jL7ST2GYuwCqwEDkJn
4CBZEXrPxZq2K9sZ4OcD948Aq5iAdeGIlRp8L1RHimdks9ST/haidbkRr3ckjb8ZbFE95jhx6RgS
Z4t280M0s4sYoNX/YUkg31EZXsv3xg4OrQ5b1nQ5sTmsUWb3VDKZMq21DLhvTLZ446taDBo4e2wY
Ks8f/uXxNEWyWLboH0H83NtsmDo1RGVDltwl29x/VLZEBuQvaQ1epPWbfFm41x+Vz6uueNG/wKCe
OIokqUaYd/ZMMl21iOzYsOkqyCozJxIBJYILARQIo8YV1AwB7R/3zsDh9cyErpOD9UmeSiylc9Fl
5PUxM5Mwp31WdRdbaGxUH23bnmN6A8owT0QK+5XaiMXAUV8eka+hL/RjKp5GwbHnX2t4RLAPg2LM
cptnPldRWFat+24k3CJSVJGmFl14hmoU2FnvB8U+Vbx3H3sRFZK6UKGoy5ogiknl2ERNZobsUJ2G
r+82gg346BaeUcDp68cRcQy63bMmf78Ubkm3k16nZqRyGQLONcmq+QvdjmI/eBXwrGYFJtQxLCvJ
TAgdrdYr2nxmQGpkb1+ufQ0jNIRF0eVgGI4LwaEjB/9Ndd4VnBI8urUHIjTgIqGWNA3TlHARYlK5
Jsg5VbrY+W5mjiV8Y1bk4//O4cHS05QkDu2O1ztuwG1oEjXZFogP6uqLSXKCQhtfoxsbvK+nPE/a
/7O4sDvh6+37u8yibewgIp2fd97cXB9E1WxaTBrNniuUSAhiwN6eAI3ysdV9qgLDwu8Wr/Xfm2B1
UYURO3olSnGwJIkg1WnFyIIEQG/Ydr0r/xYRQ8FwFtyGx2gl2iLMdmQi9OAxzPUHEu9VdoEh2s/Y
GxZyydzXG+ZiP26YS9KUcHjJV3ImVcxW7KzHNpqnP8+q8Ae/xFoO2zcKAguUqithERFD8VFyyj4c
fuDqwZt5Qptgad7ZLmnnDQFYoVztxIbkJQZIYE9vT8B67xeKhWbc+VmiPaOOxjpevUtdu0TRgHYI
5toNvAPvyG5hXRQ79UAtYduYFhSenAnxW1v2DB9XlojbxR2bNLrVqfOfqMWH/+1ZncOv8JodJK4K
BaUETNw/GDo2/9t4cyvTQOHYSPrJuHSBz+7ezMviemIWvhv3fmrXDg+88i/s/I6D43AhcBpd47RX
S0YXAIM+ORd9CDHKpjy1AkM6cpYpAPb5/Adbgw8thr5JnhGsSHyDlSfsov/nqzE7YKuZ2xcjL2dQ
GWP/98EOm8e7Z2p2uZ8LKTAT/QSS5ONJ8MnMByCZ+DrUnxTy47TrMtqD8G2cURe1uhNQxHRlEQis
m0i0G6v/nDDbSCYiKwRo+ZkbH5EIGQxenAO/XgHEMdCIQLDotHnYQCC9GydBjeiXhmxIatrlaOvc
ABh8TaZta85DQwxb6AgFucJy9GmM54uXUruOCkwGLP07KttNOcoUeSsiDk4Mz7bzCaREg/Ay560f
Vzw9lBZxYkmkRIZxi8uTcgTxHKapanmxkCP6zyN1sDv/w3nrSyPIvlfvNalcdQgzStLYYXRUv7p1
vBdQR+2JMaPjleOvvv6ottN2lAhLfhs4OuaSa1kxhJKzztgWUusil9EoxTqz3drf2uuGkDmr1MlL
DNYlfIix6x0Gp/cAwuNb+bye9bz++j+E7oerDhKvWgPjIzAzsQcF0n8ALdMSdQUr46p4OFUmY3RD
o8nYQOB+ICGlWqk6oXDbemoGop691zJ7crXp/roKGvMgiAVlgU58BnQVb7YDfGv41O6Aw+ofSZrd
bAQmV+owJUOv/LdaRYEtyImaFaWW9BJjJydLUUsm/9tcaFbAQUvYJzJOa79E3oCxItD3GmFNdXEK
rDVNK1SGjjV7L4naYv3BPOEkxOG7aIXgG5Kr4mwKpiPJ8Lg0JQqVB3fm8tuNSkPlXVo5dvdqu7D5
3RZsJr/6B3J+t3jTINW7qVniR9YN2djUwRpeZ+DugDySsdttmdKM9VevGJ85Syw/68sFVcs/F4rx
XsGsj3WMzZ9KfYjqX87Tvj1cDYyM5CL0/QJL5XaOsZNcWIV6O5LYpZBYjnGeWSUzWc/JJZotLNuO
ez3fEcxzfucQZpCOu2q/yIrRbjJ5pA7ZoYByCNdYvviDf/Xauz+ILEA05wYljPCrZtaNCrU/rqU2
spmioMGf5vKuDAQQXFOzBUDZiRKij8PdjZqRTT1d00KFw3ybcQ0yh2Debi22JnJlLad89ID0L10c
4NldzGthkYI/Vg+9K5ESHzbDW3SLw/py6YDQJ/r7UPnHUoL+2aLxYJyKBq+4od6bl8xPfnqXJcal
9kMSLdhlQF/QOef6CClM7dNWrN5EodLa8PlsrDX8h6D0Krz2+Ys68V0vJm/GyAnUatl3uieXPVh/
cq2mNRgAA1cyyGxydzDT5KlK8t7LcqglqUM/BzzFPpAIsdV0bY7Gd28RGeeVCnOQbZ4taIRut8tK
4wgg6X4HgENIPSb3l5rHqMeN7iaysdo/4j7xw7wuntZxyVex+/kdZe/BipBqyB4ygFIK9YNIjJz5
1V0dBTrrdkXwBHSq6uwK1w+r2s/i/uYreaPCt+s5OnERhqzbwNzBBSLHXaKp+wwUrToub/7QWmGZ
vfAzbuoBUFO4gdOT2t5FwcLd7S8JUZwGHrPPe2WqWI/qg9JwBBzBj6G1mij2bNHoLR3XkZSogwSR
v2ZnFhY180xPKBqpGOTMMW7cc4bXNKyCIuDE9l4OswRSBuTGBIvFMQRGYcZSqG7krAPwbuUqAkbY
NjCOyNVgDnhtekwHjwWT9M10GxB7qswBq/MGTIHr9WFT7awO3RCuvEbodOSSjMkXOQXYHvZZzjbE
ezfOq3DuEURjFK0i25JsLFVmPdu6oRouCnK6+92ksI883/otrz5JbEMKgaIT374Jl5zUyUVO0mu5
cJCK09/Q7Nq9jPuGIwSeqDT6WIMF6Lxz/Unu2iIz6YPH1NtX082lfevgRWYIfgULdG4qAyS1TsTU
6O2a4AmJtaZZ0vIyVECve8SDgE8IdU/wabzdzoGYxNfgDG4AvGULT5Fqo9DkM/oIBItdhefBEFkf
G4MIr6Z/vAiUJ2AHlLjOrmA60xDs/t1PN4qI2titqi4xuckqeUIgI40ycWELQDsGt9SLG9lDFZld
D2e9MCET6agokQ8cFTpm7QK63QtP8pwG4BZHtXxpEMLH3Lqq/y06QFNbrWIsQNVD+iORxYSfeNkx
4RZTZ5xYaF/L1lPFT0X3as0983lmfhC5XxcetukDLqLdVl6eTmZOGaRO3tOgYqRuRGxlPsTqed3h
0Kv/65k6yWjTScdJFG4g0SGcQObVjKIs0F8ULXOoNmVmoSN+JRvHlcVwxdxga7TOv1dWMcUtdO/h
liIABW//CflPG5szrZwTmukDi5n2tyrQKadAnDsK+NSDRKnoGH5ES2UrWntcyw9INdSLgWzTmDGv
bpqnnrLvppA77OoXxuKaFGcw9J9/h1vGUe+6qIGrsYWB+jv8BcocHRfODFlX98Gi2rvshWjQkJxP
aGJBHY2ZSUe+HY3luNyhTB4IJL+zysiiQzLV9mJH4XART2/4oHYn6nVMpBq6La2UUEEN5fIqCJEK
HliNrHExJ1y6U4qhMAeH4YWZ6FRNMVFc/NIGuRiJ/YQrKea7A68g0DvhZgxptRK0TKZVygNoXs5E
FchY8RDwPN3lmM3ZKR3Mnjfb/2ch1HbaYxtYZhRwRaeDZAs2hErluDcVJ5XXpETee7LO1b+33hz9
3hbWeVIW3ERmi26975ad9kaZUj30J9B54ZxuCkH6FMRM1r73nKY2df6mr3Cj+fL/rQlC2NqYJv4Z
P7cNtL7JscGplfnOY1IEbl/3TBgHskrP8loA6BI0iG2BYN7weQMLtckSBp1ooMAvmKvmdxfrnSRU
r9KzTlLvSb/Tbt4iKgLVv4ALKHO7WdMxqXiixvYTxoa4Fwo5xjbZ6TOGvJSDSIT02jHYuFd8nL0n
nJxP2LmGdpzmG2bjpvFZz/bUpkq1lXiaRsbZn4XjkQ3VG5ptfg5yUInqWBGDzujg6jD7xIQC5Ns+
zqVDwgBNlUoxUWKo4iQ2Me0iZSVnEQl5fPN8GqDnLFMBWfNWG72T15j/hQMXJrjaQYzRXqRlxDFd
VP43yG3ZVKi3ICFqTSj+shgVN8m2sYHybDmh7xU/crR+n3EXEGD83b8K9tT3V/K/W6C186o9IrNf
4jQEjuv1NbrAgx7ih9k3cWt4ogUc9UtPka/GQqeTGDZgvsYn9ZX+AiRjEgXc9tId/1YCRXIUWbJ4
so8Yi6AbxstsFO7JZHqY4BihNddu0RKGB9jb9KHPaBkh7RPQDe9lx6pO0XrAbL8YvXD1C00fnLEz
aAameNbSgQBTBCdwVEzo7XPxu6eaue27rnw8mKicqXM0QEgWCxBLuWh7Ck/MgIYxpqHVMNpfTBJC
w/8X00Zprq7GeHN2vlCQKJAbaKaIowLR/Pb28LzrKwi55Ph5xooeP9eEeDGYGo6cYeXsI3B3bTGZ
sUGy3cO0bdJ3nirtkrrSlsJ5QRZIxY6/al/kSg5RawkyyfyQTLFV52BlEh1C8EA9AlkhKD2SqDDZ
izXEq5hCutjkqSrsJzFngYmYlkmoYbrT28t157cl0ilV03Zk5Tg8HduhckOVIqlMoJi9xWFjHJko
UqY4OK9hSvljWexRXwXVMRsUD2hAmRXC0QkwgPqX0OGpaekVHEC9cEa5tVmXdJ3Tl8a9NmboVUyu
G/HlUx5LIi9cS7EM2XVQ2sGuXIfFnsgmUGLLteNefRLxzORgrMOrLidNwxfvODM2D7xeZaQ6eXXE
Yma06r4m/gqGYDox4ukbQYBE2eblt1vqgrDYWR/IxCEsnWgc3eDs3Ai2HUmoDWQmRTjmGYEJJhf7
amNcRn1qPyjkvXa/sorfxi6YMxeC5VBQDlFYH0nVO/DmsdBZPQUXAypdrfW/pV6Q7QMgW29zTGbU
UUb1vNuV4c9dNKb27AOqO0tS/AaX+j+178O5s6oQ1q1qQf0R5I22baFaml4PLZamqg9osuUCdt2m
CtW2d4lhmxecF+RRxSBm2lK104NmsGvSwzHCIYJIxCFtDYSMNjEP6J1qPnjXfGe7KSQYEE/kGchH
NXKF77/J97yEKXN4f40KV8H9Dtdq0PIg0diVjNAZgkNDWR8t8gCGsXX6Nr03Gp3c0NV4lBO5NU09
RthYl2nexmm5N4TiIMDISphedrkVahE7ZFAvnwFfO1NDeIJB3E/3XFV4UjSM4gSYyE88OfZECXXq
IHsXBBNsfJck1MJNowUFOlkDlCsjGFLL6qIAS4O9F+yJBU1mFwH3/o/7WgTDg6Wsi9Mw+5SaM6eu
64NcpnMBhAhdXuOUfIP5EwUpbO2UV+E2AgCzmMN38bw1Ne4d18y/tV+UiybTht8spKZ8gDfjOXfF
0nUo5/MvtGbwo2osAT1zlAXmVJn1Vx/9TzYMxRrSl+LEeGRZhvYyUqmGn7nmq8/RBlIBNhHQAJb9
tdW618tY82CCpbqCQ0/UK1/TrtTnNvTtdD2jK9upYAZ1X/2S7aEKUF8Qf3JrYkKPFmUdpv5AhtYH
cOztHoWJsG2vqKRRb9D6fOj5bVU0HSKj9nYGlmYt62BjRLm1N9dd0M8/+Qq9u8+cUYj1VwIel0XA
i6+mgcET3FJ9cTKUB0tlog5UHK7mUUoYQOHcx0KCcVzvxF9Ypg7MlLK7nclgW21OkrCA+4AWepGT
Q3/vKydO14+2D48TkCbkOI0GtM1LFsn7QNw/PDaeImte9E5I3RlUEzvWT9DHcv76LjeOfgX2BRIF
9QJus97+QB0aAm9JUjeBEWXFr5qV5DFwPF3HdRINzULAWgMz2Oaqa/Ny3o0jjiqV0WErBos+YmMX
Zdlr5XfEq16Cd9oDALfrqb2hJxmY4/kDznwuSdGQNlR3M9trm87gNRpn+E8+IesgEiQ7JFcsqcO+
9w+vI5lsP8SS6aUeRtyHEAMAUN+s9lANuWhrPjRfkzs/U7WfXBDryXWsz+0v5m7ahdkfk8HIn3Kh
4S+1iIN/MemJzlQOLIWwmsWqJYZnxleoY+ssr1cqbv3QMY90OBYfu1q5sCNSH88z0mmqciUHuGpb
4j8gUbIdU6+wMdq4s72mKZBKnEuzPyuS8RYeTikCaiUEXV+bhKoPDLDPSd7ZkO6oPSSa0TMeciKV
ElcpDXjSI5C5KX0mJEEfTGD2N7jwcLEPUJyVl101vx/0UfNFPfyvfdKzvTEqw30521hz84pf7ZvW
YSW7jU+AOMwB6NOyjEI0ZpYMBbNwPhep+tZPB90uimJxIl6eznc4t5+l4GfKtJRMjbfDDb7fqP7l
LVkQuRDZWXZaQDJrkaufmUqghLC5ygvt4yzM8HczxlM/QcR3+9g3m21iGo3HE6qHBq7dRXnXpyec
9zxFWKAqlPkU0TBC9rndHQJfVAwqIT1oN6rhU1pyIswM183n5EAtd158UzrR8gR+ZEshySsfFTYJ
lr9qX2soFHgeILYKgy5MSxvHOhfwfmYX9+mHvg2iXmsXq1Avqu/8fiovO2VYbBe9tYce/VxNs/Km
55bCRpR3YoeEDateF1vPN30f79A0kBHaIhqlM6lDl+cqcuKZEbHsmsLYD7dGQ+s6JA7NRErdbh3L
xcbKjOfXf9TLXmL69D7qHrRkjBXB6qhTXwF52KkcDfMhfYbtN1VQn7VqXpR+LP9dxWAg/mkM6f8f
ukmoZ7x5Er/AJsHBQOHgnbNYnaF7166js2maKtZKNkY2/xvj8fRfOeBcphkTGFgbeC6RRNYYKr0w
6ht5Hh5JXIY90jov3RsWFPOESuFKEP5Z2PQ4OdcOK2lcfs8SG9mAQh4gHr9U1mrymUxW9hFFD/Hg
ynfQZtxYUkHzDsp1lMHAEjid4Vny57gQbsLl11i3Jvbs5/LMZEwqCLnN0xCwNQoyXp4svxgIV6Rv
36ASwoD6+tF1wooRX6ptttzF/1B3i2NmS3NKT2+kaX874lW7zLqrtkO5vU/yqRfev+hXmqmGzX23
2ApxXs7EaANxsqLE9YqERgUXO9FRyab1p8mrMVP6tw23zRVpYjasUxykjhywB1W/qVXkQY7mMoln
NpWW8qgD0yTuc/Vr0kw4HmoOezng3c7vRaWCWtowIhI8BnYjc171KJQlaN19ey5/C9Z92cwLw32o
ljqdSGP4erjh26rD53wMu3JA01HHTXVr3e2Y6Rj1Kj3ISFGuB45TsFcsRhM69t9GmgytyZwFV08N
kWyhiMnJskn69rAFgxZAJn4NcWSnKsEc8ULYsKKFhBMsi0C1QVLiXahV1W06tgHg+U1cZIQo8fX6
QN8hLA0lpKfl1L/NETSKbhy2/b6t7l/URw/88TwcE6Ef2jXtZzWsGNwjyD9l//tyFzuuUAt8Wqop
z99P2/NtGmx0P5oB88CaJ9hYyldaXZCJ4yvYq7w5rnJhdILTCmZIEuogebmg1MNfbhJj0sYEpbFx
fiNIwQ8ujewQtr7d/T72zjUJ61llvg1KkTjzYfHRqy2cIRFP91/2oKjfyWWwEdGYclBLayDpLd7C
KF8KHi5WkmJJzxdjzjYlueMWzLMPxrVz+wMqp5y6e2QPqFnmfp0tqgvj49KiUGJ1Sb8C96rJA0YL
2vSJGXPmmo82gm4hig4MOfEujPPUM6ltqcTIvbGyTOumKD/yKKiZyA0OBpKqoK8UeXphNrMKLmps
sS6AEzOjchJC5lu2S1Lo+y+VdwEm3xZNVAKUAAj73gc+Q6b0XcMxeyFWkhPP8kqZmjBaR9wOKy9f
qJyEpgjcuEdt8SxDhCAUO4M+Z9G4+YHm8bLD8anFWj+qFXbsI8arjGPuFfj7ZRANhUU3b3HsQ6dC
4Y3CPm4CbfX9HIm4Hx8MZMs/TK0R4fV0TkDVwJIEMrZCXmJXj512XBBa5SC44R9lozva26k6gyZt
5rkzyrEIjvR8vlq2YqN4lsi3BR3Ib/K4T6ntpEqpo8NQBX5ONgpxoS90c329N+M1kx5xPEgCbp8y
M3c1Dk0JxCHnENnCVBQXLmMOSSLwYmVW7g2NSGebwcxuVnWL6q5ScouVMG9VO4wuldmVqGsd2o+v
ofk5uVjS8RBbOGID/+54zRKUPx9nFFCwcS+V01xwZuCx+fx7wpq6jZ2g/4wEF0VRZDmbbDloU/ru
orLeY8v2SwDfavdzz0W0CV4PQj99cPJ7Q+x24yyrYGDcLkrP0LXIYcKM1J6Ho0a9f+wc+FWNLZQU
sqQSmq9Vt+srPMIKfYTZj/wDwCMIZ/yJS7kASeKzSMZ33264vi9X3TrRzB8kWKTmc7GrnVfAP+Az
yrULc0GitjGKJ7obTwMJ0elcf1fCGoEw/GjQlMx098uN0RfuwMxBdsefHDEcnzVJNGOcdY+F0yMv
YQjgp37alObQJrvJE/+VXfZtTJnTRuExwuwCiKUlvc0TrtlZbKuBvlpd/jTOU9hJT3nL0rovUOoP
3PtMM2IiFquKwtyNKptCXOyINEBOp22hBXyC2OYRMjhXz9LKU2gpH/J9eLJdp2vYkyf53clmvdiJ
nbiwM8A/rKdwyajcFSlHg5erhdBrDZDApohud80DbJGINdc9euk8P748sE32bvOs8XsVLEWydmj4
C5eYV/3EbpUDNalbqGv/Nbj4ZmAvP6kaMLK5QsuTMKIXsPv3jshyOLAYAK7a3MeIqRw3eymRMpIP
FLAX1hS38sKjui2U4iE8kbUaSFZ+yd6XkOfkYNa+moiN7EqShvSF3goB+9mULZRS7euO6KeZDy68
5KatuJduCUGW5x/VjtSBqxlOw23/fiHPatRVnjzDMsWkEllM0kzMg9SL/6VMTSke668aAvZubDsl
kK77ZMC1JbhT3nGhpyihkWmaN/0AjseEDqbGDYsXYTTInYh2z69coZ+5gPRa/xJMiEFpXKGC4zEB
y/MsxtUTyEVh++XPB/BN2ol9OlAHC5FLca+OrbnwNzMZPcBzogbX8b4is5EMit2UZ17yI+6bwHdn
aRnTpZuO6236aUsIWfyQEbL63ywwZ4NsOGDjIIlxi/2paMcHSy/gdapbvfFZv6f+T8+343io4Fjb
xZwnTzgdaWQ/ceLSo9ACBhe16QAcdsQgyUZG+mhpFZu178j7dkB9gccS1zjsVl4W55omo2l89rTm
L5bCR2FesCVhsnmpOYsRbfotCSh37cqcyqcVaAoG7oZyAHuvNFlw4vnYLeoTqaaCiiLRrNWE96FE
kHbWSyJRqJayVjK6DmwXeDyEepE7dFu65IvYOoAMClSqBOFrfatU4QX0sPqFBNeArEipZbnQ8ClC
Fdk/7Sy0DrvEc2MryY+rEOC6M3kHXIAbRDu3U7CmTRP4u67UA6jMLh4ypf04Hm85CEKxyPx2Cl33
ue4JNdumdrk5qMC3v5Zw1arDXpXU0kpKSmGlmLVuzupqbhNbAVT8/CA1Kq1nffdJxJ77lYGGyVkP
kHks43oJcZMjZGkf+NsZv+VYKQW64qnLn/ZPZ8Qc6shwLO70hSnJJpqw54jFNyczcDST1MLaoNgu
02A699lOSK9URy0upe/XA6BI/1sz9y8MnUJoUghnp3hAF6897Ql/8HabcpIRynh1++M1aNFI4NG3
DJZQGlqWZHjUDz2vcuqKItWhTk9SK5uDp/ATQ49QB7fF88ce5h202Y76JLARaib1WF87gtVJbGAW
ahLrF+RRvw5i+E+VCEqkeuDgA4q3Sx1eJIh76ulmMlxCX2HZnEA3Z43OfU+pxk7X8VUSZ2TIVx/K
9RxfH3ssFfPrmLGQR7CLe/ssL9kAZghxFVRlfwnVVJX9Z98qSe4gPN1VZFILUXK5UVX9etXIJ4ax
OOdYIdYyRZZmxZDgC2n+Q0BIpiSkpoM7vY8YaGpC8r3gIBPhruiwfOq/vxkSrpLd1tIiz6PzAUjd
fNkYu9suzB5CEVLeB9lXD6g6rRilPm/JwKocmmiX0Zs47fZzkMn9EliUW82YXTCa6u1TTxwOb/Me
tNn2J0WuhfCJ+lFl/Kq6R2zCrWVq1/wctkIsR4h3+xD7vXppZ6BSPkge/WQ1hz9odGHdlon5Pk0G
Iyz7mZKATJCpCER2v1Hb5z8uPrGE6vhl1Nvo9SPUIy+0rXaeszdkA35+CO3LlJtC4p9cg6q9jNlJ
4DiYVfysRpkxzk8nCMh8gHBkuSaFBr4y+ArZ/XJtGWk0IijM+CSW6HhwKGhZUT2r4thliHJ9MEhx
03LuAchU9//Q1F5FMJTdo9cCtcoMNmRiYje9hMug8Vpw3wZUXUYS2OW/JYbNzFQpOvJSEvbfew/C
ZQJYXssSTg0BC2II/fH9ZcYlDP9pb216FLflJLCCFEhM3l9D2762YI/UA3MmMPTHIdnfz2Wsdln2
VlGZiX/rRpJbkGnoEDSBftV2ruL8GdJu7PQQjsqowrUzQAl2EAuPJomIwID/fWXawJWQaBZB6YEO
XKe5oZWGxclBJgZnrFEOOYuB3OTiRFg62q2hAGUSTwel8ngQtoCh5hnUTDWEvXnwjXe4v4XpQwEm
eXlSaPwrV7bqsCSStrFlwxQPl/kQ3igQqFOP8UDhlFoK8EyB8zaT0lrWUWugpvRw0fH6dVJxNDs3
YA2slbibHLSnG1GTpTrayON+bb8Z36W2W6YWaVQEnKKKPbKErPzV5PZvVRkAi6iAd/XV0iCtoKWE
G0h33BvXerHCfUZxZt4dkVeJYuaEsUHZilan8IU8x2I7qM30eafZO0cp4mLe5mPCKMvUxQug+Rs0
p/yBylGZzVDd9BrSoaCh16yDMI7Ovn6UJ+rHc01T7rgU/PLv2xcxMX/yIdjYsU/YBEVWljqmnQIn
hSqtgIiTsofw1wBTU/NCrkEmbFKA9F7YsqoZ1iJ0Yox1T2QA/zPDfqUSXEZeLqNJMcfYl35/TydP
heZklTz41wP/UkkMnfjy1TZpb/ZtBBI0FdMHHUE35D9VSDDsaWp0l2TnEpRdxlAfGbBgI/o5xhPu
8NTf5unzVTFRI2ftWaDp4F4Ubzay2X1xtCy4YJUH+if03ANnoDPg5graZ8a4Bke5aAAyZ+qJ1wfK
gSHkNqyhyJpRkzGOK7TLT5Q8Ig6mx5GMqGfG3MLQh304ldpLT5u84+T2FAnid9F3j5LGf9opEq1G
G4esqbE528fKArDq4E92AiyJWrvAh1a4xDwsi9aloWEzei0WRodMOWWrReTMvqbZLXa58W46cKFw
2wuaaLmzxWn0ZDkGwCzzfqutanu+4esknaM0Zd8tmTh6yaNc4JNNsOFWjWA6gHfPnmsfIFGgjPA1
U5V8oTDBMSW56htmhueb2zCDdRLN/APTK4wC7ROHSXhzPJqawB65DooxiA27MfH7ntfSMPhkIrO0
ZJczKeqQLmXVW/+cmnFd2m7DTF/dE+Y3V9PCdEBAgOThGUrayM7ajRM0uO/pSTkbD7EOLuspu90N
FAkCWhnilBXUFZbY0M8S9GS3Pa/wK8wAd9bm6tebdBPNDnP/xbPjzZTnmtG0QLoV0LPCOw7CYxMD
PzWkuFUuPaq4P5RiGC1Iln3I+1dnjizGOADPSxhQDtOvB5BKHxerKVE2QypReWnqpjmiZ+qVvPPu
v/Rj1TQjVnf2dg2RzL0Qm7uYXz9GO04PAgNrp2woAHiFX37s1O8zKY1qvQbWmA+JASdDJ1dDT+9v
LCJGrYgoID7VtSClibs5EfAESRWb9qXbG6xXp48wgrlHPd+QZepRlBtbkBB1U8CiPLfAYyLnbGHi
e2XJ9I/WSnLuXrHWL3YT9O4qlsk/jT2hR5Sr1LVcC/wyiggmWEn4jgfvmbTiDvPH9InzrDI7Meg5
hBZJtGIt6AY2Z12CRTrM4Favf/11RSJ1wbP3v2iOCmOV+JRIrh14oBz4KskLxrA3Wpz6qU8Uf/T4
QmXhcgNsdqyxnQqa4ISxFbLFosCChpLy7HA+lc04gqwUKOchphW46RcPLOKO2PLjKntdIIz2F8Yn
TteC4HP9oSob9FvFuSZFl+gGc7hDSd+SyERKZmnQO/ZiM19MtqKSyCnUBp0aTrxJQEhds2IhVs70
BJKqe+X0BIrUFfQRrH6MCelLJodo0AgY4etEJSd25g2BY05DpHo4OG19nG5xaFW3b40NG1xH+bmi
LHVlX3gLNl5gfYt7vyMWa7cIru0FmG7zGIQb1tHNjHzDnX4J9UWLn3mPe3xnBnD8pPMk7dKyGopw
E6bPYLaKs3slmTZ/Q6bkz8R4OLrT/pd7MnboRif/ZI+gm6zQXNt90ExXA6NgFuRIiPSQ3mibdhn0
h1VNN9jyMfHORC6LD5TYcXLOorTxX9FaLpTD0qn2RELvjIt6kzNoY7g36+5kGxQopXx6sTTmrlk2
u0UkYmmM3sOuDFcmOEYnMdQFLOBD1qXDEPSElfDZn84+5ClgIRmZC5Mct4hltnOj4GEqNHM6qOlO
oToil3CvpXRusEauprTWX/GcgScV/NpsH57+EUbNuxmHCYHK1qYvRsZFssADOb81dDruklNSonAV
sx4LyAZMsSsgYZIyVlngscviII4oqeVfORCEoJ0/GpaSLMfY9N/RfOFVEr5ZCD2cfPirqytjHgZH
AdKtvkn/rfGpae31h3JYLxXkY1chyIfbvx6FmD7yb20x1ZawG4QhcukvBiZU1GyJDN2/9Rk3hoQV
c2S5AOPnegs1G5N5mOXCIgsruUDHgjR7w3TCvJtLhF38LRPNjeuSaX4diaRzwfpRivCxtqu06Evk
/8V9KAYjDW9Qw5cA7yygloxe8r2Mp+5nE3/fLkz5n8CmhwxaU8yULHMqWNDNcZ670Y21XtuHHz0K
2I2YRNlA97LyVEALmRCSeQKKoi4+t58f0/hqGL5yoliR00shObcPf3TGbPuCfCLHdptY2nSPyt0t
mPtf9xoVTOpwhtLDLbJA4FJVy1hRoA8s8UPFDT4tr7Jqoydi1EBORJMnoErm6HZVeOxtVJ0fdqy0
nWGt+cA43SuyzogxC1pTyc/bwFxKpYVlOiZ+PRPgnG8EHu0PLJUwtMUwESDwxgBoxrJJezv4oHko
xMk/GU8m3LiMj/2GZwr1ZJA3YI6VfRrwoSgVXIFpZs2oIW+wVXCovu+BSzzU2QDrE1ZRtX6gn7So
gBKsLxinghkAyHm7uHT61cdEiGN6QTuh3D3QU4w+uymV9nLxizX5nGXzVOwrnlaxVfj95vVsELpK
zJP/cplnSkHOo5/9aoFpN2qN4RAr3iJzhpytnXZl3SNokrnQ2Iy0OkEXKr57nscoiHlrNLDZ0ZT0
bcB08ZNB4i+BDbEWmNu0LpYSATcs9NZAgd7YgTarBBXuLQ8LLPAEp/H8rY0AoUh6PI8GwdL3z7PZ
BKoHxGAYZZtPQk4bGwqgaobtCiCY0/cgCwYbPGB8AeQZimW9yAQj3WfudztBZ7UpYYeLzpqQ0ZzT
xtx3aesV6fq6Y1UBs9ZG1W/xCa+VruyxL44SC4LTmWyy8/2967+LSrrUbH11rjX7c00OSCl07kV1
mT/7eqnT5jQUo6KHmF3WtI9riIrHhzq6myXV4+2aWSjP6djd6cetEE3yh1CQx5PwUosPC2y8QjBe
bsbH+GTVheDr/Ry0HzjEs6yYnOJv5eK658duA589fBFP74lworvAXyrfC56TIkbgDhzJmNze9Azq
j4V+nVm6MnA9gwlJTkd0w6GiGTOmpQJ8694jraFMR5Fe/7S9zzO0CAMe4hKS8Oi/C52Ki1Kju0GJ
nb6ZO55TmqQ3L8uXN8OWMdijStkXkIYwMipvtSoEPZH596XOMLtYoPrYXCjdGSIn6Q+0ST534c8d
8fFaesmfSrd0rpx9JdXCkPGkwyZgFn2cgUQKvCTtLbM6DJ1nJVf1/f+XoNyoMQU19AAuIJ+U3tv2
TAs+hvXQosUuW8rrRKqd6WNofSb3HYdGHRV24EpF/nw5PJe2ZgcwohlaNABy2f9TGOefU4vZxHKE
VnDPGIHd/uf5Q0KuXSETK5GkWYTuvrHP+WXKfXuX9iQo01a67/Q/U1zAcyWzWUPQsY/zJvuDdvKK
tprjH2L6gRoLtA2H7yW2WZKwPq3cbvbsYeneKwDRbKzuwqnziKyBY8yL+UMm/9dO4Yev1McFQjMC
LfL/j+914riI7Lcj8eONPwVhTVtaNXn+Q4OkotIqP8oOvgHTtyDZmuUkKHoe/YY/6LMVw1r/lEES
t8fk8CP+MEfH8RTcfJHPBoIL+VpaOdaX4zaEYSGNAFrgwEeg/VwlaWyaE6/VfVy9T6tp+v2dsBxu
Bb4TJDOXrPsZGOmzreCBP3Va2MWFzAkv8DL06L4GMJTi4dYhJNP8t+EbX76IqvWO6pxvqZ3rmNsE
FRhpkNKlb34P2/5Yj5Br7tYcFZ3FkVCRXz7iqg7ZTdmMtJ3UxVR0erGojH7utMP5EdKvS92gmyyR
E9Xeq0efV1AbUSsLs0HYKbukbPpzei4dTG3dCQeg404XOgdbN75lqW3Qqs9hb/taE+dFJQt066DO
Z8hmcF8U+vhKSNMWUHsiA6YK0Q5PDi0vXqoDLSVctOLR5UOjbUqNjfdLB8aCKoDYSz/6aJIQ6wCq
jpivgXWM41JcHhc0p4ieOfE3OeugXfUfx6UsJdcxaB9z5XbPMzTsl66d44AMuTmaZ9mYVNIFLpCI
DyQtXr3yuFkv8yKQZwF0o5eLDNt4Flzr1zpUbwvfyHv2riGVQrNZ/+BgAJUBpKRaz01J1SMId+tn
/wmrkLj+PxLYmRbZ/zZassSLGA8QEsbT6wp+DxZvg6TBUbwfUntacfdYb7mKikOzbOZBLT3++hDp
5h/dFBHBePg+3U8y5yMkrQw0EwYVzuw7J11N9BNMS9R/73QSFwSaZIAdItZTVzS0XoHIApCkgR9z
KvZZ6zLAWhmwg1Adc26C/GkQSHwNfxdbU59tqjEq35Www8SlNTtRM2iara2hN0Laj/YpD9LFo1nb
C+GBZSZ4TiQQgxf/U4XvNDceBoSKUK3ra7tYBAJCQkftfVN9RHHmxmj42tj+gGegQ3/GUg08Fg6t
TMg7pKdZ4bH8TBE0X+h/7bwJIQDt6A6Lj3TPkqfniRRwj4/wG4oq/fmTQRI06ruau00t770vMBFN
qtXyg1yBNGy4f/s5iDHy0LBJB+s5G6+jZUvY7azU1VDvAr/W4/12yMgu8CoK7IHpKAUKgfz0cyfM
UtP9xTKxGbzd6Qu4nuqoie6U5bVPUUxioZ6egDdfpgrPw7A5ALtH+bQ1l1bDdzyzUPgq8SqdMW6Z
ouO7KQdYTjaJP0U4QC6ha6O8POnNhU0WqMq9r3nnY2+4+x2Fg8ixP5olKX0UX71joXSC6Vj3w/EP
UeNcHMfdQRmNE110rb5VK5fVSFeP78gPIhveZ0A20Odacxd3gRZFrOtP85NA2uAyMyygVYa40o8a
B48Dr8laugALeoU5ieH0KtpSBn1nsDUFuaeIteWcWm2pYINRA+/dxtSo9hp6wooPR8L0YxyWINP/
4SQ0tdfa5EALMFtY4/92GcRIOD3jYaMxDpf1ZsCdKgS8dZpc6qCoqB7XI9vZXSlcGUREsj4xMxW6
QXMz42zipIVByWXOpjXiP9dr40UcMalnND4IC3aoVkAQkZYvWXsYlLA8utyjcpllzXJEEgaGlSPM
si1toE2cP6AnjMX0RE5WRGmRy6XVAN3zIxfAUUqHaaL2sgHPjut1lD22/rtTKfoOCdsaCEKBi2NV
egGtv5+EdkvMoBlQbTtHpbf9lSebjiaMHSwfmyUcE36eECsV7sbfN4rcrt9beIhSWhv68qr2qGEc
uSZV9RiRY7kHFrasKoabwndxyQ1DFE/Yxv3exXo9ellsBJ4DYoDq7kbu/oVoRkh7OClL/1DmpaUp
qMtHDAa+ZirSBnUB6tk6jB5qvgZhJiN4pVj+eThNX4pNAtvflluW3dfr2wrD0m62b9blxBoh8G47
vfi6c/lRk2wzU+rJd4/AROb8qblL1IEYPaRmLhymcdHssoXEzbEMDP0hHoEe+GFza5ZsCErnL0k0
hu84Q9v1+lTqrU4jButkjGIZ1KZJbk9pbumSZlifB9A71kJzgxY+bTHVqorSLYN075BQ+q7m0Qlv
mK79+VxKzFMSCBik0v0Iom0Po71XgsgE3nl1nXD1yCEamOrk7lPAyh/+jN3/t4agAux7h89QToaV
YZf6yPdc/9XkTljjJ05S3Ix6wHIvLt8EXdN3lo3giR0Lm6GsHQNx4TzkMfXSdpTqJkkTm7TlWufL
3CSoJvBPO/Z/B7lzV60F5ki874ZPYBPp8qtXLoTzgbg/rbTZM5f9sHU03wFOTxCgFB2cIZCC7iEz
u5CXZ8rf1Z4PUkTrrQ5dsm1RNQbJs8PhBPHnyrHMn6E8tuRo+dofPW4sW+Q4dvdmBNRjvrY1lb5j
BpHcjv08JjKNDvOivyTDU8J3+4fFwM1hyHO0fq1jk5IhUxTGg+Ozz76CX7oUqvOTG5qSytOA72dw
xhDdh9IwIJxvZM3Eid0FY+AoU6eQVYpjnmitB/FPMHKcSunK8ZPaDto5h3FIZ1tqC8yF4Gw8op9T
1iksBAK+ZA56x7olVu3ks7seT8WEMordaG45vAltV3swbg9ielOVQkfB0mDnjeT4L7xjugvm8OcU
UWhgmKbwd4HusFXATIRX6V2qwa+z4QY3ubZbzCGYzNIiIW30lfaaB9qPH01g6qa+cgUPyhyVrfYX
dnrHxbAhOU0n/vs/MwwinpiS6jt4U4JYj2a45A8DfKJ3lckEqr7PJVpKlGjEG8TtC7Ixn0eMRtP5
nMhR7XFq6NRrJTwJa90208AoZZZJehXUBuRZN6eJS7fbWuB85RqkN69REVr/XGGyTsnn1eNkO4wl
0ms5ADpSJyBAg4I11o8efpifUEVJzQVre1KNqvpmAyhfq36B1GFqYDtK5y2aPGX1r2a25AMgf2gZ
P48maIWqqvQtWezwMHo4DyGd8rO5b46PE/XqP0saFy+oG359U6PvE0zPSv27oqfrBvurNXODVwQH
GCQx2sccFrUeXgcD02f8JIJApRSfDpaktc57KE4HOdAYW2vhhEb8swK/d71KRSRWHSt9GrdEawgm
KhuZOLlNvEylq28IUI/D6xvdH9qWg+KPVyrJ4NoEbPQWY5+JEhEBvJVEDFHSmE5st4BdAEgFLzfm
tRSaHeHl0SfNmJv/6VcfLG94EONV2WrPvySFKkGE4lZhuWa06D6QbDDx55tmgqHCYh13bQ7kTs2c
rGIaByCHQ/hzp6RonVs5HkxAdn6EUZNxj8gDVbMr09Kat8xXNpdjqSYGgSWxyp0WmUyEBnwXP+ve
C/b1X3YQneZEbX1q8AE7ysracdaE7rs1vX9SnL6+NQcUQ+ia2iMPfQZnKvx9LqyQBzDVw2/R5hUT
ugROJ6XmFqJKq4Yp4jaDVx2NaG9MKob+4Llwip6ez2zfwgu8RRpvXnHh1Ky7o4KA/yYTVfMUkFR+
vtsXkAW8HBbTEJHHZ+xs7fY8EOx2Yw/Pes23UxCstPWKZj3NWO6tK7TYE5x5F+1Vuj3qL3uAwkES
9q6aoWxPqUQeMo3NHnQbaYjmeCblKYqLtKoFyc/BXxB6XYqVBNdCN0hsQ5LJYVkjw4zjEF4f18RT
JZSQ0gHi3qqqQvoI+FEgzzBUDVoHdBIBabRZJZTbmjixCmnh9scE7H7zKhpxTPCpt22ZfXwBipMq
0AFD1YrRNucFN1Mtt9qSY+Zm7fuFMsV+47ChpZcdsUugwPird8LPC/IVKzMev4T+BpcWMiI1RZVF
a/+ZLjMMvR0QkJmvZzMSvejL0c6JOIa6ldZuIpSdhn/o6ChuRrEQrM80Qo/pz0tKcrxMH8q7iIU0
0U0RyKfrNaa3gG24mT3PT1W8HTl6A9xYTuPpjNYVBN8nzebsLkrqGpWKz4jE1/AnaDiF15EHLReW
edYWLOY0ANy8gImCNh2yj+ZgQSkq48EUt8p9HV/AAn429vy9KezgNliUAou3HXXSAY7k+gr4cAkq
quMb1P7SqN8QLBClYeHWGOjJZyz/QKe0g3HvAiEFWV8tkp/pnWawOqPEsgaIHbMK6SlUjY5236IB
j8aMsAJ7hLGr+15XwY/zubj65uPHtenNRRDk8tmUzdcwqPxSTFH/9WoQlMjpSBvIvbzARlhadqLQ
sInr4jdxVd6eBzsnLsQz7zNTSogBOOi7Vv32nUP51Rvxhd4y780WHtulsGj/xcVDvZ/+dh2Mn0oM
gFcH6mPvoo/EMUevqKhTQT/CesM3l+LbFPR4mn1HxBrCeWh7jmFwWErzrC6EgdNtwIQ/yX+jRTCa
zF6J92dmSJM+afHeuwW+62MHBohYT5+x3Acw0B7GLyisW7Yxn0MKvtTd1/c7Q5JBCuY2rUpNivFi
BFty2MgbTQWyaXOphlCykvRkmVXQfh22hGbqU8kV2oZzWi4WIxe67bjuvPiBXIzSVCl7Ifm92kWL
TzKcWTadEsU9XGVmznhjbXbwWPoYlMZdE/QZMyyCutZz0C5SlhiurNUxKmEBhFvPpqCPflMhSvgG
ZAobSlgv3exolhlbhBSvlfnX5x1V1ZQoK7oPTV72005/A3QyhKoAStHQ5VSPCD4VJSOVcgFb9hVn
KKaVXd/Pj0QEJywxdlLOB2zkcVt/uyBy2T3OjQ2un0RkJ8RfsYgIWk5M6n/EdWVcqbwsiUtkjgxw
sZ8vBcBDZvT/TFibK2PM3uF7x5VzfzaPtOYzwmKNnMHmqE3OtkhRg64mnMjy+VLwNn+S1nj7z4Kz
lkNpQX5WnciJBDhIvOTCHKISdOvnqLZsbKfXTkql1kxxioJ2G0JDN5XA9C9NttANavNo5GdFyc0k
UBGM29KvrkeordVAG1+qvSg2Fu/FKqxl5tpKaOoiuuzmAH7eRENjj4t446LF+4FznG3SXLw9IH4z
9udp1ykQSt2gUGtZEsvToArZi2mRPgyrO+INZmPos9q9r4VAkvKH60DPZX+y8WxWk6P7ebYvBMHY
Ed89Vigtkl312pBXtQzgwAxv44om0w7o5cfsn41pKuTcklHtQ0F1LPdLI3am9m3pwtGJFuLzBgDY
CfZIt8e3qRBhGVveyRcY833TY89IjVMKbAlr1jYfF4gvlt0hfScESDzWOTxoKmwt+F08slQRlDll
ba0LUerYXTTfBx2BaXINOzSk7iPoZEaUinZAKkXEgNbLJTn1/V0qnKYRv18OeDSlsXwWXC7Lyqha
VT+m8HQqj7BKB/RdCg6UcNtGAMgNljEpjdKmzRdk7ot8Q1r+PO9Dzzk/5qAEAWHZMfdZqkTZG1Un
V1yVbE/AjJEdikM9pBozampIUJ4MMcQuuRyIdzgUu2TRuniLjoOt5WFQOmb9iRbca0kgTmwMJR3j
L8hv5PPn0VoIMso6NmOZ+qW51v4uBmyPBCH44Z70psWhp4xawWi0DgO2hGXZ0csoSdRGF5cBZ5SQ
qsOdjKhrJrNpf+wO/n1HzF4h18vf8G83WLuhMa5bT2OSvaxV4kS1haxcEwNuozPTgcAOsT0Ks5u8
mlirugKlDvsDB6vaVML6Kdsfkfu1zcNCBug5ufUYkML86vXUkjC8nWDj3D6rzFkiOdDC4M5qMwRP
AHQ3zZHU7nSsxVzV/ICuNngdjVhQROkN+vbQ4vpxM4IOYtCz54c6VNTZvu8uO6kJUYngpKp0UGA3
YaaSeWquK3o2TnFcJUO5mwsr4uiD4w0/yQG/xuXrFqcPrmJ2YUT2am1sYsTEUwYAn2SBYE5siAPp
9ZnfLSbDZJ8GoyzX29oUijQIZHoQhTB9KTWRD2UYOYomgJr+PvpMsc4jhvTYq00aIcJX6f7p932p
/CR2hlwu2pu+fHRGj0tjNrOK2M59LWB3iFbgbSd6U0UAZlR7YJiDXAs0Q+T/d91oO135vmXJ0zor
kNSt+tX5K/oQSivMt78mT0ZRUiA3OSyLHcX3F4cUKOH4pBuLajBCHVUwmByOV1nPN9AIm2w3eo2c
RDho7DbjhwdWdXr/7jp5xdDnXCXs7GSlTM4/gAphHbMOx5hs2gAIyq+ys3iKcg5gLbDHjMql6xof
90Cmx+X1Wdy1ojXrQ64UZqivM1Qu0aMZRKqPI6HmNC+2qLnpkr5J2dLcc/EsfxsCYN73DOV5xra4
bDz2Kv6oN+PmQ0Uh4L+QXFD1rSbENKWcC3s1u/FUOkVyW6t5HoXnj3PtdkGissFPEXP2ETxZrc3o
RJqpMYWEVPSrieg19YfjawBGwNUm+5amppBpbGs3oaVO2atpazK7bLEwdYKhmZxScrfOq+5UkFX7
dmdHl/LqA06yuXiZXeYR5TSRAH51Q3CXHurDise5Ep9zFvQ7W02HMmcweNHsqoOB4WjeqS0hy55o
cVKTEX2eDsgC5y32KYQT2SvDU9kdWm/bIFJE9VU4OFc3xwTHoTMtmznZoV0Rs8gjXdBBRbVsMYNb
0auh+x1mlXWDxSJhFO26WECXMO0K73cG62OBooHMs8dhiczW7FzGxcjtuCJYbrFYwtxg/7AUpwP3
aw0xt79MEBA1HWVQUdXXkuVmfS6XFdX2IZI/E6I0V+j/rlr6/S21HHzSC6k0MdlXj/upd4qfHIRv
p8ML42z8xh7xYmylyXmS5ljqIIds0WAHqNN+rEE55KN64RjTHIOOROUUgZtMTIk4hU0mZ+LH+VIa
vIg+bDDUt9yWWk0p8pzVZynlzLD/OugnrFaYrYVZleuuZ6tg59NIcxQC73Pw4L/jamtMMcSYFVdY
qNgsp9JE+Y0DnTtxvk4H81owMt7Y2YQBI2uS/p3mI/I28/NmIxfmDqv4Pz9Qu6USAVkqXNU9rNXB
UcHt0LVKKW1MDETYnmXeXyxoslphxY/SzcPNqW914OAoM4x+HfVA6tj3xTLHeMmehXnImfB7UwxF
jt3OhqhfbIJapgHfZEnL63Gj9PYwZXo1Pw6PN5xTDaLkj8cbl29+9K3maIj4MvZ/baPN8IXuCnU5
SuTq/ufy65lJckzEoi35384jvEVkVO45l3jrwE+PyfhK5gTvpOkjLXXP8mxjfeM8TUp2jkI/Dj87
AHMVlBRA1N0iK2S5XAJjPCOkPa+Xq6YYq0Jlu60gl+XjpXBP++U8v1sMKeCHmp3YrZqrs5WZ61vj
8ToyVV3ZCgcIKsotHdiLG34zpKt+Rk2gA3GlQixcKFTMGpiWH8CxFni7kxj0ezroqbm0ws3ELtA9
tSMoL9AtSeX+ogAP70skGfAnJklly7HMjgy3lIZjcIpzPSC0eRcfNTs7Goq+StJRDLADfFldasXf
GbOt9V4rWIUjXLMUk0rrOQIrUN/qSfs9pjmMgnPwXOjafsmfEqpw/NVSRSV4dd7wPRTY9uB28IhH
vGw664K9gYtaRzUaQZrH8d4OGf+J8xsihF5zGzgiQeoNiM5aCmGU9w8il5L92auhF9XTgxtmwlhG
SBp1foGRISGu6FJOyuzFHQz+X2TXnFtusfdfuMHwgypfAjcWOXUd6cU0s/bYLBNyMwRjSquWH24Y
w6QPCD0JynZDzpQQ1haIZh8y/iRDoAN7ntoSTDMXZU7tLgM2AAgZKFIVDhngwN7ad62/wJ6TD0TC
fe4Xqnb1oyNqwITGTeKW2/r63fSMUEgrMqAz1wFb5YoRjGmogwGfo/ToEixsXK9IUBVTQ7rbjSee
lQleoctlfkQeZBkiYeV1+Gl023Y7OQssHgYBSSWE46/S7HOB+dgRAGzqwFQ74uXzhIdOjvPw5f77
kwcLRjjKHFyCH2QzPzyFwdJx89CKyUQy9MZTHZZ/gT8ba+JSA8BMYi1taacetkoZdUbEJiTZMhpP
CJwrpx+ZsOTorVYDcBK3iwX2KGKxTBNZRR3zsQj0+ZbmoZGyfFCIQPnRzD7o6gyBBy1RchogEr0x
tnADWo9u86v8PIFk2n2utIH6t7Rzv1KOyasleoxkzZHwLxpVJMSqAo0hTt6g1Z3+CA0l0UoNUqbB
2g+s6VfyxDKRk6AI2Fh8kCSPvsqIdeeZr5GSimJmqHCaPrw+NAROu4aS3IZfvzCFCC42/6awh96/
zkSPO4H9FR6mFwnuVdOboHSN56sUjLQyLl3+OxQ/uUjQhoYPNt09CzVOO3+nuCNdufkfFk8cFv1I
W26+Uo3NwVHo1a8uYEBjJA73i0Zsvg1Y0wc6UnXeD4jwvrbvRGgzH/QTgRMlg5xaoJjBwsExjnZE
7M2uDFaMCM2TqpWBQmqIFy56ZQBrH7jvcLWHqfdQu7CfYvH/lZCHLFEOI9WC8byeuBUrQqcHPw+f
XgmQpIm/lsTf57gCOiwKkErYHRfwsIiaySQQZcAt09/whtw1D20ygEHobqcrFeocHjCErXSFbN/5
JIWtv+3oKvSdgXA+1p9Kfmaw3g+ZZK4l35dRXEXLufr7SQYxMhTqRX3asINyQH64OCg+ezbJV1oV
ZrDQy2Pj+w0KUWatwfo19veeyqTHVtA1PNkMrKuCV2R5o4aSXT/Nwww2hoAOLITgC4NwbBmTq3N3
0yJh2TzvliKSCA+qTUTjNQG7695jcVF8l4X6vKYuViRZwhZhU8Tn03NqvdQ6aM+Y3v0s7u7qBRTC
/8YuVhbLq0B+O0T4IHyndtAB+nY6z8Uf46t5HnGXbXFX9SIo0uFFmBerMNEZKikh9Ajcmn4BG9eP
0dUK+hr0wKo8OyW0/4hjG7xnRL3jndArCb/qssYgNZ/514ZcPlUAD7rkLsTn9AZZ0WR3kBMdXeoG
K2lYadBT3pUUAgplbpOswGJ9aupujGL01RTK+nFzY/yNP35M5VEPb60YWMg+AkCXYFeEIqzC55Su
wMc045l4TGu8Lc2LNlU7bkGEUlXzeyY450AORU6ADKUAKAuf+EafbaxVTd9o8bLaQ0dwEzKIBiKu
g7LMqVhQPxgMkABy3n/p+lTUv8STn+gnRJWr0QQ47A6oYXhMothCG20wm+ETXDxiQV0LOZtr8XwA
b00kyZIWgKzqceOHtsNKjTc7ddmc0sVoD91Yb4smj/wZPjewhgMMu11Xt2tAC4vlZ5XXRTD+Wzds
Qznz3Ur6H3z25rit91Pcsh9lvgFdzemDy1I/tIYNAFrSFp1tHb/EE7CGbpz7Vy76FjS25XbXIgC6
DqtfgwG8AyTjgKfTexVBlgd+hmWShppD5UvjWGw6F/tgCjAEjU1XNGOL1QnQOT8FgCFycUFP1DCL
Q2WznYzTsKIAC28DVxxhhDYh8NB/eznwMDUOen7G2i0n5WVplH06XqGr9w0Ksr8+COzvBaxSv9cI
RDvEUGEvGweDW2YbPeQ2oU+9uSdZxXXmvP290haMXOzsbjT2LyKBwirGiAGvJrbqAzIIpA8XZDEs
9a+Z4b+ahWu9AniFShODA/wZ05iJktfyiM4GRkp8guI54qthpovvJHSPwnsUxCYnI/1p+YyS3Qk6
X922kRIcevrQYP/sdwQRdDI4xMdhCIH0Z+PRmAcE7/gaR3LdJYC1rrN1u38/kpREzpp8viJDYL2f
kqtMSCGNVijDj5qirYi9e0TMa8eGRk6pgm2BrkK1AUGQoKg2D77/2kNWpRkyIRbNB9M6MXrJ9kdJ
ediOE6KI2uqSbgGwgZ5e95ip97uSnl9lAmnmtqJs1zxUy9/3oKPR5yG4hlStcs/GH1IPIdQjF8W8
vg6v5KzImF/baBqfV3G3i24ARmz0BKb/IlTKl4vDrK91hhd0ieVbX+iXMN07LeqMV7klgDmTCxS1
Ws+8g9o3obZ7dQn3I7Ql+vhnVcJqHpr8oXD+VQKddrjXFK1u1nXP3aXk4T3f0tY8WTaoawnHqRxp
uPsK0hT3YqPDGFaotI5MkS9aqXN5jZYQJDG2tIS3b+EUqFibkVgV8JaqleM0mac8aF25EtghCv3N
iYnpNV+APwf2OQ/4hR6cy5RKGMDB4kTG0LidtUwkNW5WpUp4/XzYT+kbfHf5fFHsUwzA/KqtCMgr
pFIh5szNtkMmzqgrhdJux5ZTdGpeN05SB5pA+CVNyAuLqlfmyguNAS2ejC0w+AUj0fYD8M7eC4Vm
Zy0ctttLsq3lpcUTQjBSNXACNL8oHyvB2Rmh+rnQGdv0BzxbzyZKmVhNLnc3ILmzzbn0owAHJLC9
0IxwMCJ4BLhfgEhyB/BRYjWufq6HxCklx8AV3syZ4bIuQJTBAenTSz8hUHYgDHi9y6nsO3cFWn0K
Mj1Q68gO09rfZ4rt/N5MSZCWLA5XRP+W7N8PyFKbOKBEfjJLxjLnjo4BtTpDBkoYUBVmDa9J4Avz
Q/ZL/MABp6DmtcMN8RZbDnl/DMSn9kWtphLavtSLlm3fz6P/yWjzolDfSSvsiLDqa+7SJFjmcqBH
ifNpylvb7jKIWG4CMOQKq0joBjGr3RWTSiDPFbamJ8kF9dCn6n2XaWv5sFzkWE83FQlkt1Y6x4Tb
3E4gWNfg1881L21Fql5hGmCNpsW8UXO7XRof+7NiBI2Ifuw2qqNgQZXWOWHhoaorm6ovLlhNrVs9
k7mTQh/HfAeVfL7wBlBOAu5fUQvcM22QA9o0wlrMh7nEhEsLiXHNNQGn3EbgnzXQJxrcqDoXo/Gy
/lfp3y6JeJF7/os75o5V5+3RxCihej3afg8OJxKNkZCeDHUpobWSMvYN5syBnpKorM0aYwTtxMo4
3aYJoau4e3zH8OFjb2wQmC6G3FlPTleH5EVXDaHzoXjciXFcZr2IWSehJS0qg6PhbCEWRY2Zwo0T
ynF7TQZtoTMv7uJ21UEgs1NcIerobnAzEwGUOB4THKf6dVerSJaEmW6V0YIPgF/5AK3NIgXBkYuP
OFJmxG2ZLLZUMolmkwWIQUtFO8NM1EUWO4x2vtkA4sNv1J1+X0tGxgwbdsUoyPuJmqqNBpFH/w9B
XnGLBnRFI7FKkpcvY4rZyG400+JP5YP0wVjbgoUAKCiLMsRaxXrxJ1gFza+tReQBiMDpSi9JcRCw
DzDnyFRnVAZNDolcvrW9gWZg3QKIE5qJvsGF2CrNZA3VTSq/xDOOA3jfOhxq1i4JKcZGnUcZsuM5
QYZVQuNhC/erEUT+DV6+TuSKVc5n8mMnREzrfbq/+zKPTEJhD7A7nQX5lupX7iE9GiXzBzZ2Jt3r
Eel6/QsPWoNX223kErKy6u9Kjkn88pU7zr9grhRVqvsGlTENctVoWKikXv6qySX5hBuKpRO7LrFk
d5miOI6lJkmXcpzfM4T4veqU4E02FNFd4rlzJr4vDkb1bSrNpH3Gur7dUHziHXsoidoKdhza/ISV
aorDGyOzCMWsOkxwj7RK3XIvM+DFn/Joi71NgwTFv1mNL9KoWBNVpcRdreDMOR0LKSPEQ2dcl6EJ
NMFwiQo8vvbHVHKsw9hP2X46YT/S2rA9rrBJ8v/mLZ1FpUshKfiMPgKEgm8lSUbP8jJy54cPC960
lQO+Dl5u1eUgfvfH+oSXUbNGbo4mY23ZvgMXpNIdtSINWZ5lzgvIiTL6w+BLCc/rsTurQSBOFVA7
UqdsTFqlbaX3JipovsOiKxWWKwLe3BlSf4d4Py3rwOlYFcbjcL9aCkmOiIurOZ5Jfe4IOH1klpb+
F0XDx4/Y298Cu7NtcEDX7X2RS/v5vpyGTcOCyMcNOKX1foJi4C7vFZwGnRr9PaxOrO/7AnXHB2o3
AJcKWHYjXP0PDUoUiA6TygPnT3E6SYGTM48n6unJOg5/OMrwQ+plvwk4xbcopsoaIJL4U3fC+Or1
9qdbmGX7JHEfxSXlW9CADa+YEkNV7hgDHdISVVInfrPQjHUP0PObK487WdLNqPKWJeGUh1R4JeZo
uqU+TYfrdf4aP2Jait7Gsq5RW09TrAIlxwUnvnWiyAogBlk0/gK19l1JGJbSW3J1zFbZTmS2jaeu
T5iC/emKDc825NrBpBmhCsaScln8vLrdJA+tMBP15sTc01rQNlSIOayGGWmrXvtI7q33JLZsveON
eEky8oXMv7ihf1uXs/Eq8n+ltPL0HUExCxG1Wl6lwJJioocdsA1hR1iM6obLnGQluEZspVrUIeXL
Cr1v8jxmQzndfdJgFa2bu9+BEQftatYN0rU55IPdMYkA5Qv96gUdOc/NY+yYEhSxYLsseIJw5hdQ
LFYeMwBtCSorC4V8FqEpNw6fg0t0zJGnzj6fwEJ0JekVV+OREwyZqelwVls1nVI8bPqI3FZlF/tQ
BFqCasn/Ag9j2NBvFXeC3YrsucctpHQNlu2vk+23Up0W53JEKLry9B0mHB2TJ7RTj/534yFZh77s
hfb4AVjlkFs70QmxMXZjj2goQWu+lc/NDdflxV0Om/KlCO/EKjeyLO0wyxE+1knT0/Oqu/ZHhm0p
TSCPRL+5yaowtu/0yDmkXHNd0ny3LkqRjBHJmOtYXwoXRUJKrvhJ6CiNkXbc9W6BEoOVI3LnwoIP
vasmWlBqlRZYx7qZmWGqdUbBpkRtM1QiDvJa3POJG4Z+90RfPqLprazIUS2bv3INhdRub8U8bU9D
4v+401TnmOEf8eqLEpcTi7kLMnX2BV0gIE8mo1GuRUBRNyIU0fkCMDr/J0q6NFBE5QEeyPgvDxni
DEC02rRGMmHIdHXKeVp8EjMVnny6Ju5jJrh8eLiPFq4sU2MsNO+fGQolgqVPkXSYjoZq+Qrnl1SX
Jzz61Cuxy9ZIU8rw6V9IceijpQhFvU4ymdf3KeXcRB8Dy8jme+v+q6E9CyBXxEW4ntHuv8FGeWC6
ALRL67AC1MHGps3Bkneku/vuzdbtr+/0kQ62ly2eDf/+bpnVRGWXNB1gNqvHLNaw7HoI/WpG2At7
ujSZxRlTR8o0NUdI5Grrgs9pAdA1Q2NLWXS+6Ll3bFayTARfkwZmrxjt9CY60RFjTqH9Ij0hs0OD
PwcH/C5joC+nHL9R+ZVxqFfSOjapSYtUo7oy2cqmakpxdIdsPb16O6qXY/fxPmlMOBL1XzRCsWKj
oHgun5Ac/2gX7+v623y7Qsl+7v983YEuHj2UiLojcYgQ+tNOTzY5Xsfk/V6gPoWkyORjMkjzEySU
0gno+XLLFPXh29q7iYKJWP6iQCaykvjuLTVepGvvD0wrNlsmOtU0oU/jJUC4/ZkpgIb/0wsRghh2
TrP0CMc3GGmDCKda28zF+YXvFDsH6PzpLlOFSDEetlPz1HPMwbGfngNjU5ye++fwyZeiUCGf03QX
ZrJBj5z24TF1p428lXt2aMJcujHmxOx9d++izMO0+qHcwPxNB1AR+tRAOEvXHBKQlAcB4jLr0GNr
PfK0CEvAXhx1IBIzznIMgtfCNyiRUzdzzqWxKRx2IH3CD9GE+HOOUnpIKYb1a37h5dfqsqztlSgB
fcvBAdu32jP5dD9WcAMpeXDyThIYC3qMiJQzrW1gE3vE/1Z/vJ2iFf0H5qEq/LgFDWraGLYEvxGk
uXIvaTTPM0nSEUfgbL7Z0UI5+SGox2J5JhD4nVi5dFAFGaEY1nI50pb3ERWXDqT/VU6bxzskXZ3+
mgoKHysMgUjJiuFzeWt7HyoGNgnN9C72q1n2Ve0+fMRUkp77c0AbzQJ6GmZPe6qNr1aAD3lOJs6w
GSNf0rXXIt6DS3HbAQCC8qbRtP7QzoT6nHwFB61uQM08v9vJaj5dBDuCr7rqI5NKEJPNZx4n6FvH
dLDnT8JpgF4zE9dfWXA0Yxva9GxQcuxM/W6v/CztWRRBF1aHd+icX1EeSK2j0HATZA65D4boJKQ6
H3faIFMhGnP650Bbqpn2+iRiFm2PpDe9tyaihQm+PriS9D0Fn1P95AOy7yhgCIoIE3ouVG5WbJTu
96w125vJ464YzYRNanghSLVWaUfS7tYhgc+CHyYFf3f3m+HqXjlCTo30Yd5+Mm4hIfTQBC1eOPfR
tg86qcjwJnUDLIWYXbMhRur4nod8SP3s5uIEv4hgSxD99AGKv/wLmHZ7d1mosrKXCzwo1RZWlhAq
wYCXhFl6UYMuQLRnQILTUoie48kEAJS5ZukjFOIL/XvC4IP/R2QEXRamxBZSBhO2IaSvx7wUjQLN
EIjSAEpagBIQTe7KpfIFeuaN4Yc9puk1HB8TmM89b1JBOZDZhBvzbl0jTVvE+FbZ8jU22mz1R9m3
5sjRrWyrKcErUxTbCayIeyJJf5YPQUJ1nSb29I2TISUISjbJZQZq6J5rjIBPGoIeXaD4lbY8ayjU
d5We/07sHY23zXKcEDi56D7tz9xZS+AeJu1pK18RFDx38Bti8PApy7p1TP7i6J/KQaZ5amDlzWao
fSPpWRbASQRQ6Es9rrj0rK796S4vhqBmgSc3NTXxL2WPYaq/RDs9Uwxf9gAb9vgOg0BgrOcQxtZD
La6kZaXY9xHfU/hNDYmX4Bix1iuaei6/ou42j16lWikhlXb9Zl+p1ASMCIgbremP7AMgcDqwPvXn
+G279cLnubfjp61E7AEPjMl5KTVy74KiFd6ISUwRXD+e089ayt/7KS0FxtxqAc3MYuPJtL1zJdQD
+P4A1q1YQCkqDzTFovgcNiAHlFuYqgUVdtKc6DTO2cAYPOplmdOYD0IjPu4eNjqhT5F6ORn6xkPa
DgXmiYi1++31C3NLGq4yLhSOzmt96JRNPNqdU2WrNgNw64NXU7gqNuBV0Hs2Fyxph4YA+1bapvU3
E5NfRRlsXRc+MNUCFZSNUa1yAtPS4HiYqGTdJHC6V0eFoFcuCnICiriEnI/ZvCOhxYOUKjCmF553
jwn9STzm2aaNXw1FBwghKeAEHzCSpr7XYIpJXYgV+kmgEtAvYdyG9Tc9VM27ZpHrgMishYj22nKY
Hyui4kjm/BerNYFsPeq9tb880zpXQZUHM/Nx/JEsWzcHaCj+wJO8OOBYTNRICpSpxEZWdxe55DAp
/axokBuoRsBoU+solUSDdr6DpFnH/bwYZ5mf/RAmJq0eYEMcwkH436aEFmnGS81pLAJG/7KbAB3g
Z3McHmqTG7ffDQxsjxVSW008WHFZJfhJFFHwnw37auhvLMakCJAKifHqnWNwryIJEiniXxnMjlax
OCpW5l8wa7Q9JBxw9qWIjUNtdmWRrWwcNPptj+yQ1gzIeNNEM1o2oLmL4Y1V8xUE43LpNpXjBi7+
vBm+ga3PJGxh1iu0R9nwzRJUX+n2DucIXQDgq8Fo1VblwF0Q2yuQJPksB1ghudcQqzzAJA1jrQxK
DuJeWeSEQli1IQJ5Farc+84tkZYDJja8Ep+w5fFr8XjxrnaIu19597asujJZVVQZh/MGjrzkg9cn
lsWyFK7nPytMnwGMUuh5Nwcs8vZnXobUAfPX1PAF2Y93W2e40kq8d2mkmCCmAe5y1Y5yrrt/LyRg
JdR1NVukG9HG0EjRnIBTsRq2K4qVVmUjQ7n65CTWspxpQ4gTwJsRcxV7nyHHb9E0LEgOROUv7FHp
YwsRvm/jx2u1wpLVDie1E3IE0Bv34Cs+Q8fIPDw+KrdS2+1IEbasigQiOJF1arL0iny50EDHKb8I
MD4OEWTelPkeJh2zojFPXb7rSWC7f6RqdjvMqP+FZTILuSkZtGfys17nLjNr0sPS1whlMUF6E5ZV
6aGWjBKNGCvsIHkNlBTeSDRbWQYGJDD2m4a3E/8bYboRq8wrZYLtwYfgwTNDr4K5MoRKWVnt8Y+h
tm61OC/I1F0SUu4YfPf1Cdl3lQdPwjNWOKsYIcVcn0Sv5G0KdM3rVpUltddbvloqPeuMpULU3rQj
ISJPDnSEoWQzz72VSm78wadidC+0/p8JEW7fivu7+zRKRpDuHeFYnVgIW8Z8roWwnULPT5SthDFg
XCHP5OXD5ko+z2wUBGS4kx8pEXJUSp3Y0tPit6Tb/UheaPkqjgXM4WLdK1cj2Bqoo7gb8+kUxj0d
3XTnwSXJrfFjd1oa7XvLpuS+n1vKDkd+SaPleXiNYnZpssAuEntujRhQvfPbNavHxouqLP+2F5Ii
dOSFYqkJM9fhElWqT35uhZMe/BHVnE2hoV29/6YzEcC5SiKsmWWv7/uKTAjXtgGYgrIf5bKKeCQL
NQ6tldfk/aht8hiKHyZUZ6kJUIxxbncHFcYVa4pTY4dPsF29bBUKqD6DDgzyop8Pjfp7Kx6qyb12
6C/X8YxWk5cg4Yc61FwjWwh3Cu8z9ipkBfIjlxlFhZaPNznqIyujsC/Kba/jwTNiP3Zt7FQkDGGA
C9ckN+GTYb75o37Lhuo/vOmF0Aq4ipdpPD3cDbSmI8PnSQ/D1E6MnRKkrLtkhO8yD3G7hiVYcMtc
rci7nbpj6AOpGBWeqzkTvgTlAJYktFMovCZRKrPeLOxVggIwDzxFcORAWnyg3NLv+uIETVwsBU1y
TTXlTJmW0NPXjfP0AgXE5gTNd9Suk1I0p/eYElb9teMMKbbMmbI9bOH+QIxZJmjSzR8xbl8lv9AT
QiQ+Ou4x3eA/hOLMkp8FUwKvwgZXMMm/1wbelIzx7xSAl6cxUOQLzW5t7J8aMWSPxvP7MxWF7ty7
2hjvUSgSv1ozbJe2sFlBEQq9MTGJG/Pwed2YSS+6wOFFiNox1o28pWR7p5Js4pptEqfeSErH42Ck
gOl08WxXDZ13fuEorNVCJ+uyecNTH7WaSOhGpeOhnFQtulDKrRLD/YzKhC0iD9zphb6W6f9x4J1X
IekmsGQVGigwnMbKCEfh5qnGGo3HBfSRiHd5M51QI0ruOsVZii9N+Ff1ETXarVet59mDeC6nGDCh
/xyT0HBEsDZAHhgV2S8uivWHnfGMRSOMosqVTbsEgFdWArbDq7LG7FQQqW9vBy0hFTpaf07JLyeP
Y8ZXlYSdegK18tvqMugUZ4eZ/WjBnfVeRJJnnO5OMtWUg0Jxry8WWSPhzTg8ErJqKw6/6C4sybpM
5e4/3xFDYEPWYhwJk4+rjBYOl+QuZX8p1xy0p9I+aCibrwLeFwOqgVhRZXr65kDBD1JPQP15oxrq
xF/0It/NWGU+WU3TrJyXKOLBHFj2IorKIG+x4Y9L2QRkAFv76OyzCnmF1XkdRPS7xySCQnk36lfw
srGXXSiAaelYZO4LskGY75TxT9AWWbfti3Rpq4A+BcSH1RAwM9/MfWeJuMHBG0B79lecDikvcjOi
4Kbm/fnErC8+eWF2O1zIjr2QG550aU++apqC4lQRijlsc9SWpOwLA2JSzB21I9uD1le6jVsG5BTL
/EJpx3lVR0/6f4WhyrdB0lNa2NiS29siWrngDQZTTud70I2HnERFhhDs8UHPBx/i6RrtpFs1juNQ
8ugaeIozJtFqroLSprrNC97PcKByb5tV63Cn50Sxg5K8Cx7VTQ/LRgSuMmbLhEOI1tw48fd5lwNs
K8LPLZ+8VfQvng0aon4oz89DYoO2FsHR88BijuXvihMmB1VaFg9Ys3qzFNi4zCPL0eDODrfPn9HT
7iljW62LYgJsmNp61YljkvdNQIZx1LNwB4OmLfu6ETGQSxXAJVWVdh9gc9gY5OyFC609lt2cTeHn
IY8KW4m4yaS9XWz6osDojlcfcyouAViZLj/EfmWQS0RYauAOoLFS61e9yRXvvf2V1vfmbMsPOk6k
15kUJTU5q2zfWzSudzvOjiK5LBbD4Mhp9t2YzbVroVf2BbEh0iatSK1WnxxzBu+1g5Pb9/I5QYcZ
opvSbeA2RNeeEn1NzlHjf+HwlfjrnVCXhTnCAExJZmOHbK5FKP4J6JuE+Fbp3sFGDkLAws1kZY4n
Qq7WVO+wWo2h8wJWTimdv4hI5hQtCDvUAGS/bg74B13uE1INK+ujudvs/Un2mYXkRdUH8Ly7N6c4
KnJfjw5sAC5TswEMMV0U5YcW7kxNmlJaYSq6xM2VcBoeypMqY3w85L1u3PlHVrfTxAC+IIXlMxSR
UVPDGD/+uDUdMtIH63DitG4ZsxjJ4DLbQw04T0rLDXjeu1D2X3Cq/gAB+OMvilQi0OKa9nYQtCy4
0R6ITVZZIxzzXH8hK1mdsiWEZEs7Ke+ZySKQ89dwtah3dH0rCQOc1yh0JydOI5V2/+rNOI61KTuy
xwdvANwjAW5BuRo9XrLBNjmrdJS/XR6804C4oauuJ6xuHoI8qr8SR2o1H1SbuvrJKJCjaqYA/lvG
SZfU8Ia4D+W2aB7y3t9kQIWjVSXU2JIswt2t41wuha/rVmdx9LWUHDrWhPGWsZro8SlHYWKTmM8K
rvIXPuvAQGRkbeHtYPNV0ozBf2/N7m/jmH55zpYqvxI1pkMNHHQ2PbI1YIXtRwhDUbYaBUQjjWgs
gRzHTomigHqotgN/HiIEm1bOr/uhLSAiOWYkzhmuRvgGJK3WL8jdxKbZi3IjbL3cTUOOt0qEyni7
7KBNlRg7wsVul+x4AMnh7sKykZHFDPJyU66K+yRTT6bbvRLNRS9Ot+mYvGTUyRIozUSgDo5+Hctx
dCzSMhvPD5c9DIBcYiYrELjdVelAj5Wr4r7dgvOv0ibgyOePKkUWQH6q/cUdttDzEgYXc40Vy3wy
QOdxaAQMOXQ0Au3vZcdAs5ka7YKVEJytkDotYFxNf1bHVoQLpn5kE2zoMk/7hAeAnIkgEXD2OGWr
zA9sFtgOUvbKdQpjV65owDd/TTvp64COH5l1DnN0HBq9swXNAfTYtkZMntO94OZX+kzew7SEGdQB
0wQxo7xuOU4vAvd4s1nV5ZEHNyyHwSQxUOJhfAIKemhU7ZJNbPdXq13GMvbRFC75mIKMUgk/4mSe
YYj3dqccYE4giWB+dB1ms6sMh8MI0lp2CqSixgAeLxC8RCf6sXSPKM6DnMWUPW9w3oN5q2IbC6z5
YiVMzXQ1qzD50X0HDlDz1gh+ErgQa2a8As8xLboewqklnOL+JXJdsK7OvKFqyoONt0/cwF7C3EK3
p9f0LvLTD8jCMz60Xd82Ykskc0T0H1F9VgrGtGCnkHvAcy4A9mL0Ccr+8Fcf9H6IxNKaspMipffP
/hK8L7B/iVqX2fdX0N0KBNfryfqUVOmvlxkGtWu8JJegvPM2018Jmdj3uHqw93LKP6zJtk48AD+o
SKlayyXjbdKFVglp/zOl++Assoovak5y2nZFzlRTVOq5/2Pm/nNwHePbxQFqO2LDFXklmPEZaqBg
tmKjD3PqOYjUCiFEEZ7T5aBh2Q6cYcjpNIXG5JrsbQg+wIVA9+FplGS4uQiuHb2q8GBby20uqVBC
R5nIFxzVfstiL62bdYhxjgqA/O53+V8+yVJLMtA87sOv6b+MJbArnaQAiw8mNnaSGsO7+Qz2ONYe
0+zqP8ctFp57THqqAONF7n5XM8ZogKipbTSJzSX6i0w7ty8Bl3yYWWEIsTLvbEt015GdV2TE4uIZ
Lay2XOyugUGW6WInPAdicVMu6FoxdQ7Y2prJzPa4FWs2Sfv4weHkD6sI6i0mI8+pv11xemaYXbKW
ch/SaFJPHIUAnsaUCIkyAYj3Is6aZi+ookudHwhjWFkrKt8hrNVpDK3DGZYSP0BrYFHgR30b0phq
iIEN+rb8gpn0DW/jDB3X3dPf6xTdjnYkcrJ8mUIfDD9MgYFmu1NRVqS2q8WC6KCmCl13Of18V9JE
e6toblXUIbpJcCzgReDXSldqQFxXq6g6xY4Miifvkyp2JJROl7dYzfxUvpB6aMuIqE/f5uzhuv3L
Qo827fmw0I5uAG/ouAuxIZbVffo9e3Bw+HIa7H4vSxzwheXZfRP5yv/heSVzgJ4sj7Q+HMtUxOWT
LuoVuTorSNL6Ci3LMbi/s67Gl9kY6/NuNaBCB6VtisTwXsaGk59w1wIoILwvzMP/MSguUR5jePVX
6+Fabvxk4By5p02pOhvyk+dm2JSZYi+SPZudscNEp+j9qV/VBKBG+BtOqSJnZBUZd7QgMxz87DSy
a/oq2TslCVi/bFv+mTJbT+FN2dk4cfKJQNLjjmJG+BUZKsL1vIN1dLPIEzZuE73tj9K+77dkh1KC
ykVd8RuvbrgekQ1752wZQX6IZLsUQKB04zO7kZFcKaVcOr2Nf3uTzSP2udqyBXLmD1AsCaqBj1SW
tZzVMjNVYPJPt8rcweucE2jo8IJAoldRWRLZdks50i6XaVKn5zlqpMaZmqAI0wHlFv/f0n7Ucb2X
gDm29V+TSx9w7Mbbfu+/QVj3NilJ3rd13OGl91GB0YgKl0EMIGPqGIoLVukGfeA8oPmo872opltC
es/tp+MNnin+vvTJ3ark2aqMqaqQEXHLzol+JPfWjeJTIhxuV/oPNVEgEerafHoRL1jd/tR/UKl1
qGsDeMIrQWuqaItVzzsC5KDJYK+qYMlX3a45HdV4YR859FEEqExDiUveW7n7Jq9/ssE//Umi8CaH
/xJ+uGAfM7kQnN6Dbt2dzZs6XiAOJGPBzkNJXKV2nunEntGlOf/JixeNVa2GzRi3GmwINv4up9U/
HR/Dlj+5jzqPp+WO41dLdmgiBaki4roaBsLjVQ9IRv5a5qQexxUESvh2kBZSnInLMs1wHziwbDy/
x/HgGMYdHw5gJDZ/BWGQUuj2t+OnIgktQOsl3ae8hW68ehLJDgAPRIw6+93HmjlfRXzkXABF/pUY
sHo6oAyyYtdyqIfdxooXx9ROxXVp63KhMM00I+lzV4BInSX0JJJkHJb293VsGX85/kj+NgVgkojs
e7WzKKJ3B4xQyZkmRi8nAEFwgv2oq8lBy5SIyunWtDU1kc3JqQ+Tzbmccg4gm5Mby4MIb1tyb25g
7fDXAgPOJnOvgakaNhU3Fzf1YS+V2RrW2a513EzqWenCFwxScUiuxpgXgRi3+a3eELXmNUPu6X6W
IBk/Y8uHfOruBlHCoMTABiNvAh0XMSCmo+WwLB9BHkXXOrGlXXqJKpCe1c8yR7cEFVL4wIOBJJHY
m9mO1WhJX6LlS/mESyQyD7gipVf19LNUQHOK+VwzLVlaAvq6qpIpEIWbVdtTDUaFrLbzsm456C+v
THX8q8EilJk0Evrbfj2hzUQvn4VefOuax0QSVFnvXsd1ZK0CxcYoXI/30AwVBxDVyIm1tcxUiRiQ
cdl+Z5c4WFlRrRbmoL1Fhd5xeK8Z70SnaNvuhJRigjb27XHrcJTwO5fTWDQ2p4cgNteCaJw3E6+B
RMh/EnBmNDWBUAwlnzdpSqSFC/uL1xNKe6KpjgFiNOgl4hUwroNB+J+R5iwdm8MBtUa6Wt6qSO+5
VjubSgqoQacSvHe8PwBCFy/9ww//AsPI16X3AbriOjgKnZ6MugzLoryM+tXY2ZEagsIZYUbZe18Z
LWolwjwupiXcG4uyJbTYesladjdFAEckYqG9g16MqvBGnZoDC03BEwTQ33UlOutPn+3iJmllql44
x7uyXO5SD413iLBuewGX+d5a9BF1l1WfHsBTI819oenJpCVbZAjud/9VvEcEtjyuzPs5zVi+mA/8
gAvnfy3llrMU6V31Rstzsz5wIvixvSyqZVsywnZWRqxrSj8xtSZBvA1e2v3rMoJn0DVp4DQAmGkH
KloQIyXDe3NIRH2Y9j1S220FjAatbZgHdekZS6koQAblNPlfM4fh3Awz7fJBOX2hpJviHg8UqEWE
v+ljnCyFw/HqKgqP1yQEEE4RvXYmPtl0lbRUWWfaipbWcaJz3Rn4JZv4R1Uh73znM3CtHabLKkMd
MDaOjYvVvPiEA0VmQRtOANZJ0QF9b/3FQ3QUjTD8t0kZas8Qi4g344N9XyWqnxhZTy5xqzc+8xzF
4As17m3UP9XUbHmvuGN8VCCWpISg6wa3VKNASO2U27puxrTsQc15a0hFpzdyXdZ15WLncsfhQfFX
OoMxpbJdwAE5BtnMJP8GiTga2buJx8Ouat/rVSwqrmyRleYybb4vH5jWd9SwYdT0h4/hodGyQ3u9
fhP5DuSY3MefUqdurWfOBWmL9ehcaaToRamGCatJfsouv4Tlbcr7ldgBDuRe8KUXyMZs2Ovichib
ew+XsOG0mA5mxyhYoBiWp0EHTIzKdM0NF7lZRvC5kSiii4VYKBSHKE+ZZbD+bACWfCC2RLuXF3QT
J0RUjRwLIyWbKlSA2SjrP/w+irIsiFeRg5kx5+eBZtSXzFVLaBcG0GUHaWxyyu7YuQ2ZE2oSfItd
OTPbrycQjTFH11zOJdeceZaWmCbCBlDdDqgqST6iKpDsZB53ic3MplSwyDhz4pxRE8jUhgUuHroz
e+HW66yiJzX4lRsq2VpLhT7WoaxmC+AhqjiK6mtoN3km3+K/fJUAv+FZFRs6SXSq4ovOXBh3INu9
FiDuNImScmvk3sh7Je0qWcIpyPgAcvEiNIHWZ4rMIhYf3DeU+6ogm1Lvh43o3+hkWwqr+QtxNaIk
NNzqYy78/29Pse8t2TXFCF6nNTKgn4VU3MwjTduOVaGEKavX43qfky6QhdElVpP355MkkD9Qh1XY
ttpAbc1MfhTLPXr3S64qfsDPnFg11ix2XHZJdsXqESM4NoHvGfEKBRJrCXDQN+Nyt7QaSO6qQUpp
AlCANTypQbMp998XvdYdypwW5dEKvLcN8pDF62NFjKINmEKI7V45ZMJ/CDkNKHdbxuuzCZZjuRcv
F5R2uR6GcWj8mnpjPuYLYbDj8Um8oeXX3yhetIWvowwkPi/n7K71IWQffFOv6loAB/jOb/xu71DR
8ClC2zzdk0Xz+5Ak1zfFLW3Ym9HjRoSXZgW7UsYx7xfY4gLYdAWJfZ1aN0eZGbT6v8powXgZgtHo
SX72kv9O+fep9Tqm90OX5HwPcKtQhOBI4mpCjlgXeUnrOWy5UxLvwNKmBsNjrUZSS7JIup2QEtjK
WFpwrFdoUn6wLA+QmkHY2PKq+qZhzz8yDoR1uzXEazyUc64Q5GXdiqFaZckgD9GUVxXcBCv4B8Cf
J0F82fXney9qKvoFsj7nsXLE9gKhuCLgPcvnnl0eCHTlqMD6FmwqqDXOllBjp+H89SOvZ3398GYx
6b5bn1wiILReGvquaWMiIXH3zduu9/OdobMa+wnCpYa2n+LINorlnaGkCr3xjpdJybej7wTVqy4p
HVJ6KqyKU5TFydS5fN96dzYnWEnA7Oa90J83JNAqT7KZ+4jCitvdRV0/ALC/9ZGtnblC/zyrvwDj
k2RRo+Nfi5x8X3ZdRtRQ910dMESnwGY1oV1KPq9I1OdXZrjJEFW5+flS31DgoivklqB1vK6yaMey
2nW0Tkf3YxLmCb2K4oX/wQb/RtxW76cByaUcs+ts0KIxCodXRBZc8pIYUdsnk+5IwL76JV0dAgVu
df3k+K2pU9gH73yGavCkPlgK7+GBfdmNOhk3Ig4lhGNXmZ95f/0QmxBvMKtiwYHiKcW5gYiGTY9d
TpVxBiwSaUlt20PulvYUJ9+4wDwe4iEa2f6fmwdEweU1276hzqK76PT+TjIlHDEUCH+p5ZjUIuG3
8OtQlE9lVaDNJkHzzn2cNWuhq1GfcvlDzFh03vTLeRNo0ktpZfrvjhhTQiLw5GrTuGzW6cLUtMfj
z05e8E/QGVJKwsRiFDtornQ61ZWipagxgrcBBxc2ijddGKb07B631+LtSAjWoaAXeOs8gKRFOqZu
3foSJTg/cteBB3wNgC3TgLaB+mgobpxx8CK3NHStbTIPj74CBpkrW3o6v3H3F9ahqxcQWc/tpj67
udkovbt1DU2fDeNRREvQRtS6Rj2heQD+zmWUMYehXk/KRxsmhlUGkzC9jzW01eLy63EwSq+Jx0WL
8uQE6qaIvNZMyueJL3od7WC3Q2g+DMvp5W2rfVEsGB9v9s/C6iTe+aTL4m7eI03oWlyQZJ5DwzSc
cxoz0mVi99XLuI7WdPX/NZo8aRWoVZNL3YjmRnucPw99saSXSfHgldFumiNPqNfwQnukdzGcEuJz
9LGdAv05yzcVQAveB94tQH7QYoq3BOIjDwqhPAZsdDCs2DrQNKRqJACPsv4ahJw7cG0V0qECbJl+
Zr65rhne4L6+rLNGjMUYWsLoQjLQYeVFp6t4hMz0r1FBqIHimRSqqUXIO11zHd4ReMI6O4JSvz5m
dtx4CWNRQ12WcxFTB+19Eze6YiwbGZ86+0zUHh39+RalkweYqSn6HBcPs0KjQIzwHhGWGY5jt4Ca
ew0rqKXEP2OCm2fQTk/8d0I1414xQEScZeVIwsP40IzMaT/dy23TLrI4gQ9rzObD5oh7rvdBIoXI
aZMGRfEJrjg57z9O8saTw+iZgkgL/U9PzaY/clPm1yvNkJ3b1Co96juh9a7m8uaEORXzS9+eHmVJ
pe6kvpk0XAm5bv5mWqc+PnE+KvSHBDaXybmnBZD9qVZIkGAoIlR8oyWZgWJqYfX4Dk95BIp42wjd
7xyQgfibItD3Gk8J5R5WQhleL02Dak0Wa1zGQ9nEeB3/9JjOqFO7wHP/IIA8kGldIkc9ZQBiRVeL
6ud6cOjyrfJC3aVn2I/P5iNUCZRAdX9WvTDQUkJ1Te5efg+1LPjuEBBQ/N6txoBFdepItmsSwkC/
d8I3Q6Cg893/OjQKB5YkOYvPk3/j5wqUEMTKZ/8CLWqTzjTXxyU7OFVu13TAesldtOlRhM9+yDbe
FDbpqMWfucT3OOtaXZx1ixuHptrnzT8ZKelIHzKZRlQFqS0h+Mu3SeuTlQIoK1g3yYSBWXnpsy34
lLN2CMArLQgzQxQ3YjTQIz7SiSoaFm1KFRz/ZcBDC4jHEnxJ/FRuxpOehEBZy7t0SMD4EmZiCzBQ
UcLm0NVQ8jYC26BEzwyzPvZc1M8wjBdws9ZRdJW7d7khrHS8j8+tl9vS3X8RcAqvZz31ULJuDZgC
60ZznMCPMxayWfVrzhJfsHWbGuEE0EiZQn9Gf6zCzKWhxsqEPQpc3DxTrpkYR10Nr2vWvNcH5XuU
lQY4joHc12PulsX8Uarz/tscQs3mrWDzI8rglPX1UOQAjtzw8llDfs3hzNDyWDQUsiFXwi6Rn4FL
WRKiEy4CHO+cgDfpbB+jZWss6KBjINimM/xjcJGWT0I/p1GkYVBBZKqAkqPK6Y4S6HJPzSXau/a2
P/cSSFbssZBIOz44IeGYmU4G/WokyfJdKLbIuAAzyukDlEq7uhp5RxyILVO9KU9LGsXTjSPAiFEj
19o1VL2O4B/d4pHGjkfHt9UuhgjedecS2e3YxlMpeK6MMDCtH98ULP+BJdcIK8Yec/iPf5L/qChx
SHvgnPgXuau9o2nqIjy+slU/ucvU4XDBnWgtiGI48nz2PkQpjSlJlgxFuezLZ73XyvTccrKgkui5
7dkGUbfTjr39v8OVgf24/+zn3zZAwjaCW3cGcaQs0AoC0DbkE8aP+d+CTtaRahuSZ6Ntx98ecVnt
IBB9+SzJWigDsFb8x9k//zO2oa13QkqIW/2caFbdfq94DV54IJCjaXIrD5NzgqVlAUNcgVWS4seD
tgDcab48RzEPxTYOaDKta5kZY6ChqrApwZDOc8MrWLNdwM4O7uYn+ZPaLFGmbQQV51OefsD7kqou
vnmnB8K2qevokWb9TfhpCnMOxE8B+QJtgNtkrcb3F+6LchZQqAi1gUB+VVXmsZGd4/Zws4sMiAMr
i0qQ+Htw+5qo5E7CpPdPu3mW2co4yho2OH9QePelnn18HP621a+cvGMUHMe9Jro7kmFMVMgy+5um
oyHd7q8f5y4/PZ9eF0gUSQ6jfOJpitnmRXRDqdsAw88uI5rWQMopuYPM5OCy3V/5Z9hYO158l59q
BlP4hid5H/IeiwPwPipxlWWlrzDj7+LK/Sy8ngR7Qu4na/0q6l/33vDQ4x+KeIFIKe9IE/2kKdDX
SZUN2TSuydeWpBb/cGYvzqdHA6tZj3IUhtdkxL8yzW/7cEoVmlizRHhxSTdbkk/McLtLt58sZrtu
Yl4pKL3XMz8dGKcMu7sTxz28d8+CdaS9rmW1Ke3OeV8xZut+ntlBTHbeCqUmX0GBpkEdN8CJ4CJb
fIkfoctSLveiB/1F6EeJ1sLCTntXRXFfQDk3d31jqFMqVFWqTSv8xaj/fXhEZEFw8hHovwesFWqb
qyrr8LD4QTFmKklGj0voHhB+0g+kq4fSjjrtEbz2dV0JHc0eeDbLwDtBxbXokIm8MYcAKGcoaC+w
ztEhYsCBk142Yf6aXiYHfvgCcTim+k6YTPn5KKh8nx/5ZqDt5jrahn9syORTfmdvUjCLca7biIlm
d8iwzGXtffJ+AETukmGXZ3tdvIOlImdsf24e6R1pwPMkOvh/m50KMQiq/NpXT7i1HqJgbVBCWEJM
eFvdclUVhKJWharBIFFHlN65D/CXWJUiz5dKmNxCQWNKYSQvc8YNRkfNkm59g38rTt3yWYYrhtts
1LZZBkyNC7dA7UxS9+tBjLrlgznSDUNLJ1CU442Y82Ct4msB6G6IsHoUeDDclkUtFuRPN4AoK94v
kbTllaif+WRsyo6SWsvtyX1QVftvU9OJ+3fHmfZw/8rBCqFpH3hUGBtRLXvTrUQPR4t6C3wSrOZ3
XxgS65hXs7zW63P8F55/0UID3omWwynJasvUaT0LDYdJ6BM+4LZ/wuxibOdnoPwb+ViJWgtj1Xnt
xYb67kpSrkV/rNoSGdl0VtHlkOniYK9A7yM72d+CJrynZsvl7Y+QDPtsVkzUgIPrHsRiiOYr09dt
NnXm4XAGKPaoEUHa7uMhidCdJD2vHytDeX29Uyf6Sa0TSvBbOIJd2QIWoIuSSIohU5LV2/cbaxpb
Tkbh//kI/cJ4UnIdA5JB19oivsuR4TyB2hbJmfri2p0tBmeOLiS6lY4w/kj7y987VwWz0bIj4uin
XgCKR5lIOx6NPTlnXV+9hUOO585Y1wwVER8rEUT2H57+yMQ6oE5Jcmbp4OlDpQtUyc+5jWtm61dF
2BTHBBpTRnmNBu0kL1gqo8hAAxhadvw79VF+atcjHgjzQEo5TxqumNdtb7En3+wgWUhJ00PEYRwH
kCvsta1GYljIaQATUyov1/NJB8q54S9QxFK4GN0SFBWAy3NcA/2fP92+ntJN03yJzT/+X7mC55eW
53FaFirwJhdrL4N/gCNvHxXE9TEVMd8popH3MZAiWc2JVGszi43qdSlt8rKR1YuIghlSfDqHU3CY
wx0IpXYEJZe9YxSEyyHFMHPHRWgSQbokc5WvpgiqWhCj1gN9tq7emZm4ucOfeTRhGZem7pE9nlxt
Vmq5frDDuXc/9jHSKV3EJ6uu2bBMFBUo0KuyUjwoWDjL1tMjJV+QiR4AJdNCy6x71vIO1jYfDbSL
rW8FrrSkT4vwicHdDGOJd/jeTn4196kF2Rcd30R1G2BWAvZdN2p4f2sGUPsetBwbABPEvVa5mUOI
ClBqkU/BR3Uzb/aK44NvLctr4MsMjPgOEAq+ZGPb0a7Y8YVyW1ZPXvaJ7UNaxM11gFXyyTSzAntr
tjdjlDapog1pZNuCjsZ9onuHtVM7x4EtSy0YqDlNXj3GpmaZQt0R0XAsfUisFB8ss9OOFjp6HwPV
ZdTrmm1g28+RcPP0JHcadN3R+DaYQOFiXnFe6nPDOSIoWaXGUIp+FOpHfoIPeIblWYjAHic5irbj
qZEN9zMOR+tfTjwv1urUn5lB5u30LdtlRQ+qtvRG2rpZi+kuXTO+JXELhqABx3khgVxFrQYLYxT1
z9dvSvnCg7bH/S3Nh/RGi7jAZ2ao3bhQG8WGNzMUEb6Z2aEe6l0+h8inJmtjChlQ4OsoPP1dWGxK
9z8exsVuDGWHUFO0R1aLI3GKCxF/ufrxIHYrDwBAcJzaxT4y7YASk1euXMqyU3avsancjBWXESIE
JVHsEThXgVoq9oOlhT2KSxFWPusGG2T2Zt7sydkc99/gzX0X8gczdr5HVx2Vp5KEFkB8vHpwaKI3
IyiOB5tj04WDehDagI/q1V7+BOWszMS0pn4Xm7YW+ulEMeaPYn9h6qVJoOce7dRiGO8ktz/jnpEg
awsrIFf8wTmDnmG1NQRD79YSkPGKNcyqP+wfwYXJxCfs8T/goPiedtdfG1QtYlVGnPyXRfCMOeUQ
eROycx0cboiozMSMLrCfSH3E/28COorr5AfHhqDvVoko3vPiUOedEEgv112idgQY4QYgTbaq5rRl
vTHs4wGTSuyOI5ZnJgpfvsUZEANX0g1AGKgom/gceRIi1OhSbOlwjKauj4IHpsvldy4l4tZxp+53
zHo9zERX2de1GXJeUaCd0KHw3RkXvSrUCTQ1wN1hgo9no/iaSm0UOwxGBy8CDMNlUYwOf6WKAAax
/xm/YIA9clUVFAMRiIm7ZxT0rS4qvwxIxfPrMtjavTbk9s28zp8HbE/23pdoDnFygXVuUtFHrElg
KAATyOT0xgdUfqIXtIWQsMm5WT4btZdAuk730GuEs2MH2Tw25suhbcfOOdz54VUTskJeU7K19Dd6
iyHU9RsMjske60gfuR/J5BSYk1KIW4RnglGyLZJUg4iGUQJNb0PBgWao4Otm+xVfNQPH7i0r7K/R
NwomQliYhm35XyiRWtj6jqEG4vQFWFTYNMoQ5jMDXw45yVX1OYkYMn7Jyd+3g4e1hUP9r+Nn18YS
wjo30z3OrjthPVG0UjDqYEiZFZZ4THH3jMaa+3FuvTH1OeQZ4SbwbE7fDxR2RUu6rAspavNRgldn
0LucsimWBP1SrWI89wk8K+xLmO1NLP7dY9D7lgGwKKWYwe/Sn8DMrIA3/JaiDPE9kvTL/DJPUg6g
xhrra9Ao/en4irS8NLFmVC3NrWPdJrBKZJXf+fUHM0yz+2sp9UGU2CnmHtMAHBHjps8OYzBpsaNo
PYY1/e04wYXbJFGENv7F81SFObimvWYBgJkX7ZMZGWyupWPe5y2/o7fz5OqWOLCSa8lVBOiNS30q
fKAONrAykT8mmxi2xhqZEJUx9Ry5R7m3+r0BTljBo20JrBiilkusd5znG8DVQZ7tVxtE4bd3WvmZ
4N4GJpHz7cZt/dkI4989RoEYvAB2vyoqNZ+vvDbMMH4bYN3felcCPIhWiRuaCnFq0WN6Xvl45zQM
7OTwJUZQMbxhhuEA4GHEnlM68/hKcgLIsx2qtsT7zoc0RDY5j2FWFJm7mRqWJa83+qKhE9B1Zz+4
FtPql+SyyjZn8+G/RFxgNwE/BHShzd37hMF34eV/8vub9Bpf1YMfVx2NvBUYm75jePaRCUbGZrca
UDFp35V/ueobKmMqAwIu1p/et6bHS9LPE+0zBWXVUjSCYTl66KRTQljFjUKEPHG1vEnymTQgEC6L
7j4C4YqXjDmW9+63bcKvguKFkVohrqzrNngWSBPE9Mmioqg6QXdhHrlPDXlyRcOKARc1BFceS/2c
9S6f8bHOjoyYy2aT5ENMcvu/juZMGLu9J+BMhUa3OVYiQ+CmmBPGiqy3blZMF+ENj7A+49QawOvZ
G5JkNrFUZi1F3zaedsiY+mMm1APGGk8Iqr3fV61rCxtwev3SernvaXeRmNoWtJavIAYwcYRF5lkg
Qbz8KgnBjV9iTubsBJxryNkhamyixV5K5aGm3A6WIqT/aVZKLNeF4wtwrPvzRZ3Cj2xmYrqAEQEG
uTCTX5JjgemN2o87W4pSMbg+d87G9ODCBmgr8c+vahbs29blrUpUVqxpyFdT0Kvg/jbpGZKYDvn6
DVXZITKZGgj6T+5luAdBRenDdMAgGykXHWjyiyV8v5xPWtkEASGq3dhEtR0YOkuBIaQhNiM0mWqS
b4z2Hj+SED/x96fVGazzwLYwPWvVguOi/i0IyR0gkRIu8PySJ/+QFUJM4H4/lMpSon10Yq1aOXlF
DzMK6iZHJsJ6TNyEXE5ACjhkS+RFNESINGeFSWYjwZQE712zghKmFDrylikLFtBvaQv4pZ3E2isZ
uVM+Xt8Bf+ipjl/n5EodVMtPEGvEV3NwKbUntPTEdeKnEKE95flzZ1pIfLxviEUt0CuWLRH/voVR
t91jNzch/vLM7f0Uzy/wmAGL8+ph9Pz+eC1cIbgWsCccEJVGJbIj6LZQbADWt52UpQlxIwgVhN3X
BF9EVSIxcCXv7iqqRHijl2JLQVccUSW78JXF9fUVE7fjKnMjSWhulbX9/VIfbc+ZL3fT5V9U4q0d
zApqq9Ji18aK7fR0OsOm+GOFQjFTXdmscDivKSunzN3nTOL0vyEYRnuL72ShYlkqnzgwbTiIa9K0
bH9bj0wxhW6l20PEvJRyHuW99hq/EZmS4eQ7i6CV8o2070Rldp5WqGQZVhSyd363FehetMVRiRbw
27wckM5goSBm+ukhL9+n0OioPJYnvDHiDVR3hjfQJ0cMTo6IbsxrTp1kvM/82Vyt6LJOxKnF/KWc
n2pDGPrdlQK3epTrTnJkNd1mKNYZXEg+RPEqgi0X92vm48sv4UHvvIf0y+TVMqL/lr+wEJxIHFSY
Nq11eBTZw5dQ6abz7roYU4SJt3KVg1Y3E7fKMTEb6cMpoJy+03ThZBfnmCLo7OJqQs7kbZIyMOh8
L11BLdhtekSV3Kv8bBgkqzFBD9V78cfJhKFc+39zwX4Eh12DmPqPH1CF6qQNBnp6Z5viFqgtHQrJ
71aHZX1BroHWPV3iAwM2JG6W6vlmkRu8FNuV5BqfLWTozuLJELGY1FOKJxTubfcynlAiytQsmyG9
6eRhMQMl17h+YKmMjLXz3+4IB/X2OUq4xJi9louQM1grGGt3d1vmoQP25aQ8ByuTSJ1YN8mj451r
D7158dK24eHDXXvuVqaBSEETJ9dkzkemm8R0z7FfmVgJvlZ+U4y4wI1FztJ8PKSR5rayt//MGIz1
d/KRQR7Hk7bDt7SPSO//Q5sYKkLwXJvMglgtICcrPR5uGwmJMU5GMTVoSZn5+uJSoBA6OPoWT7MD
3qlkkpKS9KuiuwiF1pWr4qbBkpqfgAoRWWWN9038eubtXEacPo5EyDWhVML4jucxCczZJf/19oH2
NHaKOiTUQHSLfELmIzphkzptaglVBcq2TUXQfB0U4EApi4AEQREimJNTzdZmOjBlBe2vGCWuR6wl
69CJ0Q5XrlWz4IvnpU5xODKIP60QdStfu3HV13xbU3IkUMYzFS6BvadT/FjfkPnlyk60jmxR5m9d
AWyc9Gr+E5mUoLP5PHXeaFVpoClT44CPtdW+z8TSRqa7Oo+CwSNW3Am9iHocI9GeFhSNXDTzqBqQ
5YLxNm+BonYhGYMpoz0fVmmb6xZBr81tU5OJjSioh1bindZ65lBL5JX5b5sWPHoTixft1PiQU8W5
Jw1GVo4SUG3M8ednMGYrvX4ib1ncoYUJfxem/gqA47NsiJhisJcMXFJ76zNyAPlMu31qyflNYgVc
6Ew1PwB6PmJSJp5VHFwTgkuyXjJ/icQA0vK4RMVYcTpxsxziDTRKmWoJRrrNnj3jnwlwBB8OOWwx
w07Jrgi7y+X4r+mkL1g3LzDe2r48bzvfIuQXt7W8tkYRhUzgTMWmJWYjZWg5XpXbkymoOaxqqZqn
qIazSXjg0muc2eJUZ3lPKVkcJF02j4G/rEMxLHAinc2xh0kPcHmbTZSdHNmRsnfLKn4cxa6G2irE
ES6M+TYFVhRJPQIhM8PThQ+9NNdoQYRxOAj1BTqAWmnBD1AGy9xgA9/CcbV6L30mNAmRrDBusLob
b2q46uFDwzpiI1bQHtY+JllMH8fMKbEVt0KkgD6enVfTE6ds7LwOg6BjAke2oEYlItcU8liAqdhu
3xhdkweaermwlKDTNklrzmCtkxvG8ncN2uyIZqP8igTrRFWSREwHeE9xgA1q6DGNNAN0T50xeDMj
AAKRUhyOwSnGwzew0DIVTFbYRCeg3FE2th/mG/nZaNDETRkfDvNcX2uvyxD13cOsvukGqB1rmwCm
RF+qvCkKcU5b58zqP63vXSONfEvNUxGu0Gh8UkvpDBHb/1SA1q4yqGKLWm7i4CI/vwffO3aqECFr
3UOEJ1JDwmCGp/ZzAc+EUBe3wSPpPeEO93EtniE+DBl12n6mqqIPIWoFp+Z9CPUksiNPS5zwvwwn
jFtR8h5XjNpZXL2hctVfqCreAJBmupLMmlvViFmlmElLT+grsDT84ZYsFe4/YeaY8FmGqvq+JUZZ
wnupsk4/Y9H2TReWD8Mm95UKf10T9p3+PKARP4fa+YPp0GaQP3mmRdztCTROpQrntxiGjGOO6IzS
ONeG0Mkpul12zg+HAjxbLwk8IgPdz8mEVrAGs5mO/PWrbq6y2Xj4eGgo9jZ8XrkEXir+zsYxUdq9
znS3+gVzmAhpHeRRZsJ+CNgI8mWnEiWEmQCVW0jFgDbqthOd46YkOQb/QCW3K13GXBPuM7Xf9nlb
m9UfJOu6kBkMjArszhgOxTkXxBa1D8HAWHK6M3w0o3+gaooWps11Y3A6ZU/7xfd1x7N+RtMXUk2P
hz2uXv+eY2JMjsyWBiiOcCb9HahQEga7DDhOsege/lCCVSC+BKC1eo1Qv1rdesPzAQl7lCmPiyyT
tPvxCdR2FHkwMdxLyRithYX10fIKqR77szj2FYwQ91QFJklcUiX/o3fV1Q3AFmoBzDVVPLzduLLb
szQaMH4H54HYRNlD8QLtPz2Sqe55fAGbIYXep+gmO3YQGidkFCxOGHqtmbwboVTmNG0HcBkU01c9
rjRolIebUg309UwG2g/2YiRWDUYGUDSv7rGiCOAbygR9JjUsDxLizVtHvrnmtpPDTFiohYFjZtDg
q6+pat3Fhj3mnc5g0mKMgmXpZUYQhuQMFSYzXmXdAteqX16ZyFrnl7l+wyz08l3fAugWZa1lnhKL
LD60he6PVGTl4QKCuzbnThi4rtObc/Y+r11XRazgaD+3LzxNmcc4Ufr4KQTBWpgqnF5EUV/wcpRd
iMHd0n6nmybCe64ovjX3hgjcE1lOJWf2431oP5nF4FssbUWXf2amRxJsTxXTIeKxuUYFzE1IkpTT
kNrv6LNnjBT/jWS5EkQfXoYGPpvWlodPXh+FoZMH1QWocRqq1AvxJKOEtmft2VDX4/Ax5FbcS3KX
to57v6K9Hs/DH3GOAIKrAJoMSsZBS4e3YNpNNP1B9l1WdUki/k+QBCYjugEuG9cWB2eSo08BwMD+
DspV6NJq7qZ84gVQd0e43dg7RNTubphuSc43Ki6hpgfF1AUxupxjVbB2PVV1lKqsqwxBf25bQAYZ
k3uzMdH7ylLdJfzlWN0TBn6dLlVLCftxOYsXOmr51kYjcyYkRjDM/q1c2b0v8VcmR410L7fXv+dU
GAnHRxpUAY83VaJaTFIz6KYqol8YIsU56NI8HsW5Q4dkqv3mfKWj6V8M7DSlZLV+yR1yEiFjyloa
48keUmnbdxAoMREXQIjRTnTgvvZTY0FSeUdAGA/wa5GFfCiSnIMY//SBobNbGrIpKU7XHW/lZQJL
XUi5UaWeFf1d/lZT+TBgJ/tEm2FxSSCxucqPGjLrQ2O/ho5ZtuUkV7K4xqOCc5Fj9pBvgE20qn1F
UMNhiIkx7ZFEtQujByVWKjiF6tZQY4s8PaOtj/Oy/zGxR0WAc2x34V9S2cHgJz8+Ww9ZAT1gBY1t
ygrOEeAgTa4XjEmu7+3gl9p15mezlK6O+kJdfEDvBvA5eZ/I+el5zCKqAvXP/WmAy2eifhKRDwLr
YmTBH3NcMCjTmfxJBwb+7m/Z2DVMcu7nsfg6jukHlEZNdERzJPnW4/b+PeXfR75JVnOMPj4K0aSE
9MXe3vq2Y4pKzmvIcfJxa/JBUb8dYHlg07ahK/8ZV0A9li6r9eTa2wPYaMPTnJxcLApB3a6LarC8
T5h1Lgy0yLCyxs0jm9jz1Not+bOfOj70+6xmstfD3EYsmlFNmx47X1pghcbWK2YJZ0mCuOLJHCzQ
meiMgfJcAW2wIq3x5p8F8iCP5wgmYTDBxL3McsBgHOTM6NoS34FxVKumKzhkR/1enhBRcqPbY8aJ
0hai6sGGdZ6teGdKjCt0enfuXdNpGY0LUGM5FLKNIhD+tnDgwfTexd22myO5BSigDNRXURyklSET
pCFPi+nJARv+rysYMIGBMiaFSzFrrlII77xmfWdvqjks3AiGs58qcARiT10fGZt2iNyANHJH9qiA
Kv7H6PI5JI9JyKkNJ/jKotpxTn1ZxLYYmahp7NRv16V7HaJJ/lYRwGSXxY2MKoS1xy9RjcLBrXhQ
NbgoKvsqyfhXb67ZvnFrQ/KmbOrQWS76phNNxi9fJjR4wzA6k+0j3cBNtVb7eLeYCQJvYTqt7iYl
lBp8d3RGlKUi+gCSo2UvN+J/4Nq2ppvU8fOOhVe2pp5zw6+872Si1WrwF7QdtnmhYEBSgvEUqzxd
iLc0H6h6piTVYr+zgZX7Qm3rwG6B9duPqnLQoSXJy83lqtHVhlsZHVsHwgYWFzr7zhPu/sKZICbY
dNDJSZgjD6kWbNJXL8rIE5U23/jGa6HNqXhQytxuMBXyI4UzJLQuJWBqVELtOWPHaxAuSWvn1jaw
HfMQMvy3rWxl/KQuISOi19Cr9t7A+2NaJEXLcF1rwCIBQFQ0UjVl4ewln7Eke3LGCSan7E5CTUNw
Ol+JuNPzqMqiVgTH06nJjBmz03nFj9kyMwLRwy2pGWG/2VOvjurZZD+iaFbKeItbdCLP/CMxrLd7
TZ83aCx41VyBWzWAG5cKuq2Bwxxjf/BQ+hSi3s7r8aF+3Vv1rLUbgz7+n4Ie7fLRP+N+2ZrdOVuK
tfqxxcrJmp1ReGBwDeiA9m/K2LWa75ZniBXRD66hTFu3nY4jd4JGuTM7EOPBKSS96CSrHBgCXZem
lTDmMoVxNzMumwdiFjR2Z5/Xv/t/QQRo/dqUJ9+uN9EdEBo5qhodrSRKfy6r2WfVDKxIi/7w9o/g
9s/4Dv+TRonCmeZ9MzRppQwc0+ZtvOLJ/ZMl1g5iCpg2wE008gLFRFLZZG+pXWNLoX1rhLpWE8PY
ZLlfum3DVJ1/uKfl4j8jh8nriHIn0IEqttz97d/5xlNc681MwkotVRjwki8DsecHx9FuQLZUPOhS
gi9jm+8w31L3kAbH4Qc1rCkNimoIB5ozwTsZ/NPVa2F6VLoisYMYsOlcDHSp1Doa8NlQ2OOo94sZ
xfGPpbG3F6Vf8axBeU89FwRWChXJlD+QGRiLwPENpcaN1EYojUd1pEDRPJ6WuNEWUc+65SvjV80p
P0a4DJd9ArPCWWM2CbZJnfYub55mYmqJr+7o3GoSTWaKym41Yr/9MGi9PP2wKYGxy69RR7yweQh7
WFdCDAjoVTgh/eQtQgXn6n6sJ/uSQsdirVcqdSD9N9GX7QqNH1Q4ApTmRgwWXSNILD8EScWuTyRQ
f6aCaKe+p8/kz/Co5X+GQyec5jfMXCeyoK+zpHwx+oJ4XBfd36o9dfhM5/I4IFdGYTmIotGegQHl
Iz0BWax94rngSokzCzXiK4x0eSzsaQQL6YFBJtkQ93Ak7U5DJDo9qqLdVvYDXVgMlEUY7jyeW71O
s09JiE8tfsnEj422An23rAhaqk+MJdRxkTdCSL9YvV7DlD48mqhp4BAOY3GTOrlNp6+E5RvpJTGU
SQjBxhu0fx18/vKMgsNYoVkvMWgF/MwlQFJ6xP+5BEn9Wv502GqmIKbq3C5FBUi0pYpOsdDGhBJ3
Mug3H+dD3ySWGVJufd75ShUiIJLbAkN7kR7VD4j1fOYJ54uB2rTCM0preddH4+zfDDpGqKRcwhIQ
ppC2KT23Eos/woFtNLk0GZ+Y47SsQtm1JoLxhZj8fvxiSHeIgnpojnf4N68gxoT40cBxRF91+abJ
SgFMEV9SOR6GyqI5hJ/pFIMKpOh4Tptwv2cJQKFbi9tEaE0dvnpndqGfBZgDVav36kV8T4fkXsUR
oShHMBKpGkVdS7Kv/eqNAnrumm0HI/sWtA7EsBs0a/u6vRKtL6nEDbRiHh8ROjLQd3sVgS4bAVdD
UjEfxPovdBnNB+13HKDtt9GcQ3MVQ2Lv+sYk06dlQwzfxXc2Cg3hHp/4RQkTXU0ZINS3RlNdTyW+
GnJkXB4FC1HuZSD5GpN1zwAnu3QxybDuchsXaIOCc/s0g1AMbikPsSFwHiXtkTiGUiSDJbyopB1M
+SxKFf6jXMqG7ZHIcdGBHqd7qgfokL6v3KmLXeXEYZo9EmKYOHbNluLVNCBUFpVel1YAW68Z41Rk
3yvLMaGYrpE8mQ9CNEROjxUX+pi0g1rz6/ldKMrvYTutfPl7BbKi3r0utkEcyMUDASPVZ0h0DKSC
I7QK38qQqrM2bzr3EXCpMdLYy5snCgumTJJVz6cUBwaVxiBoPXPF46IKM0zLbyBUPwWt+HSXs+up
P5v0DIEo+c9f1JKLaMPNEHUpGOnGyeoyEP2XA+J7KOWTbbRAA37AYw9cNdbafuKvCdcHTx/wYR13
MUUln3PoEGTRbxfe8/e8WZUsdZSdtNRy6aA9uDH5yECdbf0P8raJivJ1mkhUxYY62Wdu9x8FWiNW
yep0nNIea34iFcqzJU3QYhQBmNJ6TA+PdGH3ANpOSciFmjgfDjL4lNQ1twAoYPazkU1Tao/mZ8CY
OQECf+52BZkz526e0BacVAzM3ycz4aYhSrY7kwWUIb7XR/rL/ePCsM/FFrbilEtgKSEBiKtiBN3p
Kn4je+YHMjKvLX9+sI6PiySJDfX01Z9GYqeHnKQgcTqpatcUhcT5Obd6kKiBnCF1PXlvze+o67wH
iK6/lh+h5Lb359neUbvGdZKl4vUvX0LGfXPYOQSJ5PMM+VQojPoesIwPoAGog8+EmNlEDO4xiAJd
8JXZaaXnvrtJODRmucl+KXoVvKDb7fkrMRsMSE2PE8KV9AUTG5/o3SBCPWKhsWsJw7MZOWKzey7w
tZ9V85hF6PWDEa8Zri73PhCYm8BxgL/I9Lxlqq+77kWHxA4aJHcBPsycPnCx425TkdloYCSS3qsh
eaSBZb45CpC1mqbUnPU0KIWOhaGmQlcEiJdXoH+67xqpPx+vCCB61gi0BzEgc9/fqNScnohhq9uE
1UkdzyVnt1yUQx77LXAoqd+qK03enriZLTwq6muSIAKagMXm3LMWN2y3ChdQdEFqujLLoJCcbInW
7jahHMHm/pH2esJdhflCdGmFf6tbqBMA/bV0dm5tpNsnE9aXGV3wbJJFOuvSESjYXlV6SsEqnqJc
bcapgnA457eWGuc4gW3Y5X5G9bGypX7W4OB2w39EKcZjnWhlHomDcobYJOKzHHWqNlblQWx2yCbn
zZNIw3ArJKVWCbavvQCICbhL3zEvKSAGpuCKTs1jcVmtsgKKKG6vAxwJPMHzNFwjVbPmwMMgSLPt
wp9w8D9Qv7TQAHS1H0Tk7lHKotDUMFRA4Nzfl4pOxCiSEw9QPuYZaVYQmqX8+gYAoTCp3R6rgbfF
epDbUUG5dCcU6DjALpnLgY7+4VgmZeKi7h0b5Ngx0ufT8rm4hN0KGSZo86pAxO4Xg9MuCXn1TeiG
Xy/+4c4nd2txSQNLVILWwC/N3PZH4ou0T0uQeRuqQigMBHkqtZJoSRinh2a02gvPXwLMbik48NY+
MN8jdBTSNOKDMZ+NHRklVezQUVT9j6rGGAx5BPm9vbttQquYYGGMukCDplluTBHjV/0sLxdyKC7n
i8uM7rvnmFvyR4X0dIB9gDziIHrsghQwAeuUaqQ0txXkQILR0jchtxmM+T2cNMDSRNBSg5wlxEsw
h9zqSr72lmndAZScpNnuh0AEKdxlDuufBSNHZ/gI5nALOqljxHBm6syB+1qBJJMFHq1bRL3866UW
CZQVjfNR4RbKRBJp1Tm6R4TCebyRiGIq9dYcHoFjt4N1sHZiX5W29V/pBafiKEqiUnkDBzZ/eAQB
PpPI7ihNTdSqtcSy2o3G5ZS0TUevqRWtnAcSF1z8nKfhXur5XweHbtFTnSVKQbYMw//NksY1jvS7
c7vNMtLxOIWV45PiYGxRKT/LgxC9PKuv/Sq74knyIKiUINVLgv6R4mKUtQsyDiVm5Sha9o/PdQP2
Czwz0+mle7+BLUvud68UclVH3lXGVnXncoZylYAcAMl/5rME18c/I8C/VKeYGjwo6VBp6D77PLx4
t6cecblt+lm7uDzJofN71oZNw0g4I00G/2G4JKE6ASTD0Cbt9CHPv0BMBsteHC9adO+fWkBL8DV3
nUAhEYySqwWVn16PJN9OdTxRO0SRaRmYLd20uOPVQj9f0kMdLjzwLYFcsoQbF9q/ZHIqkr3drnRo
lV3mOM2jfYKaW9lAry+QAnjFA6tbeLLpUvEgrlcgHahS99Gwgn1nJz9lGr1eVEimT+TUlmXqKfSp
d18i8oggbPFBVAeQdcA5k+UticjRCvx9yGCSjgJX5wW+mNyisoxG+DA590JeIyWnpFBlPsQz6Zul
FsbzliIWe6roQrZhVgydHr+nrDFbyAH6vZn5ZgGADPhJcJgIv5fN7DDQu/6567KMF1RqXfNhLmbB
Sw7X6fNGfujB/41/qQ61PnJtPX+T9wW4vPJ80jffISPufaXstu203oJFHTVImi5qotUGF0aluJ1r
n+j9wRROn9TJjX+ZLmRKcerMefNivDbR1SpPb22LCz/pGlR0/S461YbRAIp23n1ubSJtW5FL6RWu
du8REUQDQGz2o4uUKvjnxYsVj/U6hdtj/5b/xe7gpUsBYEn+t6qksOmor6GK/P5jDkhYwk2euWOC
NDBsFPQLbT135mAsHxdWV10um5BU9MqYAdYX1opnu0HNey8QEiEZG9c9OfFWLV9p62No0dJsqF8v
VRGwadsT3pW8nRP9B+VGi2ma3K7ZoSMJlarHIejIYiUp+kou7i780Np/5ktUDiK6CtP/CyF17RoE
EasJzexRYJsw8I8qo7I9u9qNRT3gzwD0GiZK5RV7cZtuAr3c0X+uOEGbX7Ob4Mk/TWX6xXZYc1Mn
zTURdZFEOPi6Ludp14kDxQ2X8/ZU5MoHQDx2+yz6h++0Reg+YB9DUiOgDzfxWVrwavD2j39/hNdH
ksvzpc5kEcmNdcHrzeyltwlrrjrsu3wgt2OLWsILPHDv7/A6KiwsA9u71JZzuzUaL8aZbDn/PVEe
eEIIqV7W6lR3y78dPXKVsitPrWzJryqHDgApcLvHyKBcoA5TG9J7zMxA5vdEOE7indrdz2X+FegZ
d+NdsooRMVCzvSQsNijA4Bgc3O0VkHQLs8KGkSYpB7enhFZe5i7AsM7V3gLKTYdKgjiluNCI3HHx
keN9VXMkYSJfGvbfBVgPfAtYx4VplJJVK+R3PARpByUtYP+i0yk4t1gl9eGiUtNbOIznVsBa+fJr
rG954FLJDH81X3kqNMHJmM2bcdfBSN2wOQyR33qsCCkwEs7yv+faqUlOFgH5ua/HRwwyVyraUq34
ZLdtPlxMcD+gcnYsrB6mvzf6RbsD0lzJiveLiAcyh51EpufLg2tt/0qpirhzoPNhKeqht5kDTNlQ
t10HTH2M3vB2YYz8S1mNj8e5fOVcRN/QkxYyfCg/vJEG/mKRI6Dt/tHjPEAgN5gJZ0vz18hvT2ii
KB6s7xmsEs6bD2XDoclvro8bXNe5DdWho4pxxswwCGlWtnvVKDFzZHgD9kqFK6I8SGQcoMFTTln5
vr3ryFvfnfbM5wGhH/ZeKyAyZNAaEHZdScX9WEuiNVbjOSBTyiBOSobw1c3Fgil48ukjWHt3vvpz
KELgadPfo2iW0K4P0yd+VTxxYbX+9X2LbIJGB4iHsMvp0bKeOsdER/F0OnzUBC6beX/08ml38kwQ
lU/XJSzZiQnj867hKcCS+3wY/Q4vRI2xgCJ3a0VldEQIfGd6mlZXSbnKAOCLfztax3vVF1W9tiYW
cbzypRMF9bHyfTMZxn92q0338nW2dexgv7hXFeVtODVg23w42++VsCJTksVq6QS0ZoNYrjuH6ac3
pka+4TC9G81CxRZNWFRPOVvQYZmcIHuMMFgdI8Nq6Yt+WtsKyD57j4n4ig5Cx+prU+lWs+/GH8Ai
rPiEEawIcEkeXHdYhJCWg/iny52BdfpeWwpIpykUlYFwx/httS1GM3iI6n7zJHt0vVb6PJCHkWHT
w9jHzV6igByzU0CbtIutvf+89xJzXDmq/jdS/ydQudjcer7uxXYeRPikhIN09JY0GeMZJjNA4/gg
GrBebo8KIUwMofKWlygluFuN5lI3k+g1a9c6T/M7lmhqxkvvvH+Ui6cmiDgnDgQ6Gb0jyUXGawEH
lLhGn0vaf9zv1gzbnm6r5b42jPlmZd9IXMsuGHegBa1XRC5JOVNABjLcHqSd/bWJV3vFBCKd8OPP
Z99NaENdPDKK1+C1FWLwV1KhuRngHUEmUHFyu1IbhUNbrjh/baX7Z4Z7uJM1cuusvBdC3fZ2FCWV
cuvLYUaEFY/o71PnCVm9mCQLBdfFhiczcyqdH8NOEZMn0lrV0gor2OEQXSw2eB+smqHdRgtz/aOw
eREklcyeM3+0yP/R7NV/PDmPXletsSsV3NK/MB/WFZ8PqyIPtTe4UpWnVq2wGiXz/HSmIt0uop8U
uA88p0N+Q+6oF4Xx2VCWRdZH2GRku92SNHH77vEIQmBuCl4ZzZkZheitGLbguIAcmBIvHYjIFjRl
XTNkKNZdmJ9U2QG4/kVf7WT4lUS4NJJka9K7zwKyoj6c7J7HycQMCrTuUjBoDYxNIeVLiOlhI57U
PKATp5yE61Otv4+pYzRMdX3BdgyHz/4wSkJR0YRvnM7KF53zuWoCKD52zLMTfST2T2Px3UXlWfn8
dWKLpyrU/NVA7U89xyWkgj153yIfry2Wx5lfLrTsXDNJYF+TzFFRNsZEOqrQLE+OwGx3OePXnbVy
xVXBBaIa5hNo575fjqbHcCMpo+kPAHP+TUR8PzFoyOXy+aATj1+/9GLhc++pKuafxZ8h5cITSzxK
4xVGxiHlN653SaVC4HU8VgQMUmdOb9XrD5jxb/yaKbKtMb0ZlYkUgzC15lNGFVObGWZDxIOWdeZr
x4XvwYVfNCJYWSjzE6RkHk5ip9chKW3z6uC/fkuWEi/EC3FgusQQwXmPzsACChF9GW3jd4Mf5TJ6
3I+s4C9WaXGdc7QXCkhAUt+xh5RTchEEyX411SlRHqTGQI/22XA3b5WzdzvFkrqfDOIRY98lFTet
iTrGVm68aS+tl49sdFjk8/uhQj3EEHYql2tK8XvNEYC1W0On3ej8XN9dBfPLu1Q8sKYNb+cqM6Ya
r6oEWmkiNXJPCpQQ55YtmT5WSXYt9mzaYR6rGI4GLxDEXjSktyULp/G1veuFjvZpB5QHFDppU+my
6plMO5ODbymKDWIx1Fl/MJojzq6Ro2OYmYtmqkrXUgCgoAC10GMqRLf6kI0J70kHxph71rVKYvyQ
kxEZ4BoGonJ/GzhNuGh1TwRFvXakUcNpah8KzwGZPf8CLhXmGql09lRHJtuG72Ouiqcd3whSk06M
uuuNv6tWJG4agmdiNujintXEopd6J0DWCP5pEE7b0ATGpfqaU+Iz0lJIW0dNpENNkRynfTyRl6iR
fcFB8SMa+C9PxOssCZLWTd52og7HtdVgBwq+eOeJcakQOZVd5IKSvfdQvUeuwaoyYQd0yVKDgj4x
E3XVgJkPK3aX8IZ4BRtLV4e9Wh27xytrec97SsJDo+IcZszKDWdyPvhEx3vlJ9daWFD/7M8eMtnb
iZaE0EXy78NGzomJLon6RddQe+JpvCr9n2m5iXo23L4uU2EHL2VLCpkPoCnQSscRiiyS7oD/OLlQ
8h44+y1YuHLZt52iU+ntRNSxtyRZvzIZ98eri/c2PeymJ5IHrRP5bOQhvxtfsUSgQhhQWAen9/fI
HcrcheRhCrdKHwz/wPye/fYM1YTK+UJLhV4XmXvzmQ4Qpdz/GXfxUqlmEUw5+f/6+RGjhQAiFMmM
FHPB7VtLjK3XqKjSTfLbtZpa7U1eFchii29wdvFA+sL6w8KdsJOfQydmdjSdNceOiVnOL7Bbl/aP
jZ876MNDyajx+/StBhnssxv0dZ01TKysl/wrDkdFSCasdJ+tCpw+5JNrYoUIKJxuw8F72/mtJxkx
JH4+DsizwGCF0q/lmA26WSV6LUfxzl6z+KcVtkYGNu2JJ81WLFEtydi8eLGhrYJm7Hw8C5iQnnTU
LZk2QQc+ePpqHPLWH9pR1Wuo/GV0ADZLnK/7+RKLEE144gX3SJiScR/QhttqoFBBTGllN+BGqhWH
vql/eJD/KoSaYAdv6l1aq8fm2TbqUc0DOiJotm1BzhSIwzl6MkeBTujOhMyAQKf6UG93e5lfRsWW
w/pZCbRn2ekEDjiyv35uuU/RHbzzPNHfX92g1x6CN/Lt52cTHSWFuAelKdc8DyXJkrmy8ZeOi+r/
5LX8oL15AH34JWJPseR/zKCNtsYpJK8/0XEGHox2wIElWIplaVxmS1YMGD5KxfGekKMZZ8iCe+G0
Jm9L9DmwcsoYQ1lX2vDgLaB31Oxq3DV188PrU1yww6oXh8wvWU72RlEJxE3/imiwbOoXWBis/iJ7
Gdy5/kPGt8BOipx9RRVOwiPj4RSicf1UMSoRVNtflzVg4PcxsGyVpKJyisGRkIlo2XCzwrrsmaoP
7wk7AROKvSef8h2yl0OkJzaMNmnj3IgHgnLoWOuKY30zeRaLOfaR3uz+fqXI7sStd8g6HSYTlzlg
0EXanedG6Uy/s43kryg3CihehZHofpbLBR5219ztn+kQqP/iewMUWBSCh7WL7Ucij87EgsPdHKHg
/Ww4Q4wRx0ZDdANzyKIx0QSeNpyKZsxzkacGdCnDOG1lKyVYDbgDM50fZ4I7bZKJtL6b6qwxwfEW
MOSOgkCaXW5EM6kvTbSSc1l4BOGqNtBeDm9WdWKX4TO5WkL37jBausjIBhujn6p8iOW6jeeoROzK
IGt85nmORrDsOcKGokEeN0yr72eiuhBJ/aP27B9/fvOKUl0hFHlzSni01CUDkXcShXZTRdbyZzjH
rszpezcc/vkpP2Te55keVJsqafPt7TnoX4UrKRShgtvHpfRAOUiuB596aTHa7ape5XuVm0FvOc0C
RA9XJwYkMzNm/DElNt9Fa1AUS8U+B5HZU27QEOS640iVWR4nVoN46YAVCRyL3mTCoZCDcZWJyL6r
chBeXEHh7TXdgSl8T48UbrthiGhj89bW5aV+PEM55Awjk6mSqOQBSXhyTV9rLUNbh9FBVIuC7BID
A2E7XfrWzdca9qikAIVT7uWFAwrU7vcGKJX9zDhziDdx/bnMRQG4LHEbbH3wAg7mt3uBZtnWUdKw
RHxPPar/5pYA3SHCrdxSfLyLpjDplcXSSqqV5dfwYIpaD6QkbBM07FKsY1FhAWeB+uoouqj3oUOG
Pg903wEtyDKYIQ/R4tQrHx9bKJhtUn8jP0dm5nRvq6VYeGnfM3SgPAnOCgh1rhwFXUy2Oy3aXTrM
qk8h0n+vgTWOeJt6mVFZ78ZxcMwsJ4EbmOD59Kun7EtOEufcCROQwCy3lTd5CRqP9iOrHaAxF/Yl
GUKLXYZJyklXsZKAn20tT/01+QfSFbv7BVfzXjDVMOXInsyMJsbb7tWcsm7Vt1i4QKmRhWQut8Nk
jl2NHw+U4jdG9b9gDwGtvqeXPm7n+I+OYp2NDtIBBceiO++eGXBcEZvSG3TqUWV7QYnEqCYQdNM2
pgKS6nO6GfTHzYkIz1/YffxP4NrKRZ04HPV3ilrDmhdUwPIioc/9CZkL271cIEG/igxPvHQV+tpU
yN+P1zSus9FLWoCMpXYmkjqbL8VFC4WfQGqxDKKsC5axaVdBPpy9oIlFS52edvJBMc/73viOKpA0
QSs8PDcWq/T0vDkGP1htQXABe97yazfdItrYHEeABzbNE1+ds+AaMaOE0NwqVxrrIe+qT/itbef7
S9ff6MWwXlFeg7bUec4xCdS8WcjN1SX9aysfNoLGNn4diZ4R9fujEj62ETfKxY39bIQNXB8E7U5j
jWNb23Z6Hy0+J+IiiwBbDginPl5AgSImJUKQgiEsND6SyQc5UhqorAejqowkkZ22oypA56kBOoHs
gDBT5i5JJrJxyBck0Fvz9OvM981o0aE7DIcClz4tgBxr4rNFcLUzSUBE0h4AoSz6NacDti897iMm
um7oIVh9QFAwafRaVEigpzHmTdvRfC3e3u+9ScJFhljGM/nc9rJbtLoMc2knGnMdAeTENmb4+VU/
AIMPLYFYz9wfZHYIBInHzS/UORN9cVJb7nev38DtH+wCK7fq11lazW0kuM/hvLnMiIEjmwXAHVDB
MM7KY76MGRpDiw8peJilfjn6QqENxRZx9D0f5tGBGeKyUTHJSDA9rIHP3En5JE2gSN5j4bq32FH7
oNA+qCmK/XQzZ5Nr6nmK81cLagLSSW7eUfFHzRdKi/mbLT27q4hvxY43qxZYU+M/mTzkUvxKeh3c
P+6RtMYWn+VIONBcPNXrcz7tKdSvypt2GuS9xaMmaD53IPabSL7xQbpXyr2KVqOTW67OF1WTnsms
9QvGb6mffCC+Cl9Kei56j0xcvdyDMXN/5sdqJrdto7UDfOWeoVxxG7xQQqVXyuAEGAFWufQ/xLHG
r+ykLvjnpIZN8E1tEK9hnHq8SXnQEOiE0YOHtMSXVYYUiS0RM1Ax8pn1GHdFoJOMi+dY9sYXI9iX
+brdieleQWIrRIUhs4lAHDO7NhjKSfJxLoQCbF1czJn9CbpjMJ9KXZp+gWPwVSwYOJZuppEqKn81
bsUaOAg+2qRfW3QIdHgaXj6AqV4NHFTfvHTkPrp7H3rD8H6jidtn8GchQEoeBplvYUunwSvsngqk
qnrY/f4SYv2sT+yNkO/FTn3GEzgktupYWtqu7f1vZQefhWY+JL0aHSl5BcLCn/O09r2GOqEuXvGR
8MH93AFbF1BaV1sC4p1hwmmzieb6t6LrVV8wUSdjEJudsmquIFvD0QFQroJtguR/TkigmJK06kqQ
Bu2frskIzQh0MNA8q+XxsboR+JDCd0zpusOFM7YvOwzaTArYUps5FDFbcQ1BcfCb/SB2MYwHXUKz
oIJpvWC4e2DQoaFnCDhH79cr1afPXKAzAji+HRpao8WLu0QBZE7No9Y0wcmIm1F7ji0Q+bODCkdK
QLQfDNF6X66Zvsja4Et5oi7ndWXEi/OQk0wFCF0kypZYf+2F8gBCr3JwNcyLknq4jFTj2dkoNNyJ
0Syyx8zFqzp1Sz+W5TXEuttII+d9NYpRjkx2qdAbRyy7YXD/dHv2lHq+2NfLF7+/PhvFBiQIMwmX
Yl6+QEfwpI+sEB1yMp9cI7dFR6o87J3HOgD0P3/WaCujjP/uQL5Lae6/ODzDszSlccfAkCliZwA4
jn5qnZrCP1uiTM38JoqEsmMbSPWxYf/pfkHOIcCkQqSIQPw4rFjJB5pVYbKO1A7GiB4L5KUHl75o
qNx+5DDY7ehIH7ClMdXwwbpR1/TjA5ZoIbFQMjGJRe82mpAul++uZp7yjy9BxFXZxiXkpK7r4eYh
mj2GjovsqhLqO1yi+vQSUnrx/N7/qXFXmrbdnWMgsgT69fLPRQHK2zkvQu1/HJEv9lUGN7WfwuSI
aQ4Wcngj+R941iFOmvgF4lzYDFTHUj/5u0n3/0Wmbcp7lL9MCl0wDB9fnQJQ8YEkbIiRCGb3z5eS
PbSwLYoeZ7UANfCk01WHLSOeV0gWWL8oR/AOLekPPromqDzaoEYAYXfTeMfo45e9qTKYCdKDD0GU
lZDZPZxloIiASUgOYnW2CtRm2SjDXFrvgmpMljuMhlEiU/x5enLalJdh6magBjiDZN0qX6hciAhl
msVp5cIqy/fZfBYZHGAdAch42tbk8ITzikt1m/cfgKqcMHxqjDbMr7AHQ1VONrHG+uXD//ySVW+z
yxZy4BGHyNd6Bztaav/kujWerQ0BrR09tEbAcPi0BIdLT9iMPbt2Jxid6mbKvIQgtGd2eGIF4HER
+RNZS4udI8ySs9THdefDD00/H7qJsFv8gaIEMu3/gjI+uIQUS/sWTOhZ+ZSQC89iffxfSdbZSOXx
ld8G36ATAHxzoSF0ic1g8gZ2H9+3eO2jElaMeQWZz93bXXns4B+0R5Mb7k4EYjqcD/A6Sds7t/mz
uBLVvwqmm9KCpKNhtdGrtZZgayYWkEq2JgavlhieFgqI93Wi8Crb5ytxL/JxOeN78kYzOpEM79o9
gBogwSq1Vvl6Y5X8eeH64C8XQHoXilwRXNbF6uZ43gtiR3Lkzw6I3Jk4NmDJ5TjkvZjMhcwfM9Y0
YgRjwz/8N8XQfamxDlk6e+32Cj4aHyqjkJniphMkPcnencZ+9WAqiLKosxI6MAi3XQ29xlVAqXZK
iNiMR84ubfg8qxx1pOrawSqpyOOT640N7jJ9HQXZbevrOZ50g4xiU7h9TgZW/9K3h2FHU+cL6QIx
EoEcfHbqh4YaxY9E7hougfB7DcevOZbeOtJUTzj8DRp2PdteTbXGCglUYmk7io3QbvJHcQ8ebQXY
ycwvSuF5Au7BxLVcEUYMpbBWHIeMPZVrDNI6/i40rXqVONSPhk05nm+qCadntBCP1OPTB6bCHb1v
ztoOiJaNN4cbTD/CeXagfxo73voGM6yTYgd7jkOqH2yVW7D7o/wPK3v9K3WNBjcFcp6097XuRuP+
U6DfeSZ87YXWyKW7a5MXeGNHWdeWZJ9y8wiWTKhghiUpOqbZstpe49mDKSntzJdHjWkA2fcxkmoT
2TEoWnMnZfqPCUtT13ueLGuldqIYcDzJTSBL+knLiMaJYMJlYPOWDDpfGSaT7ijKn3u5w8IUJ0Th
pYpWjAnYruX3s8ppB++kyL2CooMJhysq7EVrwnYb0G3x0GKlMrjb9FW97RMG2hKARdYU/hUSCQGG
6dIYMm/iOeQB5lYxswv9jLLpftUI3t+ljyA6glwGApFJ/t62VL79/9/KIfX33axeGY2L2gamUic9
9+ZO/RxDTkwiVIXqSrv+mxhT81mfsQJJQGREfPogaj1M+E+8KIWv5Dp3MmqQ079ps7jFCovOvYZ7
oA65C8Bx8yRLFwo1zpMVp/AkxpKhMrn5TT9FcO5l7Q+7DmuEuAfu+fWV4bU3VfcfoBJ+cSjXsjgz
wNopsby4bkZd9xrEIkjXBuiimGor/Y/TRdC7M6DeYitPvVkqsoWCEX8BNzuI2BE6KEOTAkFGT/by
16/2ZNwLIFGdPHGEe9tdkw8Nns/r1go9P0HvygFrQn70wv9DVU2e7JmXMj/ByK6rQOyxU49Ws2B3
KR9Br7qbZ3X9Y+Oq8ttppYCQJuFNqL9nO1AekITFUMQ2zmsMDv+ZHZgAtGUrnQvdIr4/vZgsaYXo
U09AtEwi1mZaevs7RSbKtSJxria2dSAqSepRSFZ6/h3LVq2mYkfHglVQ50NGpDmXPJneaY9GkAv7
iYZn3wgY9t9vk/0I7s6085KjbQTdjghKExzWGgs9ClJJCHIH8mcXThZYNt4KuNDqQ7QFitXU0p5e
RGNraNThcFOl5FPDJCs4cTSp7kyrhGF5dQOajnH7YXRPOFlnb0uNNzOjR7vtDoqLV9zm79ozOpN6
eR5XQB1nmoHW3ZcZm2KrOzFF12kbs84AqvhmmqOpgsJnBemf4sVMw94mhR95tV3E1po9AVhJiiIm
oMqaAprzkNlxHUmTMaEUrGFvJdkDJOs24yjQGGLZOYERlNfuCdOMpZNFktYjEW2v5sUcpHq9Y5Xo
aSWyZDo3YAFI3ekGkXt3oDowo0bAczZ6Am+bd69ajPcmlD7MHmJR2RKZUL1vQ8xq07PaHB2oUdgu
3PnH9EuKK3IEQGV2wZktBEL6CRZ9e+xaCFOkcZkzxSFaGXDi5K/jACfcytMoDxXFjZuIwbw4dldN
8DxnHLNnBviuZMqFZa50v3zMqLatsGrow+FI2vdIjkcKSL/YG2vtXtOCbxKaoeu7Uh15xWg4UDBQ
Z7HwzfCx5f+pTT1TfmAAMSAK2rqsH1VcRpX02u6xH9JgWaDrSbwmKdeiW/cweGEjnXt1QvjLLrie
IudZdaa7Keb+EWRYhfDno00Fc8X6GVFQCYTRlI3hrHvHv73Hh4bOu/iK0t+Li4EUKLgqYSnzikwT
MWNoD/5S/1soKVjaYbGTl0Y+ETpToilLnSkskbE1hYiLFxJX8gyR14KsgEtQfJ+IgVpbyZDrOaaa
irNZ5Gb9w78KTVc6BaTr6OK8tZJI8esKyGiTjBBXjDAquCC7oLhvGIloEK7e6CY6ojoDMrhTswPb
LxsTzMJAQEdbvavFfFLAK9/4CGErp2yTq2ALYcr41TvvkqbIA1IcoiCDGk7DdAmh3/OqqRMWI/O9
w3hnLKquehz4I7Lmamw/sD30qeIwSDqOb324hNbcNTrgYls15ZEhOFDXi2MXlcf5PbU0m+qau/QI
uVjFHsvAsxFFBcRMJVJygjnj9GFlKD0uN1jvHLh+FxcNLlOrtYRVxM3oVt+DmLw3SG+1vEDRCDZ4
/VnDBHK41unWIptM1cyBSdeBEiFkBL3aZmQDsS0/abeNXG5sLYciTVEcYynKn7DLSeE6PjX3kMOb
bNOlzisrkmdsI5YItorqZwTXmf4eS9iu96rPVvO/hGApCfeGao5Erz1F1iZBJnxRJ1R3n+l8kMHW
8hi+xXHqGCabMUwO5tj06I8U6lMrz7oCIG3w7+EXOuPNv6tN7o0VwdsAZGLcLoCYE33mKpR1LdXj
7lkf30KtpAiCXhyC/SC4gqFwxmAUUWSBbKFzHzsQfdoNVhhYq/alaclrQMza726Ml2Rr6SZ9u/ls
ipv2Ic/zc9q2m9q/HqcvKONDKoRD1OxMtncGLsR7t5bqGkUOrTcl3O1Mmglcfl3bzF8KStL8ZuCB
oU/JVyElh8C1IiO5XVsmsRJLgOqq4VFxsKCsJVXWfAJDMiZtiTCeBs6WmQLEnjV3+NrrrrAN+Ugl
NS/kfxay7s4xYFKJNcb1mvH6q+S62MVUBbCujHQzICGkJ/Hvi7F/O2y35ic5sqh1xHgeO1I7yhGG
DPnw87Rn1aDrFBjbNfnQ1AcIWrpkyUZWsAGLJ0fOApw8mGmzivEPOa5+2n2hOeMejlPuamuYk9/S
Ba9HwreX0+uwB4rXMn4KqhIKR7MuStArv0S7Xd50iNZJl1/BZjADskoSk5Btd9qlN98oF0JYKFgv
yfJU+0oWepIjVCDPhHWptpwHeCKFZzKzeFWezRYhbjlf79paCpTR5zjlwZrwIiyHa7KK/mLB2kVt
rLjU6p40x1gIMaPY2W5dXGGz25e4/C4V3+y5bNp0QDvRNsC+f+KU9cgkReR12YQUH1RydSIowKwJ
szGQvtEFM6dXzrMvQMxFV+ozRk90GdVWPQyGJBZuQj9irEz1DZ4Sf+KHj9WHQC/1t0eiA6J9MVJe
gQjzCYWU5cGNh2XVmvBq339Ca5bm/qYTzpDZUiSr8W1NrQY5OzNLbeMJ5lmMnK+5u0PO73KbYdkR
Y0b4zhOyT/bXbQWcRKoW5whJRq6Ap3MYZ22a/btQiNPGU8zotl9dGZFRcQkSTI82aMVYT2CTLngH
+A6+wjZ7f3wYi6ZxpBP1BJowtcewaGF7yXa//LtcauRijKsRuRn5YGqcu/4ptAFxq6iINEeksS5/
x0Rtci1+zPFEUqPIOfavrIJLI3UU5rn0lrz7frMIbRzvsCIspvp2Oj+c7PrGj22+hlXU+oypqkhJ
GXu52a9mNsClp/MxIbCA7LKEg+OovdP//mQ+nc+/Q9r2RVRXsU4afkKgLuhohGBU6ovhDgfiXq9y
TBb6mf8nnYLeTuqcJvjSg31waY6dmclEbM8qSS+1riZdj94MqB/pnhwde23wXtEXAiCn6uh2s4EL
1sfK/Ux6avlNC8vc7x5zASgRjjgsi7xc5zVXh5yXhv5d9E8MdsHK+9HraLDWPKNLV/qnS0BY+UZ7
xcAPZCXn4cvqlQ4ivbKVteWTOF9nioKrochXxaXoP0BdFl+ftteRf+lnwNyWTEseDr9ALuactIR8
N9oL3169QHo5gty8NDTpZVFcE/7uU4KaI8ZIp9trpb7+A2OQm+BpZ3WFIPBiUhcbSLA9ncaFs/U2
b0Q9WA6MwCJ2i0WygM3GuKP/0p1ObmZ4LxxhHP9H/r9evB0ciJcocUNJaJLLHPcRdlU9rVMjavg8
I5jbACa06RxRpoDdHuw4GG0XaBHgbUOtLB6UjsOcQtNijTyIU3cWGK1Z+2gssLvOXN7zKAIMiXO6
HXbUO2SqdTklRTs/0GAnIr4SUPdZ1mWMBfgEe/ATbFC056+jiDCwCeq6a8vAdtsCnqdOBrgpR153
oXBZGcr5cojz1cJZaBTKMbwh97EZffIhH4R8MSdQG0zo1xQUgiEMXoZYY3uGnvOne0H+7Y6y481x
tPpCzBvhrkhFJPCv8ddgCMOEWaT/DsJPyiqj1vvMWYnJWE8Q4JuFNb7xiLoqDPHaGEh/rJ7uJhFn
gLhYV/X55CYofyWjQ/11zpsXKFCirN09ZY67J4PbsYOA31SzXGiyT86cfmDJzrydXSRgagZHgsy7
Kqh9CZaLvIEcjA7BBEwOUEBm4HP8eWHhUrnOY71qxwrLGhOwAzYxVHzyc7FHvzkXXdI4Sb+WyOrD
Ot3w6KwzVC4GOATWBPo0eiDuTP2KnPD4TuKDZKZBDb/+fAFJO93PbnuLOrhyAOH4ywtYOiW6YXuw
U/13raUmrXsQJ9n6T677AO2RtTYzkJZiIirE8MPkBEKWlj7TkgxsHFCRn0ALrVFkqlnkx9fGU0z1
BRXPRCqGNdhkG8hGslE0POw38sSkRZfwm75BEgFkooIDA5M18d6SRcan8RSEs9d0BWkVbtE1Nly9
4NDd7uXfRfuzA4KpW3u1f4HO+VwinUyPi1oalQMVqDnl2olPizp0XmNvzAt7BCkysP8087J2cHxx
u0Gcjbhvkos+sBxR/8tMnHJM1r1RVr7ZCTnueGJunknYGId94y1kDrzpN4Th8ogEry6sEqWaU+oK
jLXJ/wzx0r1sEnv2MMOXtdERCTTKycN/4FnT+RaG6VItO5HPxUghQpKTmWNFIahSFJx9r6gRZhJa
L3hcEKtUn60ar6t6iwX+LvkUDbmS/DnwIbGM/sclSLwrjoTGGDzh415i06MtUo1glCJnmngfPPD/
m9VVSfFzEURvbk952xJMI6ftec44hP8OPg1VP3FDclU8quqpaOhlMRl7jtlyD5SHNHJ+OulnbqhE
1q3udbIGAPzgWhUQkNZBhg4P8X+aMBP5gM6QfuWpRtaxui23kKF2rApgNe5+DvU/h4WunAvPwhzY
hLzE+M0+Wkw1wmzjm9UElHKhsn0zUkqRNcILD6xW/KsK1G6ubBZReB5XPssOBOA2YDFdWGXIjLdG
07tZUvN0odaPhqZ69J8ddNcjGiISMu4cZCWOtXxT/qqKTDcWE8BiTghcZYpqqrxzc+gQ3nXEZf3z
qlQNzlDOcUyqMoX5I/7539Dc5KL09J9RxZs/cm3g4yCUqFbiV53eaHl7+79N/RE6UN0iaYLfYfSo
xObaCjMFlg9cFCk7iCb8+dLydfeZNrfPPaveQseXriiznXHjqWCp9tUprB5RL46mJWt3zImnIqre
kt3apLA2F8kwV2vsSIKZY09r9pcLrWDiFFScOar1YS+WK16WSI3HeYCfySw6bP0I7ffoLqzqvrXa
eg3WZDqPdHw8B4T2z3ljcymymgAjmvMhLUXCuMXv6/lKw67eCpLVzZIv1HA7rERw9u/ZbU0Nwr38
lixtp9svGTjvVFfAJ5InxijWBDsesVFxwog0JVC0csKpogx7i2tv92bf031QXB0pdqgDWwCReyXk
+0Pkyi0HX+vnu2DULACCFxt/pNJERhuC6e5x97VVptY+aXyk/GtxM2u8n2B7lFO6AkAW7Dh7GKxE
Wc3EylJ9Je6cVfLeYSD8GVycNQ0aFXuRJ2l4LFUZitInWiSO5ghbJtPjeCRxX5v95w7dcjkL980L
A/l6+XUAlNx4SL37MZsb4cv/gjkEIbuppqCwIB+1dLh5ZN9nPPn8kc5gARHtKWyXdFXnSup9mU5b
K0DRDb4EnaJzq445ERy6J32xCw9En421FsRaevxqfxta0bHXFqdpKAwK6MaxRwdCgMUKCkXuBHUR
Ie5GxOsUzifqpnEsSZbjYSWf/Fa+B03Abcji2dcsa+A9KSR9uz1ir5NzraGeBhO8s8SkQ83EHzbl
2/n8MqlGxYhqygH9THZyjkZB6bj7JawsAbmUhbKzyfIVD4cuOiZ9Tw5inIYQMDK7XtgkOpb/K7WQ
WGuZwZQAv4kP5Ye6HAcpA0j5BNfZ8//Dc5Iu9wlPbGlGU1u3q475MvvhP4cePL1eEPVW2QCHembe
+/xhGXaJXnhyi1N85DrPRpiIHyDYvgI6ZGhRuK1zdBItk4EWjSdGw63lkATQYqNz+wPgZVWcuR8C
FwQ7QSoMAoKzMtYLmObfvApOPfxn7MjtSGF0j1JaQBHcIzFocw3klumzVxo3C7/5So37vT2JmaUY
zdukWRCjGIHUUnTlj6aaB7zofyZwxpLTowct6PptU9yiaGE2/70VCq4bKP9f72P4Z4DeYzTP9lR6
RFJJ0jEsofP5r3misl07AycWXYPF+YpBky3vY0v6IiNmVoeblR3GTH8sLL/Lz1gjT/er00pDe7DX
5uaDlaGvoSt5WDt+7hWgetHa/pSRyegb8GS8mdoBoWZXF5q3iH3cYar25WgUQrOqLTNG9J/u7FfG
bgPeg0afNpyTONlB4r/9fEnaOvRG5VST5iJbmMCNR27Np8l2+aK+KXGMfOKNnEGsZ8GuG/AtFKKx
p4vNWMu77klCy2w1MGt6tifOHX7Ockvwf7AjhJQ4sSAOuwQWWwtG8HUQG5ikVVZf5hTnsLP9Izzm
M+RsRUhumK84ZFaN8G3OX4En2Or/KcZrPi/SngMsMKhLeCeGMdT3w40Mb5wNAUjD9qRD+42VRO0o
W/r2LqeOcVa8QPSD3UYucQ+CoVmWs7xz0daXxNn7O2G1c8eZ8pLMFCR4ErPBVQLSm4qBRdiD73TY
IQeL0dhNcgf9uCAS32i6NFOHT+v7sbCkI1/bhfk7l7QO5ooL5I/eS2s9MyC5q2cSd3oZHZ6gbc/7
QBU9Yw+5K8aPqQE6g/AoNPDUmC2nROF1HMols1PGly8rwLQri+56pXm4ypzVXAii3exebmtdplCc
oRNCkb/Wt/yK5KlaVuWDYrI9xwEcRL+Q8EQ8XcrosjM6pchGaanh88kDE/fOvbtlV9SSFCE8hXdt
WAx5uznUDBdqNv/H1+7NYaQiLtv7Z6ylAObJUEr5sKlfw59mZ9+oXkGf6zFT7za7aC48NyItPRE5
9M7jWj6JPVHZD2I+lPQRbKALOv6tQlG+sn3LTgn6dZg/UdPxHlIY4wL65/h+7ajhaiP/Kl+DtKru
FZW8lYuqpVllw9TIW5Fd3ifCW2O6zDYC0hEIAbM68sScTgR6YrBh53aXjiAoDX6FIQa6eEYTvqih
69jh4HzurXMq7lbw5p48d2tzxuBcSKyPjzpqBLxIh1ClTWgAyyOo1+Avy7r8iaJAKIIqhK7RsLE5
4KPz+pnXBSrvi9rtu8XyT/5HupJfqESEcD8RvV4thMMN3sRxSIzqEhP9oU2fr9xERKruvx2dnlzt
8Ok5+g43LLsiy6Rs3aePoSIWW9E/CdmaQ5GnaQIqxvHi8lB/O9/c+NMAfACQ5+W55hBNNjRma+lD
oNSKhKHGiSeAecj78NaBZKpxjwC1ejxgiF+ziiEayXuK09e0PIQXVUAYUZtmCo4T4BaCYKQM5jkq
kdE+nFjI1k4nXRcZwzbIMMO3rZcQQ8lKJPwh7qrUzeq+5+LuyQGV7fuL6ho49r55U18Sz6bw1qGA
ZqZvf+CIIsOR3xZkaIBJ367eIGQlFAvxulv5d+gsn1HU13Cm/9rRzaedlkirVOjNiGm93pt4Qpn3
7uQfEsDUi0ke5ufsmQzg97LAju3OAxxvAnX5KnnY8IX2/PjWlWBlvaUBdFkFGhsd9ADw5odE6U1S
gj3Ha5WuNWTTfxsCvCw+MMVRjsuz060IaSP9Mod3pogFdSwQ6g7HCQCFqXLC11wt7bhbDRf+3ixD
jGi+cjfBli4FTKFLMLKmTTLietAklv6bKNxzviFL3Gbkof/Tu81NZDsnZu0i1CWL+JEaPSD0HJrv
H1pLKSlropGsSP8r0J0cqPKaKXlVMnBtLNHs/tudnD8wrzupt/IAkGwwWAQFGwpyyI79OQ984iMS
gHrJ/J9fLbNE/O4FA66p0pHiLiiDvlROf3sBfBOqSmeboYkeHTU+MxCy40LlKKlidRGTaowJgbLl
w0N52lcLKzY8LFPj/iOFpzL7x6w/ELVFKu89dQnhCJmEMsYfySsJTxRuycVhdgrWPEml1M6Zf8rq
/2FKo2kCgnhdhH3HD/vAEq3cV3RhUerw4MeUZF0PukBb7G5Mnq09H2XqohIsmarUYu4G3DKWymw1
EqvALa4AK0WwrG3j1w3IMe/B2c77jnva5UvuyadB/RIYdImAzSLwrMFm7lKXjwtt+OVL1gVf7Tdb
D5xxb1qC46+xEP5g5F/H8Tibk3v4KwQw7HqtzbdK+r5SdlbtAQLHbEWmPw5xshcJAkj0pm6pRgBB
41Dg6zq7gEYd017vzXAvP6hfsxzROo3/l5V9EGCJr9OO0lFPC2B0tp0/undDE7OmQOz2X3Itdq9H
3RyBnGVk59fesqNFstQS2UfyRWfpfs9TAtowsDI2wgdxUpCVN77kIPd2HIZdZBJ4G4sIfgG9UUGm
QyYsso3EbUZeaWR0f6f0iMIjLKEf7sUuQ7H9Ru1pHKMptOtU5CKcGCMWzbt5tKUbrUH4lz/0uXxs
MVuGrNqP5WlIcufGT1gHUlsRWnE0W43aw373XNbxpOPcmovgMmj6U8+kYO3uTvtKT2kOdooGkHSL
ne7G/V+QmCSR6+4HD+irQ5drUzkol4YSSXbWtDd4OSXhp2JnQk78YRCxwXK8pJofINtA3grs+Io+
Cty6SXIKU7n6wJ2Ljgw+ZDE4z0jgVdss/pVVeisHOLP2MDXMmqfW6FN4vxP84PwbzeCXn1wvm2TB
p+rRYha/jOM7LPrB7gO0l4hZN9dlqt28v/YPXdwbjHD+lbb1psCFVebxtYTbUn/9/NZA3tvGNE5+
QRtPXtTbA8WWBe/qY3F0YYEjpK8og4OICphWru8PEw2SAKlw5k0aCoA0/ShmR6tjkZLuEz+g9Pel
loz7uIIzi2K80BC9PFC0VcqU9KkqB4Q8nUMEZqoYSi5bnGNvDBXKn6pr5rhoACks6CwSLJNGbgXe
VOeFR5QzqlT65I2d8bfD3y0xHToPBgb8kdZV33QlynxzvhdmZO5+h229e9t7mLSiO90qiaiqQ+fz
2DWTYAU5on38nX8v/fcPYz7Z1pi+grV9ljpU61qR+j6IRPhJV0PPkHCoLOxLc3qRBPXwr0LCiZqB
UkCmmQg0lkBcq1UsjP3cye1Ue2Pj+tHepiuck2kmUyiVKDIpskVZ1WdiXFIs6TxEvDRBI2zkZmGp
Y8dH+eXxoI/UjvtT0QTqa0lNjA9HTvYjTgo4t7cOU8oKvIzAd/JwosB8V71LAE+NxLV0G1tmCYWT
OET12MlXey4soitqiv2VbbngK9WiVcot6NQ903o6kRpvOV0VF6BpIFZSsMqMViypk87SA+p0NKPe
zpoOpG7J522AwTxYRwgAwtEk2eHaNOCqw1DTUJiVt9SnfZGYyBKPN8C5YshhxA9JTz7fo8QG+8F5
pStdU6T6IFHyTnT8nd1WfuiS2GblslHWfjRGfBanMqP8+jvXzTribdG6YwKnKf/iLA8TJhIKyhab
dPEGgQRwcOSY4564h/qCgug8KHKce728NlcinGxFISO6dpNvCzvnHvKhSkPf5+49KsUbpHxg9Jsy
QyFVvXO2KcGUXVISn8dKocyGDSE0tTckNJo+2/Morf/wemGVmDEPMpjrp1hJ6oXaew1mEox2eZ8T
qOboQozAUN6hMPUuIwPG0t5imnqJ58dRmBxgED1lrd6GQLBxL+bDt21spSs6jN0lDQwRQaleq/z8
6GPyxljVfs0J31wRFpfxdpZPYkn47UsNWM/uLrlZk0E7AG5IJGakHfv0Yrm2Zozp8+pYv93FbzJI
AlD38KK/F2h/SNbI7kcuHTFjFfSuZXQk56HL8WVfgkPq4KhkbFtk1dOoSocK5qb/vKIYYqV2heYT
vXAkaYWUGie6rpa1vItncpJzxuPUhNO2HnU6cA7EhOxGYUvQdiR0EPymh6lSw26Hi+5AejzCOM6q
2fsRPhTPKM58dVRlg0Fn19v8nBuoX5X+fnLH/xoQlF5AoQYnTmkobEaPf2nM9GO40sNtoEnLPWB7
KonbTYq9AC1pzFGpltl53FOZSXl41opO/4NqSUYn+ELdt3G6aFk3T+FaY+Au0WdOwEvfBnpNFLEo
YLAczdLC4wZSaU79io/fUFhJBUEB+p52/dtux6COFS+kqZTKAbEek9OGWb1jq1firqSyhh0ztBbm
ea20/6RrW9GLbQdDWYdXyJYZjRaWaJEpq6FubVJ6t/hGVQNZwaLuORYt8gALmoMyIee9ipYI5ZOU
sUZJlHpBzMvLndUqiKm9dkGyjyk79IvAHpiu8VQ8Zx1DBt3yW4zjY82PWESg1uojndCKgq+SJ11m
LUZZRVlL5OeoeSGTGaoMJQ6admiIhDsINh/ttlrJ3tQayYOn3TdK6f4FeICO9NmHr6y81VDyd7Mc
INAku5q/G8cFqOIgnjUy7GNRP3w6jaWfutsZcXjeWZP783lU/7OWzMoUJhVsMbyUSfwbkrl2SfeS
Uv8VjDl5EBKe4gYXvjKilwVOyBLF/0G7plr79sM0+22QOToHVm6A8KJWneU4LaREYuRHz4LsOnci
1qhDAnGMlpzOUSxAD6jMSfRRbXwFZitQmmgoetpR2QV/L2PTp9RGJ1BbCmdHEbttyv8jQiqbnPfQ
oI6pTEk3gJvPAwBvwmUFUJ2SfIOo20NCroYDBjzG6+XG9nkt7VrVEYn1gNqvyaerInF7yfXrSYLV
8KcQi8E6SlKzgTnKNKHCeFQ+fYpkCdKf5P3YJ9p3tTCX37elpe0hmfsNvPO6RJyi/N8MwAB/Kdrs
dmMhR4vS0uu6ETLmw9B0TqYYk3Y9iTkYkh5IStAdi4MdX5VCDR52FVUjx1FyS6uQ06PDv/SruNgM
EC/A5gy6o92xfNafO8ZiDNoHgG9ks3yNAlTH14MxD3GEj9Hn+tDVNuPr07zTXaM54GFKqLVuyDrx
dijSeFBSySnz6IdRw/nLIM+dI521R+49Ga1oCSphTxxMOGoOrYSJPrExTiZHixEDfLSCmWG8L2iy
fRarRAzDfutWVsqII4XCge/DgsXMAkMd0j/g5Hj04Xt6oBFvyHHrKo2ipo84ud9zu58Ucu+/OYy3
Pch3AXL5QjtBhiB9XfuUTE0I1jXXjogIrzCECEG94negojElO6pbgz5tttAkME0+Mbw9/He3Nk4H
HJW3YtYcBUG5IAG+Lk2/LwXiHX7uZxbVfpxjmNn9eSc1BUny+dysHz3Ook6eibDmYqtZfqUsO5hh
DT5jRkR1lbzQd6H/66za/IK0HKQR6hQ6pGtE8i128LK2ZOJELUVdUZX8iaseVAF8SxvqIt5ETS/a
wsmxXVQfxZEADoePFcaWbDNtpcIIHAgl5rhJZPQX1ycCSxqYVkqBe1rHQFDiTylb7wIgpuNhPpx7
kZ4dPFYiAyrZQSQdUTbhRUpbkfQBh9EunaXJpjrCh2pu7SBeNVCcu4csIlG+1Fx2EOh1F7LS/rqr
RNJ45gBr6RU2DZXwGKfsiq/DoPQK+wOw7IIqdua3X89oAsIbYbcS074AtEF7vEebPMeIjuD9crmU
7Jd3rUgTuv+/X+4kOIqDR2k6S/L5cYfnJRrTdJzS0kUXXxcQfSYLFG1LZX6IYslY0liUyR5SDtQS
CZiFuoSg6H8sZFTDLC/L9/UxLgePbcIJEqNr2puuH1B3w35yddcvykBJTTmX74s9UOFONYLKaoNW
V9cYWITQ7oDKfGD9yzcFY/9RUuNEVvMu5QsUoROXZEr3MHCsTgDong9uyaA2LYpE6EN8CZRSTQjh
NX2nZ1i4ypD2HKZF4YD5SaoS6FQi5soXF8pGHpeO4b8c+Qzp7jGS8BLICEjCncy8bALYbcfjNqsA
cplOUct068Gmi3ZemK20ak5g99WZMTfVezITxbfkuhOubDcHYaVARgLkB1jX35cTyhqIiU0SkPJq
isT/dFvM21VJ1SVg2WlGeH4sUHzA49ivvZxFGCBfEdl5oCTHwrYWAExZH0cyoa+kj545ocSQDtza
Thams28FBDcwhBABiB8kKccCsBLX9Esi84Ee/MoY2inGtyLjz2vqR31doJ2k5Dsl5Tv5OGHkqSiP
OxKQEQ0GmBOM8m9iLGMNSh0wdS9TgdDke7K+srgbZYtXIzX2Ykk0J0Hw5JPnEM6b2vkALLOo9WdM
3TTZUn+BQXoxfpMQqGw2AlGOzEyPRRilkFzp+D5vZcMKapouDD4pyWoYQGH9iNeqMPnBY37qnj7b
eFfqYeSeGs+6UoE6+PVFF1xemDif9Mg0KRalYRU5NsZZtGRcO2xT29Oh7cR51RpOaLKkLjDfCXGj
iZ70J7EW45YWN8SVY1mHxpV57Dzx263dyTjg+yuSkM+D87yLrGmnJGQRxvivvWIYm/oyYBL+jume
+5QpOR675hP5cOq2xoJD2l0OFsDL3KSJJeTpnWI4SN/wD5npl68R4UF85DzLvZeTWNEx2x5N4OHl
3mnUG7K4AduXA5rqRf9geJTcztbIyb8N+6EfofBhAz2UJyujfQrKksudeV5ynykD+tFzyCXpJDsI
IyVmRPLt1Hup9jIXXJF3PR/XNAYL8Ul3h/LdCj8i72+lPyRB/3zzcOWZVL5bQiV5e5lEBcZ/3wqx
foEfDEueUw7iBMaobweo4ZZOd9Qhjb7VkWaxUbGSuEUrFKRVYQefrZpwM8F/5P9J39j6FxeqfMAw
YR0XIC0QQvUvDYgVQO1SZmyKH8AfMLiXcinKJ+QAVxGE2QtX05PAWcgCuYOYjZTMEEeEpOJrxW6v
9QpQGFuz4qlkc9XwBPTOc4BPDZJ2MfBRjgVsVxe7T1DmplfnoyDL4gcpkVwO1OBwgxtKedDog8s3
FVnBrslsPoTQm1XiBTpwM631YvPm+j/WUGYgJi5V8nnHjED8pJ+aieiB/lTtauAdN1Tg8SNkA339
I9n2rPApMIpOuuSy/zJyiPMtFH2argyUbdRmrxusdFIIAmFfScuFv9+y9CfI5DbzoTm3IYXQFKNj
B7ArWfi9p7VKlau6oT9VkDLbxkbBmPQJ+2/sW++nJC6uRH10h3iKqDRNEac5+T51ml9n0qt33B46
fFtkzNdvA72jC+pYS/zwGL+4VV5uursFwEp7Kagi67BKKuar1HRCFUYVda9pwKWvUO/onxbSHjw+
55pClMjq5e6f1yTBPUOGCdI50LaaWRuLstypmSg1T6om1qq3UUG8jal7bLg8pcDM2i3XT4UTG9HL
HR02vLm7tMIduzNw+8P7NKI9haF3+u+8rjWRdBIUjUd5B5f1h15soxtQ7cxUAXlpZaDPteic1cAS
LgQqI0Gx6vp4kQLPOGTWo6keSTDQ/OT/FtxdSnN2/2cwcpfHk3YP8s1F8kQCYO/0MFzihDSwizYI
hGi8TOq9E+nJoFQUHEL62d44818c6H3/3zb89H6L26xuEtkKwP2MqgiLMHo+jTLUy/EJo1zRGih/
VwEkTaOP/qPuTrF0H+F7AEwVOMET/ROJPlC57vwOhHPJvQu5N7FsLMzhjo7S0VvBvjlmeKA0Jp5S
sNoiQyNTr1sq+8FCewOQwzuY02rYD7aZ3QBgXcHUc14pDI6JMHIy/bc7+MtU/AMw97A1ZC+xVShr
o63Cnw9utKiDxvYa0DB6uPTCcygYVvpgN2ph7JuN81IDc+iKPJ88pz7fyS+takyk10mFVkvfOxmP
2fHnMGSMDkO+Ed+ZlLHVlGjqDcX8Ip9UKI2a1MxDg6dMuhtO5tY15jWfmEBmQ1A+jsL0SybliS9g
IPajqdGJZMn9jlPJm1TofOBUyBU9wvPbgayn8OAD7YsBtbOzwWC5x6VMQtG01qQJT5SfZSZWcBS2
ZnPMOEe1yfy5Y04w+4Toqqv/OnMxUVq+mOylel5R/mTHZtZBaGgU26syMhEJzWee3agmEUqJlu/g
gZltZSqJQlRzj4HN5G1u/FBo0SMkTDbVYuNPVG0HuArN36nCQ40FMkWtAGJa1uBRtpsP1d6wQjJQ
xdqMXhIoNBA48gRhSX/S4E/OhqP8+FHT/RB+bcsgJTJ8KiMvkyiXnW8CoM2mTxjpA0oHLUEXIEGl
x7jmNtKB1EkUy0KrCnQIlw/5r3t2A4xzkjFfdiLYMrM2U6mRdJiiwBVmB6NFBTNVcwCs6UYRNUcY
nWKvXE4bcVmVEPoV5PkfQbxF3+XsT1w+2nmMkXBZ1/jIZEhfnz1uL9E/AkiZY9D1vkLMm9Jv4Z0S
uSbpBiiy736W2YwyLZUXaJiy345lHrOCw5MFAXimf822WgX9HRRtKw5UDY5bFR582n8ME8GppOEb
0E2bON9shcJMZ/41RiiXR0g5XmR8CZDarAsTNIBO7Zt0u2Dal+XAyEIHvn8EdBEYPgAKmrZ9qtIW
bWq1CJOtkbZvQhIIxctC+BPVt2ONSGXJbgzhu792HU4yMSNXFKRlrujt5wTtYBUZyE4iGXgal523
yBRxnIx1S9qeFhd+kqoPRSV3iyxtdKTAcOqBPebq9Dmad/cOMVyr9TH2wyYlADChRUu4jaaDebW/
L6GmwnI/XYowHUNi0ZoD9LxuZMUjY7aEmUX5SYrzcCrYvXVak6QhsTvXBl+YkkP5bm23rDTtfarT
nPLjpjmc5iLQTckUXt2cXRkaX4RdHP9+xlJm0psi7eqRO1gMeKFBPEmutcZ5lhSn9e/clBqXtgUo
cdGUdMDRfxlbOv7BvJH+Qva56TbsLNhVCgKuscOMhi8i3sFyK04CnqXYVCH4iDEHQ/aaJfdvvo+l
D8SSlDtn0IUBe4LLVnfuuzIZzW9lvVdnjkAELef0kL6xwTHEraErRSZfyfEKDWXiEKmEsIfP9OT0
hsoXciwJFpLw51e5TlZh0btK2MmPZBXh/sOfNiOOM/jy9p8LoAwMWx9MUqDCKIDlhvjyXvQSj09a
zhHtexHVVrCx8cXRCbj6MTalGykTY75u8JIDoz9bGS9nXTglWYwSck2MaJB6AL7GFkoHL50bFqbi
OwalXRY4LOblTz8xDg0ZeG9Q5QtKCzb44+LCIk+9CGudFNL49jcPyY6UYKKi/xWw6YHt6xt/CfsB
e6E44bnj02qfbPdAuzctJ4zBDlItghwzuu9HfKNbDHLgR8NnSu1bRhvTZqyK7cgYxWJ8i3F2kU2O
CZZp0ehODky2IaxffN5jsk5ftGhAiyCg6RcAO0Kpfen/5X3htLCUQNHwuDzi9YO8gCmVxmevGRRD
6bBuygzqFhT2d3kI+Vh5pu1Uz/FRS3FuuE3qd4PK8zXA7g1OUrMmRPY4h37UxXX2NhG+tXsWDiBH
LwPPO9jynsbDunkt7ESjiOM4ng9WnOnPmO3J4td7ldzAK+kHHWE8Arj/iGWp9/0vnJ6bDJvJ78+m
SPe+w7cQEk4hpZIQmIMfCiN6AorNVqU5pPLzUYaSlJvWMmHb8fwtXCWv4Xu8+UCVCgPTw13IAg+u
UCBcNQrzul/55MPHYdu/rV/Xf25nlg/G7T6YRg2wWArNErkh6mIsVmuXQo1w/GuQkPs4EsLOZFR1
q/q6lFxTNVjd4+OHHteCECSfOlmkPr1YAgYXKEBjXEGTPHH2Mm2TPItOYSqkraFat/ebixKr/IAl
XpPm3Rr8+QbyNZSS/RlBINlQTVqxymAkEkWw6hjS0BMIopSNJZtOcJry/WEsKfyXV5v9j2JUkfkI
a9pmBw41X2orfx3JMGCq3VTMtXTkd4QkCnxFoC73MIKvPJlTqUqR0TNYSzaHKHE5XVrM8B/SXXm4
UoJF9s+c5Hni9SCZ+FEnQ2cd89XZadFmKWp4mLrxS91HtK/UjGxaMw3pPQlRWqMRrmeWMPEAz9mM
OJ7+CqjHIqKREkvb+tCMdXZnFE9cBmyT2ZbEAE76Sjzg+yInhCIbyril+ZPJPyzoh1QTvEN7zyoE
n78MZ8oIDwLh4j58oehkEUQM9lB/MJqVA8F41qBIgTlbMxAu/36drwLyQJfgaDR/wQk6GQWNoVAC
aEGEQH1OrWF+VyYzOBqBwGSIDuJjr9DZR1n1MR5XXrpPXiWnizhp9q5GeFJitB7/KCfCsBwGoD6Q
j1P4NfO2lYUyJVAiEfMfr6r+sdnF06llAmN5AKas6I5t8+86ZE2FRKe7c84tf7BunKvsvbNxrwmm
BO0gYZWI+efyo06GC/UHZflbbGnnqQLrPgl5skJtkqEg4Vh5YOLOeX6aylYmy5rMczkqVHjxtKsY
QzeFtC14lUybqt3zgh2DrClJBPeLH7Hv/itSYPZFAzo67sI+O6u8OhzrITVEjFo34RWs7rqgyiGJ
0FO45hAxQQwBwf3JamRxEow9IRH9cwmz60KUhNv9jKaDVg1AGdhOA/0fAX6uSoHY27nTedgqjmai
egtPr6Sdocuu6f/pLwwtVI6iI2jPFiasPUnjOhG8eUQA9BlS6gYUZe0S3fycTmzUY7JhU+exVXBC
ZyKlt9euitL78KKXI5jczRzksfKnzIUsx5NSrH+rp5f6UgWb8ghE4PT7fiLbMgdrT1SHDIQ5CPCi
r+PguLdjamggm1rV+h+MUweXEGl7iqB/w3BItIMeDjBx+anUSrv+mkW49jmeVHbwSTm0vhMgmkNH
PW1QACgg2QisUfISecTLLt1BaGrV8PXK5Zsvo9k8E3uCycvDYSPMVl1Z2hNlI0FJx6N+lJClfG+I
adkp/r6yiBsenQMgc+D/RbwV8ZnRyVz1lcqz20ePj/tWaIe5ewH++5OlZzFDzxQR4HQJPb4iJwlM
kzCpXviUfvKt7dpQw8VdxN3FGTRl+zz8qbBHpATk0LRQdJn9Tf45H81MKG+YtgpZIykCnKJVuEBS
3x6U9ZXPUxOgxpwn43Q/O7bIKLciV5DgBfq7Bapm08lf8aS5Hi161X2XpCEJO3KP005PxNHiG69n
0e9E3G4WT5LR4Ro6aXvttozUlHUUUmfgGwfkf5NSM8FIkoYn79Cc+N9P1cefTKwTKehMaM8W0Zbj
Ofe5uFUZ5/L5UaGRuwcjAGpT/ZOqJTgg9ip90JrDPTPa0gAMZVs7XXuXczkJxWssZHnumkGqYihV
8Uao4RAYUFeZMluaEGDwiyeoFKq+ATpGRuJ56sVeR9bA2Jms4BYYihCA0tZFZuMrvPVhlxZyb49E
km5J8vR64jzKjP0t9R/pC0HOkMmMJM35B6rLlzmyWDzhxkKx+ypPKj0FEGHzyIrPt6K3sgc05d0y
vtG06hLHR3N58sry5Gqq4UUFxiwSJoPHnnxWl5HtWtnuJuxkBZPYxmNe8aVziINfzQpb/S7XYNIR
EFA+tYJOCFdqWQ0QsruIGVUFey1PH/iZMWjY9HFboN0tGdDezKxjsqFt9ju5sJiJiVtj6jOV6Lyu
tTIPRpzFtWfvIIlM3ExLG+Ff6tzGMsp+dSl2nIGAPND4bR7BTxH0cuuJHGzviOyt94a59bxyVzUJ
s9o9RcWI3J+zSP3PW+2ql2ehyur2eABNCBv13qFw16RBWRCbX5k1XsQRU6/ua+6y7+1RwHsUW+Iy
wVCDS6ku/WpQXKbLQYDkIcXbSVzslKpBKHLjP/W5hvitRWMAMViPD8vkwIOBmTVjwBgeiyvzuHfL
mc+/0W8nY/TETjYg+EzugUz3O4CqlCQfG2/Qq7qp3y5g9VDkF6HHBXSe7ZdYymgxXrIXW2m+xCuc
2jo9V/ouXQIPPd45Pimc3Jgs2BozK4duD9+PUvA4hDFyOineuM2eh/jVgIvlBNbzqkyvxpZglDDf
s7RQcvPaQEirjB5Layabw3PTDAGUeiFLRIL6hSZLl0JA4L+tD6C3iz7qzdMRykU/gMHZs67BM2xY
gg/C4cP0duGC2QAVlvvdEWfnhKHfOF5dTXT4E6uzjP5M7sIojKkhHTaA9y+yU2izMTeDpOwSiYzC
CClFrFRlVxuL2Q4AM0GWgvWAI2RAYYoWB4vyH78fdV2GOnREplUdq3D7T715qYxeesVOvkrpIc7D
IrQlIwNhAKJ4VQt6NiSZQbYOacYnci59ojvHlgEbMucRGO8/Wvg1cdaTupfx/ory3SL+6AZ6Bs0J
b0rxZsCFipCmUgQcyBcYpzPnKrJwkS/nVBOkUi3/XGxaMKMbvzcGOuna4Wps6ZyrRj2bAhdt74qb
vhmqJ9scEWYIONwc6CRSSHeqsiXk0tFcyhTNi5++1LuqgrCUKI4GbRLI7a6+MZhMwqQsiCX8F2lF
d3HXQw68+lqokN0E+gu2szdxXkgFfX4ijlFTvEN09UelgQpY1r7wxc/MhHZ2IqKtfTr5AfTzYTTP
mVpYpBaO0E+aqz1NO+1jwBKlzJt2ubGufsduPnCYti1qKoxHefTJo/EcsnEZ98OWodGSPKLSSDUK
bwJkZ5Hc5R794zIv2C0xGe5Hs+MxQBrHgXp7LPG1boELW9A8clTvUIBhySSP4E1c3FNPGQttUBXT
CoD0vSuDsqJvoIBLWy7giHiuzgqtIsudtaEVhW4dZr/QlJzhHYL2R86YffgmlyMpw9Ul7SL2R3eY
MSf1KiVCilqZedG/V8gahsXg26CWzGJIrJNdfcM0CDNtvJeEQqxI4CvSP9kcYHZ9ZKFw6o+3yiRM
p+1pJW8caKfgJoDH+LAHmw1rdxqZ0WqnZmUEuoPmXF5qi7otRsDHM+PprZXWOflYnvSTdP/zG0gV
/xRSv+PNcAuciFYxV0MoeCR3fKG3uk2iMcIVezXExEkrqAGfXINA2Lxu4GBTxdsOcYjAVMdo4/lz
9y54+CFn9c7NDi/BsfGod7CeBbGyyuKgkMq5JfScQrl8aljzDb4x2d/ErzK+ZQEfki3raSHS+XRh
C6lvuc3X2Fme7AHefvgi9IZ26w0JMuzMF3/YgWzpKX0Cxh/HfHEMJqPEfV8ULfnd7cyM+rfi5xGd
LzKAH1ocvPeODL1bsqwjiUoGyzqYR1bGoKzexZuK3hrgNhBtrLZpu/HNfLPCYHNqr0UvyyM1PVUa
gMfvQ5wwhQkXq9X/i/y424Y6C8HNtrS28yijAvzXgOWy9MTpdrSLnvMBi9TtYUslXwOKXn17Hlc6
u7q75jLzpdWGbSERNaFyf3ejw1TwtF5MBtutDewJG+HMjL6NU0TbAATFAZAkFDQlSs4ygbbQo9Vb
QYbAowWbOtG3ivLzO+tcFkRXr+gsFycVD24aQ+LuuuAf4IiNn1oHEhjsHhnBFVxyMQ16VwfK+5Rm
J+BT1uGLcXecDUjysQaA00H6oabwZh2kEcqiXDulqfVd2wivRFctIU//29Yp7GBw6CIFa3hCCS8I
TEhfgUcd7GhTTKJcTXQcHgqoEF4jTChXKTECXKNt8fHaylImkBtOpqhVMVLkFdtcIzA2OTlWthIj
dgOKyfxE3OL5TlctFUcCL5qH47iBu0OfAPqj0LTNXEM6GrgzwcO7JVzSWfEp7n9Gkm2KnQ0Br3ed
gzYSB++BMhitulvEToyThQhJrt3HdBSXaXbq2Mpn5pUm2x9Pay4IV1etcjEceyis7LgaKWO1LRZy
qQq77gx7aE6gZKJF2mpjx4FSJXnSyfzKs+szad/LT3zD3waLKBVxnSTRRYzbsW7TxEUNo9YlviAU
8MxfgK1f+U0KDQWv5S6A+6AoRSiBv0KqXGaJ23VEE3YMA/S8tCmBKJ7fGJ7eRnrrr/uGFl79v/Iy
hdGTGjkWeWcbPt3pGdUfIFdTixkYdcI5exFOs/Ii7EhiU+3TlexOxtH1m+iVR0uBIofetR+F+8Vy
f7d+4HQx9v2+b5h96PxSeZbbLFWQUbV3uSe39/cvqGrQnj53SzkNpMmA7n8RJPdDBZLUquy2+Jnb
otTIhsH87SEPOsiYC3nMDo6GxiUyTgwe0jOfM8sKlgwRwLQyhxippTkjSlZnszzeB8qyc3yGZKSa
b6HhyFIKHl9JSE6kslAhqRBvJyV2ZT1wmxq2WAqn5MhnGlY2MlEUEMNcDual7d7XiI0rJ28rMcWY
/3mxZW99fsSmHwowrWKQYt5PrH4c9UHrCVCjTF9vdBoX+l1cc5WCZCNJHv813jHrldoYsE0fMBOO
1S+sILtVuHJo0swVaWnOisfZvrtUqW9E/Ap9OgBSVta9ORmMOhv+WSen+m8iYoa7AtdNIOosawxu
NTF/Lwch2i/N3tj0xi2sxDVsFbqyQyDt2O17g+S1am+DXVBW4xl3RQwNlYBUhklwIZjY6QrF0HsN
teJzDNuf5ksTNYrkt2QAp7WVds1cbVbLkRpX6Fw8RDqN2GvHdb1i8QasiwzLkOfQuv48BBYd6Yiz
xI6B3NrjkH2sMMf9KwrLaoIqVt6Y970g/lE6OZEuU7QBk6rwvOBIbFK5nMVS4o4wihSNOVjIzYvH
z1KkDQIisWaOhjLIDGnlZRLF6LZkBH6pYHPZFKVEQgXifzFGVzeDOklZyU7GuBmxoZvlhK+V3qWI
4t4R1KvsnZhLWe2/QYkWr2pMprAgnwLmC0QWNkQ7qOa3lEWz+oW6vF2uvM0XplTXhOl9I/ocFIfm
DPFRQKuEbc634q61yq5eAQ5Xx/E5yI9xko4ZyfA/hpnkArFiaiscYpmdaLvTvzgcL/0mKgSDnez9
4/p/HWn7q5FbIGSGYBXXyBmIF17DKqKDnJNvSK8WafOyBy7jUf17thur9urRwVuCv+8WsUVzZBTD
ocMI3ZxVoY0ryeMqdvc886zl65Y2LT9JuyckqyqkbccP4uJ0DyQli40KcHBI/POPuSpfshyHn2z3
yeXjQ7IaIVVmwBEecfSw8F4CHaKlNMBVHn5n9eW8dlu9Gh6vYsPhcodKcnqANOZ2NcgG+NvHhOKK
TrBFooa8IcXgUOCj1MQ+OwYeY7283Fiz2MJeWJdCLP+Le+FJXdiqhv8Gp1qToFPE9ubI0vPUhelm
1ZDLLFKelR+nmY5NagY/Xm8rZv3yi29VsdUQttCExearwPHlDQ6VweQtkV+L4JnFxESZwC6fb6s5
G5rAZfj9zxErP318gFPsNmmIFbKy0DiLso3Ko9DMEfI4Onz1Mo74G/6qPpN1zUZ5uTFh2SnOhT/n
cCDjt4SdOnwY9rpF3PXgPUOyDpSmG0M49M/JEW8gjdK3FCz7APyZf1T6LvUIkI5jXjm0/lf/yh48
MkSMLRV7VGOOkn+Lq1VYqxmjPCKtnBrKx2mOIpk860STW+d2hpjfYtctuud8mWxxkyI3G1f0gTuf
TfgCYqK/52exboRV1+ZqYhYT/zrIn+RrrlfJEf6JLxaz7742MrxDcVWmj7Nf8gUr+DKMNuRC3hzW
7QgRpVNkXCixB0wALP2IquyYyIkvLn9k03hld2+z8yU3UYg8VaYvfGBzRaYXfzcvLKCormPntKTP
bn2shLjAKFaIBG5rJwuZcEa22FdEp+IW4jlRxw8kaIcwo0d7qmio3cb2s7TovB4RFo0iOXE4uQZQ
sfVJR5w8QpauAqNPVgiPEUJyDUwyJgy5q6mW9Xhz8b2CXGi2OjWDpt1GbizNptaa5YEFJ2nrrzFn
LTwcFBemTQnXn2W6zKMepBy1LIyHcqM6OYx2Xn36KEsy+57DwKmnoNjYSdRv7OV2t3KikisXqHgI
zrZcpxHtCJLBsRJUa/dWH+E8GAuJmTAaW1moh0KElCpOhGRUeyrC6f5YF8l9nFUck8LJ9Z9pK1Vm
tqzWs2Wr15Bsd7d6CmepTCE1VWve20NQwcn9zwl78ZP3bXMOA4XtBLnDt/nUPF8aaJ7aJW10UZKq
7ChCIDQC6RqDVSD21faqpdT8t1nQCaxn/ZBc7C8VsSS+j6vrg22gvV+XvipR5hv6kaiXB3qyaksg
Y0JT86iGBXPns4FGtM5PnEJ92B7G+cxn5ZN+Mq04q/xkVkToWNEiY/iU/46Jq7SnVGixJj+zf0XH
3EkszavLOQGsl1Xv2eHM1pje5k+nU5eUOvZrpwTF8QI3S3UbEvHvI1toFeFetDV4uCcsDVQUfltm
LJBFJZxitHWxR9SuUg57DzgpOJjJ9ac5ITYRimnkQAc6SKRgYs/gaUhuTvKe/otPG3aloIuipgYA
02gh8eRUOFLB7ecgK1gQR8xpZob2LVQ3taNWbF9Aw2aaxMtaw96ObY05qaw+3+SgWy5HiN4Gnf4N
kIjeWsmHZUXO2URLBrp6gnADch8pjlmoRCthEG0xXk0Py9OEZeEpwML9cvonWlocMQLaqkBmPILw
/im+nY8bKFbdo/+L6crkNlvpraNN18O+j1H52t7pvg4NvWUchJGuiCcALdDo1X9yw1ezddICOrNh
Xp8n0XKIb1Xvxj7lzxfnrc4CACy+ejw4CmXTX4ZJ3azpPOZ82nzE0tt4lLnRORUW5wcy2HOTUgpg
qHuLBQU8ImO2nAyKoNEloxKPylk/J2fgzEadQPM7oLVm0xOHLtuTWcul9ZFYgqVcih3YSV8Yg31J
mOXZ40a5DsVwHg35pD1cXn+vduztoZkK+Il0mH15bR7vIjg90D32MGMmVNKyp8tsOlDaDS2fUI9U
5bOji1bFj5PW4iQNVocFbcUBA/mk3BXcPd6yvYHnW2a7RhbyEIDfQ0x827gCMeya8SZm6x8cW23H
ZK0Lj/dL3oO68V0oKFdNC99YTaLb8RC273EYJNolIuXr3b3LNV0yQVaTI7qgIOnpdLDm7P6iwPkz
PUuR5yF4HwHkkzdG03V+eAKmAapgD2i0CLGR+p23pfHdJR+Y1pQbSE9G8LJU9593FYAhFIs8IDPM
zx4woTcGzmzTY3lfLPDfcN7hKvM0OqYw98uqxIMiwz5YnG9ePH5LB2uKA94S8HTpqigrdkoTrVP5
edXNU7q0k3ivfYcT1qIIAtFFIVRC1KrAtP8WBbmBz70+UK8a6jDLGJsrUEXYObigjRNSfd7Yko/+
ku3ruEidU+luIK6CkY1mekwG8jZZQB8RFRmU2K3ATKRomB8u/qg9pSGsemSVoZsmVBIAK2DDwR/j
SkqppK2H4EFvzNc2hpSFATf+Tq/d8oMX35m5jmOm0fApKKzPEFvf+XzhJlrY5lmychHWv3sebhxE
WhdFfi+1L2JGs1ItaY+Um4jzjc2Nq5gYlJiULK0xPu61SJ1ha7Gpj32QaeFhsIbOvuicwGxo8KHO
OJNIV3tdTP1xTvoUK4ai3OHS+7nb3EnEVt/iyohzAxDThSb+AuP/s+YJbfbpcLdgKik/WVZSXTHc
l6jf74G3GlgOG2x9Qvwc3S88A9hf6HWqlQnLJoKI0ghvP/25E49puAaRtns5tVmpuwiQLwUsxyMh
shSg5TeGfT1r19vHLPl+dRFMnVZtWj4IopDpvSJ9p+OPLDNoglE7m0M4Ept2MQi+iRASnF39X87x
yftWOiOLnq9MXw45AoL1+PFUK/D8Z0Xwn8q1B/oCNpCc37F/oBhYXq+wWIpe1lkGhiFe6xP99rvc
hlly2Vnfscj55V512RM1ysc9JtpPiFjNqF8OaHUoWcoOO46toVkQkOubUuj1dHGKeQdbE2zEM8iJ
e9Wqf/ZIJt+lZuWxWRi0asoQeGMC5OJBvQlbBk50q1dlaVQalzmsJc6rRzMTD7qalPe4Ek4jkUDw
Y8xKgooq0AdfM1NjV/KbnleCWK1JJy5aDQQ2FPLFHAG/KWvVAD7+DtxXfnzQcdu6o46UnedPHhFX
a61w7KCCVJoJpRXwzeTqoAPCH8UPWwMPlAF1dNCidCF0XO97ijMuvoKRmlPek7Ehu1LT7JaYOP5L
OkcvtvmctIVCPA/qykHzPZFbncy6AR+jwmwo//gmZ2Ui3JEoaCnx753HuHwysSGiYNX0Nf/NsESu
DvmT9PFxlUMrKqlMEhNRHwBEfkK7i/5jS2PClJhyl4rSgJRnccIG0fwP6EbuzwotrEAiv3UyKAnM
dX53iQHgq6ac/q46qm0MRNWuoDbJOMD3hRXyN2B6flve10G9oGevuzXY/j6iUHNzo+bkzN9xF2ud
SS3b9Y4UwoEjG0Hez3P4vkK3CArcT7iObUV2XPiUlDZTy5a9JBPSqIVIYbBug1yxwJpsv80gE95+
c0SzYPUwxPvN9WmkurH9ao2wkMvLwENGdA8XewVco5DG8+LA6tzTxazkVXFIQ6tbWorCp7CUMQWk
O4lsrc0Fx8us053vH+4Na6AK32ITRv2lNCkCaFPW5pAOlffHK3kmjaB69Qcr+4abXvhkn3GvJ+Ie
TOw0b1fXxS7x8a05Az6rKZzAh322XELH0KG6FmeJJoSbbXtbHLcRdi2/o3wOUUKUow9agpKcy0UN
zcpAcOyNJFZ8Zp9s7kDMR6WPqNjD4SPcHKDKWApWsqbuIpazgr6GMHQj8oNU0fuuQBq//Rs0piKg
wJ5277s4z86I/cUVQqCvFKVJ4aEDOxJBEuf+uyMbPghFYfz4qdxatRCVBh7qepOPMsL9mPBApNwU
f6S6AviW6IiW09LsRGZRSCfWJ72gomJZ4iP28iKSpl9Kd2OQwQ4v+W3HF4QCY0iT5Z7m6aMskyh6
YXug78/yGGax2f2IF7IlraaiGBCsmPJWesFFSsw1Y9MDCqYkGK+EmBQO1ab6lb7SFTPXpMzV6NWf
tAhAMT/QMJHebgLk4T2NDdyOUcWafj0fGo6Yx3vXfXoyacUQq07291klg26Icv0MTqcEtfWR29O7
c6zyUpBDYnn2KCIqkYzcNrWMVu5dOPKogvkrO6jdGMMAmGP+tWV9KgcLxM6Utn2yKSZEOEIFHURd
J2mOMr8F+wCZ2Xd6uSA5yLwaHT1zW80kP+04bBeW6iC5m/UYT1IYDPSo4Ef16wc+yrXZSLRWzsKR
Zv/tizX5fYcDbgWe47BmrBX8HVlspxnLz2ajR2Hlq1SEmH1wnsyIHXR1RmMZzt6zzvJbeGGQAQ+h
xjbvXEEL9Qd5YvsG+UAB6cPUq4rVmxVHiKL/Yh1cWR3dcFVVUMcZEZj7X9QftLa+qAMWpgGiAs1/
GGzrrrDRhtJJKTZhT3Z4Ym0Qvm0S/TJvOQLKaqLuo8PEOy9cdys1rtxSeshY4Pt0saF7MmFjlEEs
vE71AaOB0yQBzuImOALTkMyd7/liX7MzMeYZcvEKEboMfzRKm3+zBdyO0vTyLzwF10RendLMmwnd
Qu9Sm6eJXDSRvTVwiDaP1W8dC4JAwm+kpYOPTD1FHXC25NdbLu6rF2bLfTKXMEyJBwYZ2N7XIjDS
VX8JHIEZLdV2ZPY+O259IgkNfPzf1cF8/x+nwD1XjDdRbt5xxOH7Bpy6MEiFONM3DBlVIPz8djeu
+TTDttccPo4qms0e5Pbu3gOYpXH13hhWGQ7BrsX8Q+6c4uFGTkaHtvqzyLWJNNI90vfylg2E93id
X1R7IktA8zCjxJrzZcl6HtJ0YLAAU5QEvqju37+bfUwS+ImiOraGOebPcN6bkI972RJ+ity1mOET
UPZ66DYI+rccPAS+rv5GRl7Zsaxbsp37giu7hTGXavwae4C2t9xvmjehJMad7LtTzTUITJkBU781
mypr95zIf+bRzGVanJyzBGw/clQ2ypEIE9khtoHRJdilmTTQCndKDQmjigDtQ+oJVlnL3u56KMmf
TyniUMnwhUgiHy5QgQ8aupnUmHFVDOAFGnJXpPo12ojwbm6j5+zLt01jrZew/Iv85y26nfIk+pqu
BBGmB9+DeI/E3OAQvQI5PRpysS7FIog+QyolOggTxxJ02VIQNy5C6ArW2wADTzgKWJ24s1Rp5oN/
9X8FIySKsvdosedmDTXTX4DtnbwsMsWPJYOWCHrXiZApSYCbeH3REgB2NTFPrimP6iWmIPJB+FT4
09ZuB7snrNrzH9iJOFHmeh2mOvQhCx3V35BlW780doNBUv+swLo8sPr4vrlFORoN2fYxKLRgZLZ4
jzjKILSOjZ+Im2slWFl4Un31d4VUd4BS3BTfJm9AN4WqSMkR+f+tNLC2BsQ4ac4mgMweD6TMUFZN
tAZycof69v02oHUCbXBqDKkB17ekjtDbRQnyvbtLL4HdrVaijt1jNUjdzqOU6EsPvvyQQ6EqBIj1
B4G809FCtJVegzJOac4TRDkN/VUXoZvp3JrrLYJF8/Ck7ipIXTeAPELkSPVfm5q4Tr96TmsBE0QX
bN2Yvw36xchwj/wPEhkfTzAeqbgt2IhYXFfWSK6qhujHiUy+Y/FBLHKUibBWBjeZ3iFUwwKLyg9X
sT9sG21Zb4uDtP0cm5+APaSPDxAtHa6blhn1+oNEOt88mlX3ntdQkw2AKjVQtXxDAD+iRetF9vjz
Z5UlD7yH5ntRzJg1ArS377dr1SELbWW9sKL5Q5TXQb3BcnsdIvMatM1uBgO9ZxLs2KXwUaILN8T1
ubQAaeOuRK7CE+NRJSnJolYlc749bwU2Gy01DgwkJyGDLuZQzm/YmluyeMwLjmT1leRBUWkK11lj
f8pOutdV+AtjbOtqiGDk32T4guUEnA+IKm6+wSh8q7G288hdLgDPI7QE7VnymsWOltFCc0L0CRhz
5b52zbgJ2bMjHGEqepguxED92cb6khfbtBigoreXtFzH4A+m4oXcKtKgwNWstfcO0AhOqi5v3Gmx
w4d4CkHtqJBdEigsqUAIt2FUh3YYsOro/iC4By0msjhExlMdNRkqzGNkmGvDlInn2O/MoDD0Dr9u
cgR+z/tiHW6XPpKVwrYqcZprSRTq5/Kz5vR2yryECJ+4DfErlJiQZoAWaWUsVd/2rYf2T743Wfu7
3ntPxChyZP70+TvNAXd73zlGVaF2V8Lyaiqv18NduOKO6kxeoIHGnfREKwcFyfo+wa1PRondf3jI
GlH3BGwsm+TvK+4a3zRLUc3XoZH4hza8ZrJwmvaokxTB1p1R5gINSK4gzPp6cQ2MydN1L8pz2ro2
4tj62ttlXE248O4difrorN0oQI8LOKq3qRl/EKufMZPBX6PZmq1bnTb+XEjUxfMinCNPdMYK4OO+
svuCxwKvgPL0nky01wzs/EpFkTL8ha9srwEhNJwqBThqMukv1RyvBy+j+QUEYI2styxlk3G8ZPo9
m5rn720PZ3vlpTPih0U63M8EC+jOe4reqroOLDX0W3zadPTFmmuHOCz3um7qzIBy2SNtjNMy909h
Uk/5N6yueLnD9LnMxhzleLHqdKnkVsQRy2iV0O44g48i6PChch0hLwHEBHK22ix0blxJn8NcpVLl
02zZuSKLv4xnQkEUvV+Azq5SAHZv7AlalxY4qHJ89oZn97KPtg4pM14aFj16TYFUJINAOCFOKH41
v1d9y76YrTJcnXu2enZ6lUAc4XyLRo+JifWkxJHs/IqRIxgvAnhxQa2Q7d65HvXiYpF1PbTAlQ6+
oRRfYXEs65elirpMUEA+YI6sFoUIyYEMrvBVEY6Kp2bIZin2xMnfhgWZY19BOu7qh5EEznIN0Zrp
J72Xtdv1ayamvcbIV9cPbm2XMZEK7VpUNjCu9B6frEL8px9mKyJAaAdYTVpISg0rO+xOBh2ofO0P
00XkW5SXN5SG5TwKREe9ILATfp9hN/jDQpGBKxSZz9G1npCLTMMHu0KrMjn1qglM7EZTEHGaXTG5
ZTC9b0GS3P7pKdqkiwQETl2vbrrPALhyX8YILWVxgd8haQupfJ6rJPms8V0Ev4esrG3MV/KFL28E
FkLX6ZzEc3qCt540T4YH3lQO+mBAe7JlqMfN1gwSOemMXjJK/YzqIjJ1yKL8XAjszJqzHUqaFHkM
E0WSqncWNPVj24bNo5z49ALJoiJmKQDACw4EP1IV3k+MLd5bVqUKg6HXFfAUxIRXMHExwpvhtmNS
96MXFvR4dbA1r2UhQby4i/lFHSx/11Hjxuus6IQff/mInZy0FdqJiVey4wYb3fZoDEilBDmc9Rbs
vWp4CXPQeYDQXavLTeE8PVkz/dAjSjEOskalifMMj+de409Brzl9ekAX+ylmnjf5g/ZTVT5pTata
Zv2Y1NV56aNYKrk37w2OQhWEinxm/NSJjjGuEV4zkuNUHyGvnxneQbuRvFzLnYv4TmShJ+DLnmG6
oTrWz0nLpORci1+UNVmo6AmAFuVLDu1y39Flta9ltorldrM0cRhsG2w4dB3BGfb9+DPjAvT5YSXv
gnBhyed5+quXJQPhEwOXowtQ+XA7WzXxq8dFp+iHYGyV3TDpR4o7jehTrq5LOZbrhgoMfCarfE2S
ka7sCjfFOENoIhnx9MJk/gO7IGB52BJFlrV1UIT4HYgtCQxrfyKDwFoYf3sDmRWlV5QxaR0pkw5t
LO8+JmvyEGmAj82oGuVcDj0k0ACsT7wPby7feNjSYlPrEpeOMaf0UqSUt46CI1yfQQcC0FKP1Te1
0u0o9JAKS+91+aL2IiyCpPFYHI17hA5753k2JWd93zLGQl94F8RRA1XJ6I1MCcnme0SBSDNwCWKc
3A/j0JCKz7hlObvta0An8byoVTetCBllxQCnnkPQ7fuaZecLG4Cebo6LbgWEI/IOYKi995TTtzdy
FdNgryfe94ypAd53LXNku6QlJrn0xkbbIlo4aaqtLkAO8oY1VbgFZbwnMHfe9WmJJMjK/HtYGfcS
yDGRaOBNLGdgUYByK6ArUyeqdlRtwl+lJSXKr/Ul+IU4/e5PYhJEOgXoWTTOHMiobo03aY3slh2o
KOzBUYhD1DLI0MGvMn0bKkdGvuxO84bOcLS0MMWVKJZD2RG0dMI5fDa5ox1B4H6tgih2g+2hICez
L7eJ2l0Ld/KkXW5ec103AQR/fp/gw7SdLIR3GGuA6i6sETbILNNoXej9a76en0d6bYMiyhGBFWoP
HW21VfqrytObUm6pWGYeSRyT1dUC0+Zytr9YG41nMTVaL9IiRi0658+lOJhnfOuKnUGUAQyHppe0
fkGIKH7oDeHoPIk2W0nIsnBs0HxQu2ZdxkMD7lCOx3QPyZ36A8XUtrjKY6UKxixxO0MliXkVL2Bb
I07FO4ywxScHvPeChOKwS/gB92mIz38mYFPiiaLbmWiIOj9dzs4/uuVdLthAPu1rW/MjREw4jEgj
HWvu6zGzU/xwwmdUDkTjnhlO0AW2EdBRDEKsnfuj2up40c554tRpz3iHxjFB3RlpvA2Zbgt/0GUx
uHU2jecwvB0gGI/zNuxkd0UkKCbkQLDAl3pnVeyRbhxf+vzISYGcd+PbHMAygxeLtsK6Fui64Qm+
SQRsmSv+OJYUO+bZxiIaEOmT6fST8ftPdG17l9GF1oIT3dosYttboaz2pqB3IAD0a3/pdp1Dydj7
4eRCbRDjQUUoDsjSkTWS8zJMVqZmOJWWb5VjE22NtKlSqnZnrHZG5iqFxg/cAZc3/7xAN3gQvrJt
2bPgyhzq+r4+cWpbkWzYRDDFw7yWohuZE1JXdpfJA7+vuHWsiYg8kqp1yPtk/SYfTDodST+VWQVO
zQ+9wt96nCzMsSnsPsSAfZpjNgGPrVEihdNXdLuXoh4dqlVgrfX9OCyUVzFfTv5E/wlKTaYUquHb
VSYYWH1h7V9tIQf56AIX0j9vGzoyyPpskKrGbztd2v4HYsM1tuAXQu0QQOPqvcdR+SsLQVuZHKg0
DhczmEHpXBaAXYatRQ7iI+WajBqPPzd0BmuvJIQp7fC7JmaejMPVpxjawFiOI8Sk4khXV1roHKO0
ycbyntKJ1mq5dSrZoMEBg2jQx+fxAEZeQHAF2kc8cwmwlqLsmZWR0hSO9A7StOyB2K3Z9mrXJTWc
s5jHGIRo2CH82AuIBDTmXiqKS8th6C3HQlXBkCZdVEP0k2a8tTQJQQzb0WzHSrfpyWPHaN7ZmAyb
t91FrMR+KMCXlROroo5TwHE9dH086gp73yfQ0u99UAd5da8XLlACFKJFxv99WwU/htXtIZn/g0/r
i6+idoRPbIugiTVlPVtoiZNYm/FQKXmfLWdLzXRHT0V9N9F5IXSqp7NcipvhQMCTjLRcJIqn0VAq
mLk1LMSnrnpAsAE8P3F0Thu++CevVkvV6aNTTtiDlYyAQvPP3dHMFn5IAi5dwyRfQrorFT00SLKB
leEk+5LhG/I6oZ+uSiTcnXnkErw2xh1Trrd4ggytTib3O1qigfW0oW/V2iP1N/ytbLqC/olpjj52
dA4bqLPP26Mhl1Ak0fN3ksDvb8O/t5/p9KX2yF7BFfNrPCdpXsclkhVTBSxC+6abp1bykVMinYi2
XDoRIN9oODOIYIkJ9p6ntC3lHvBvoasrwNBxnzHwkx4SROdWg9DkhQx26tuHdpdVRgFu9RelhZIU
lP7pBSJsIX/7qEpAfFztJKxaOg/+0jvkLxBwlB31evZuDHursByROTIbeh0WY5jnCSzrAaVzKnYk
sSlwjeAFWAAVK0Xe4UzJrVp2GksQgByuBActxWSbvUZrlHBO6G111thWNMZT0cwt95VhfSfhE8hg
kao8QMiqZbe/fqsvY3m5virfqg3VgS5AhTpENBRfkCfkQOF50+jeTVoxF6ajUcYF+/ABVXeVKM5T
0o8XhQnovz8WFcWMa+Xox4IS1LEXOKxCZglQa/gXgSZEzq+vnYWWmD99rY+BUp3PNYKc/J2JAAR5
vutTsxXm2nVcmB/aMlUxWSnDaVP2LP2ivs/3l89ErRw+QD7oe4BECkFZ26Q9BPm95ZeMtEMsrErV
mIqza3UP1wE3fH+VuVYh65qi5C7nLd9AxyEyWB+89saABZdHwc8lq3R3Do/ovOByZ6UkyzPoLlwT
QyrKNfo8B0IsOywljGcoLs2friiw/P5+jz7+R+eAnTtErNOQu7F/unaBtSjpNbt1QKgRCUVsirLw
wixzjak1WhDAv7abOvDtyjrvRMia1IYfR9aQewSJz8eB0k8hCf6qW3xe+g34BsjbN2IzZeLlxW2m
gNcfIHOCJQ4yXqMkgsYQTdrhVql0gkn0OGR4CequCf0Smi6f/zL/rym2ewLFFULPLhVfAdy9Kei0
tXvcXA12L4jYSZVp2yUZHxZhYejXrmnjgCZiKd2zRHvCIPO/lUO5/Qe7Qxvmc4ACtnRwTYrDdh3x
his9ZuuCwgnXak/Gksr8BsjHRcy93pj3wSmUjV1IiObpC20VjydEa/RYvyfooST4PNVLYH5NOGGW
RQ3Xez8+W0m+ZsNBI2Ce0anikB/BpDiOlT2a1RxVIokQLxtFeywc1yZXv02mN85t7G3jQZ7cuPxq
KApqW/LZI6PZY2YS+cmobZCC9q6SlJhmm44ms3FJtcqPiQ8QC6ztjfs3SuxzP9On9ycPRz6Xpla4
lGuSNdOj0GcMsF2Yg6Qi+an0c15wha1HKoH2JLgHI3TuB0etOfTUKzahR1n0RziryCBsxwIrHdAC
3LDPSOQaxM4GMkqnV7g7BfltXyGWQymqscAckSZQo08Kco6jEdooyOD5Wg9cFcuPiISl+LOQ8BnW
sYZi8dWDY3FEDuh8RLLxBrRhcXmz2WjeyGTnnHzOLdHxa2AXAresdqKbMZC7PvRzj3EtxZce7J2q
y8bH1pRl7do/XCprxIMizTlAFQeezofSbPvKX0iW3QtL076BIv9EIDE66+oqclZXIBNCTQ870eew
FmdOhPphnhHohyyBi5MOXqAA1kzbJB2ARKfcxqkSpMFxJvoZTtikRfYB7iUORouBG7eg/iva0u6K
WpHPqcSDEw6mDSY4+BvanoL7VYip/LmiSrxaqgi5EhP43nZ3Cs13vmXaNoyFmkdg+vOA+MQ1b/RD
nx0VDaf5ClFuBKutpehoS8jmfyFhXbvAEJPfYr0Dzdj16p5z+9Ud9n8ZqpGHgTTIpH8TdOeyUEgM
URH+Aisqcrvw37dYJM0+CXsq7Ol4lC4NiBvTDRHJ604GM8kQxZa5c+NXbK4sLsTwafcZOSx4xO99
i+LD2NtNI/aBSdPletw3cTSDhuKjnsctSfx8uNCJWoBl+1//eDEm4khsINF+rpNYXuTTTpguX1dO
E4yEjrfu5fLEmDoVfHEl+ocZXoesndcHcc7Qzcha0hxcozXXaXgE3aRNMpjPQtUv9unxsanrvVM4
5RAumH5u4FlMObigMGuTnHOH71DumVTKIC2jlkDIZs68D8eK+jyy6uNStDT54bcyLDa3UMEv8KOA
sQFrLbbScXOMOei6itsbTrqUkt9JoA1YWhjpYxf7OTPgseBYrvWgnUxoTAVcF3/aqb1/5GON/7sO
pF3F+qBUHKWJJuaD1D52hXeypgjl1z60YUW0L9M4P+664nkHPnpg/Mgp6yIrPczlvgiISneghuJo
nGHy33r8vFvUnKIXYCOI18oIymOKu3MHNYpVCNIKe4HvIFEJW4S6hh7kKZA7/AyPY3EpEeKG8qke
BUtug28BoTL1LXqTmDQDD4uZlz0TIVoVgcnk3SIdKorRKYvZT3KAEYhNeh9/IAFHVq1DMBEswBi2
zwF8lxrFQZtxZ1zqEu21zzKWGRnDLpWQzaCLnMrkhSOOl9127vrfoQ6f/fFVkoCAkLrPubooMYaZ
XakId1kTJZLe2RDR3YjlANRvKwtEFZxYbTZVUK4tkOt4P2PLpRpirF9twRiwThkIsywnvWDB5SOD
CiMn7otwmsXYJlbZoITicSMAHrLUURxxOzYgKuoKaiwKgoh2Y4y8z9IijeGFjpFpT/4SRAfrBK96
zqIWVgBsAOmkDbifJm6iL0MimlIMSznEhyhX0JROYePgOSA47swe7g2Yd8fsT/YhV5ztCdwqnbNs
a6tLFbs3UyRFq0XxpLit+8I1FAcGiovygD1Wreokk87XW8j/JGgOnHmKRydWEh9MyxJyj1FNxDi0
i0XyBRNa6bcMaaS8mecnJOX52dEQWux3Ey3Bhb3CeOsZpzIWhLFsB/GnFw0bbHXIggJfzAMBBoX2
RMjVpTE1uKUVbLgbKT/5/ZFbA2qaOlR7ZSBYLbHMYi86hz6E+ODP7iEC+WuhhQKeKOg0O3J0tv6B
rb7kQPEzoonqCLthGXEXEjpMsiATYZg3L69QgMbmIQlHExHBebD6rflOEcToEwwS6ztxAZemumLG
2vBWQBQ8R7qzcQnFVezzfDWDJmShS/DOcOiXeDqSefUaFxJwijnwg/y5HLO+PSynx38SXG1Uq8fa
a/L/h7QJtb0GvDpVCyJGMUJkTsCt3ztlOiNlN5AyTL8/7ABXsl4Ks+zW52dV329Sw6fkA0o2Txyx
RCl2qUOdbqHioAopOjKGQwjkz9zU6BfkFWo9eP0Xxu2zcLzRXnsBynWMZLpk9DmYDf2fCgz+2+yU
a+P8Rhbd5CD/G2h2u+5sxetr25QXYHkWATyyn3nKj3eb+Xfer9plEOvZpuoiF8UDqTmjCIVEmFuY
iWmWq5gGptkc8w6l3PHICK7mp2s7llIoYEV0YLbdtkK3RHhiXLfgrpjL1qr9K7xjNPIsFD7r5bGr
gvPqhX0a7kMAgYpzSq1wWIy4K+G0vILUwkjTjPyyf+KfMErUfDnXIp81ss76u0iB6cX18H5hzeas
x6g08POzVXsaNdfbz01yHnWVutxJhXEKhpJ7xMVCmSA7ZJWq41IAhyHm9MOxsRM2duBESa14DfXb
jS8QwX3Fu/QoUKv8cX65j+6RiLElrEGndjIiOeWMFIzntFbPGcjrTbzFd/En68/oVw2CSPR6Dxoh
PG9Qf+y71mke8uVqxwVxu7xkOgJIbxM3swWOVffFTt7cHW2Lm87oXg0YyfZamDxK6wUd/LmING3R
opHTaAA7CtBFB0Gm8J1ZZ/k1oulvz51/Tdxg3BLoBpZCt6iMoGyqWVOPJ0Od1YL7vCyFFzLMBmn1
qPdW1NcpihgHJhJY4L0WqmBzveEKoXTPrVgdIaUoHrrKGaEk9IeNBu5c5ChEv9Lub11kw4XG2hU+
tDHxVoCGr0OY5R3WGdQlcqcxc7wA1o0D36tecr2cEhj08UqKK1Su2GV15r1ylKGa6ZRWvfA2ZEjJ
5Do002xq17XsY1APmMJc8eqPTB89I4E7jcgnI3x4OYVv5ctaSLCLh19XgDoVkBEIo78nNkQAVxkR
/yV7xQMrcP/oYtiaSkzwrCbtt4jSpBNx+bBeRHhB2SPWTFOWcVZGkwa7fc7ODwUMzIRKNeW8fMda
AzwWz+67AJUhSk3aFryTiZUQ2WAbMK9Cmn5MXilNPALjQCfl/X0MqqSbPokECps4L3CFyaTXpGqE
ZH2IMDkRJZlQQ7U9Sc3ffr3a0BCEhQVQ8q7hCXsjUBUqo8gY2gYCgZWp4ycoMPRwu/HihjroNUDW
HqTenMPZ211luuV2skvt46mLc5VpoC+nK1VP6IuztfoNdamVN/sIAnWnJcBO2RYvEN8zLB77M1cG
jtYja91kEbFKOEhnTN+1hzzVM8RK56pOLDNtC1Wlh+Z71NrMhJ5VEYnXXjg2/mKFgIbX96KInXBi
TUEvxN6WZLzqrsh4Al4tfh9NEhVz9+ovioT4m+Ch4EqjILfTDiDAwCiSN7mA6GREljRglY8ppB/j
+Is+WK/wQq0k1aXG34EMzwNXXqQ1LkprWpGeKN127szaQ9raBBuPswAeWcrVO+XNgMZNH4+29Vh/
OAnG9/hQbD83BLo/uQ0NYmC03e8rg9yS9Mg0qpGuVdQk9QcFRaR670fe8Lo+Nx7yPn5ME/wYxxKW
RgpfpIdHwLwrCBELreGnMUp/t8xqQRboAOFKQxSF3YFaTEVfOHTJ5DtWebWm3zv4XrL/HMHgbj8M
wDyBSCiwm/CdflAEEEH/T5RGAm6JlYLz34HL+PmfgCQZiV8Otj+SdGD37GndeJJ8wELgPXpdrpFg
1eJwdDPrW3OcVROpFw66mh4gjHbgbx2rMj2yGjVXsi5yNkj0MW0VZsGYN+iwkMRrDtAOBlF619cg
zrI+efZJjx1RUo0JNfaCtTAY00gxf16/iselxftK6npHgCHAskvqR1CdIKwCfviy4fdTdb+diiGA
zyqvXydSfVXEOXFm/OUmOd5NP1ShYVeI36WQwAfKCJzNoKzDjYxZ1kLeZjQCoDCBnAj6xub5ZI+Z
dz6LiOUkQ/0NstszzAJvA/UxxWn1vgdjZNiMo7ZSxYMcPO2dEmN2K1b5FKJjL2iTJD5pSGshYlng
ZmAmPyZDVB0PHGN/AzEwet6iXvcRHDO47ASNiBukHR7N/ssHwuK61qeAMYzFmzMD1h4fOsVrF5oU
VLai5IyLnMZHbnZBO1KkY+Uk2twUCATG3wxg3pW01kpslVwv1BgCSzLv/dRnGrMyb/dbpb1aOsGj
7MFvaYInR0ZUP9B/4Bhj1EBcx4TARWjypnbd4096c9HDmPmM/TBcO5J6JFVU17WTM35CxJ7MZ5S3
7TaIHClUtTKqWu8qiCxdA5P9OVhAhN7cM7svge8jCdrUsxpTWY266eykI/NArVcGECw/GC4ZEb8X
Z4bkJ+KUdqvAjdGZeak5YuTKLNqipEJHdpy/iB5+PQAdxEtqW2abGLmcOYruat8dEPnE6UiaOdCg
u8Cco9ViojB1zIHZupwxUgZ6IYx+MdJBu0Dchz2qP0ymKsOzj4+helaIOUDDx7Ao2sJoeR6FD+pI
8rFdNvghJv1M61/b+BGj3Abh+VW9nyxdQibNV8RWmbtfOS51twqyCi48yd0+6mhQcEzw9Y3fLTE8
7fyJNrXDHnPoDVMJeKdVcsXGHHfPsViYcOLFIQXhTYTYw8wusyvA4NmIsvJszs+nzUOkMLWSPD9Z
2LpkUzmpOtK4xKg6jsieI8fa62FGNUc39wD6a/J8H6MVKaxbi/2foHIgkjaERUsTuyQKddpeblSR
Z0oL5Mg+18lo3Nsf1fQf/yy6aNqsogQtA22f28RUG17DaTkMTs4sGmsvFF+AeHF0J5sfjfEI1kir
bFun723LnNp2jUU9iv4XIZvPkLHlqB+HzK+vGBgRDLQRjFDmhM1GCobAlTMdzanzV2FlGOqx2z8q
ecpfotSdo7TYJfVcZOYM/QwjL+wMO0STa06IMph50VtUxZEwjwA1DUMk0sWtfcITJ1oBJ85oYSOW
7F/FrXJMQWOyg3GmXuWz1PmzDgJKqu2ghYAjGMJjc/3Tl85Gi6MzAWroeLd20XRiydM5jRKkiPwg
3Sk0IqZzW7qAvl6N1JZrUdwKDxK4MXTqFHGQkWbL4FunezbL6qQXtpiciv/p+FvSFn5AHiGqugxN
tpBjN5dlkNI9cSmux5+L0tFhy6Sgcz8qyEQcXkMwNKdEZR2TM6Y43/TN3muhY0QmhUlOh9aEe8cH
qJrJacALMyNwWXL6OLNA6dvLjs7ckJF7x5wc590UB+IsJVeitEtHcirvr5crfJXhs8DmxfNjQWqE
Se3HbC4QyBzWw4pf1aN6Ol0e0SOg9ga8SvUmypocd64oCgSZVdHF68vSCe9qNpjr6cBX0Rgcr8bk
OER8XI+zpnchCD4XbsH2oGDcNGkd7ag55RLbMZ7rL2Hxmo+oxDfmw0T1e6HP0MxkI9ilkmxxLhS+
1KYZnO+E95MjznLfGod4690ZcVQSr3IjoLT4di0ggbzx2uyo4oTrtJt7zeqMyHpOQ+pnmr96X0MI
SDI6j/bkf01rbO9n+Wj3XqluU60Qp4FsnZXvLrmnq55fgUby8BOtqctLYVdaTky2yqvdLqwgaWk/
pLA38+oN4jhpzBEqP/QJUS8sTanDsv77xQLNDy2ahIh6gzfFKCsCApmhUWGCOwqEikCNmHBNL126
1OBToAhverYK6/vixDIaxiLUxkSOMDiZnUTBYKeHEAJxmeD2c8mRMnZWehSF3lgXRR8ZOdBIJ7YJ
FjbLt4fmUqloM/BZhVPcIZs/pJlnxmitUYpZzNtcU3LCawEoBSnBBKFmQ1igxg4rhtPtLIYfZFyt
/r6jJS0i+JcBhRU8v01S3ZJ6wYOteaaOzihJ9X/JI9WsLP1O2c42YyLi9jeq0NnR9B/hiWTZe/Nx
sHo8y0xypE8zmoBt6q8ibKNJ/k+x/l8vkAuhXYX1FrKoUAh+vRHH5R4xdM1zWbvTUUer4XKK99V5
nZFh5/1BJK0+dCkmzhAvDl9czu2TZz5T0ksHa+mLop5tIRcCu8M/W8jYIMohLrjdrDKkb5EcUBcd
T6oHmGyazIqU/+HeDmN3JU5lmFzwXTVhDKQx07pKv0dvLsBmis8jbM+IMVw36XCU4Ag0TpyPyMD2
2sc+5SQ82Ruony9WkuMszeUMZk8TkPox4fUAO4w60BbB+6esoFOmESwIC4E6tr9FrDSZQyVVwUWw
+GTYx6vOk0GJkeR+Nwm4VN5w0QDVUsLwdq8ZwZf1l4beuG7ZCX/CfbuduVSl1N8p9C3uXnrieTFT
wGgOvvvFDZUoruFjF61OP9DxLZPDr4aC+054kPT/h+0QG8HokOzFqDzS2gn0tqUuT0r9aw8bLJAZ
NehBqk/qBgy2kz8G7xWbPD4XO6D8hVHPGrEuNNS4xd9Yc3wi4Sfpz44apalxdOgE6R7LuhpyN0mw
xQ3IKrhaB2gSXiMYHz8HIWhDvdeaE9PL6HEtNQWYQ9jM9xwZo2PR705/+UV1H/iBqBAiGNN89uGV
b3KiV5PQ80tH2pPUXTIyMbYQ2Uvk1TCI7h9ia9JX7Cn81grxwDrx9tRnBgPmOT/mNj1fkC+gN1eq
rpbhtHui/9Xu/MDs7WDcK66VQcxrTifiC6yALK0kwYFo+owHEY60DghvLLGKS1qDi9nGBA39OCLh
JJSuLJOlSSDehLiTFNZ7a3NqDzIQyDddZfRAiyvO3yVc5Pa1RjGYHI94i6ntDukl5TgFmK5h3vGK
G3Xutfwk+bk0SbTyDRDKL3lF6LjGFVrobb8IixiPB+eePhvGxzYp9Q/4mge68UTtXhuJlOd8j3hJ
1FxW6Ew1ADY+HTNctlc2hIYl9Hy1GDR976M1bacrG695ZqTqVQCNnoqBd3/iV0ZAB1F+vfHWTep/
Ft7k7GSyjdt5BvMvhBALOy7bjRIH7RK/9hNdaCdPDXI9RI2bMkLsN3eMSV0ScB1TA9GDDQEAXsze
u/c1NzuNUdg1qXHuMunw02uGyeTaANFrK9Y2ha+CdVP9OaMF8JAT9ebHOcoMrTnowtlCbjsotB71
Ay7gzPkD+8NWl84UGsGAqaWH4C8g8XQdm/Hd5t9tA9o6Z+O2AbnB3Md9tT/iXcMsRYrWRAHKb4LA
+Uz5gwV6GqvMKQDfBNE0P/c98sf8Vjavk5wF7MQ2qq+HCiPK6ZmfESpP6KFrorKq1CM7xdGJs62+
pon+NOpWfnvxjkt9vGGSabCq/d1twHcc2B/Oy/vXprJhlF5ND3VOVFMdu4859izAgZSXmGxUkHE2
GbCtodgPiboV4K+KWqca912OhEncpRxxMUrIw22bYmY8jFcwSnSc07Y78y7nG/bGxcqgw4wEXNxQ
RRz4iG208p04ah/oSlOpfJ6K+nhSF8X6fxXfnub+YX0JshhBg9bDLdX8mEpGP9A72g8TztA3y2bD
JLmEs/Q+XffsMvhQ+QXOOjlQNazDOSXFph6zQ7zlJskQc9IIbyB379wdHIPJv1WQii2IHPnKRTj8
IhJEiZxqJms4vibn+cGvDcDnOfH+5FKYieRsAbgXcreCU0R4nt/JvS4JnuFmEshJc/CcewpVbuEr
Xl4iVMIpY45pCFLoBsjZnHsWCC3ukGuNTbdGhHC4vD6xARi9r8oKZM0POlwvgwlabaC4doGK/2p8
SpXaXhlRAC8kVPhVO18rE48SLL36wEQwjyC45nYm1F5mInY9X0SlT44Xcqm20iq63v1oAI43VqCd
Cyz8YC90PxEKjZIp5Mbe+t0lfMmb8KzOwOdvkucpkJ6MqQ5kiRqD88Wmku5hLGNsvvzEoXuxot0T
tPTu7auEN8bHUmSX5Onu1+uk0opoRVfMVz+kIvr8KnX2kZDP+JbvVdRaXAMjPP/i3shtDT7ojnhC
g+2w82UEJXvQsIonr/RA5WbkL4wbb0GFeCcYh2bKJenic12h0QIpDAewc6VjtnMYMl6TZRyQGuAB
P1IaAJ8tY25FIrymdPowLhR6u2Md56ogPi8cKpRDHeuTExPiIl3I2mr1TIhzQFqlGmJxLwO2MqqJ
3nsv7O51Rd/w9yWR15zWzSfyQXU3ycrvhyBHzalbGWXZFeF+EYI9IDrJWSV06PpNBZdGkfiSt4iW
Xr1zPsUQdF+oNl0i9vV96y+3ByIyDjT0QKIHy8S3lcBBeSVFPZlsQ0bqwXijEZ71LOYbQf50Uf4b
gFET87JkYYrfhorFXF7+fRsthpgkHB3F+sZ1JJW4oCeM+BoEzX8BZ0sG+cUcZ7u48je6CDt00Ou8
/lKNFv4dGG6fkZuNwftQUtGj0WBRIieeDBCgUSAGhGILf0jaq9OC6pywUoFBZ4+MbZARRtu1GKeT
xyzqWXrt/Re+NQx+pOfszkz+uD5BRIiIYh9+5VDy1Il1JsSWLcG+b/OWLSGTI2QKpF46qC7jBtj2
Y14XpsuDaq2G1txdlY6ijCJRqGAMMNdLepy3P/7z7+pWB16D9xfeBlb/BvvE5zPQMBMsmRMmbZ5F
Xy5t6GfULjNUAqo3VqSmaELyI9iJxK+BoGUNjpMNNrVt+wBvtRt57y26F47PWotL2xkgSoQVOcdi
m98Hk+ChxgjB8CKlU/fdo+TzUyE7QVAxzpkD3kyjHaPxjsCqEt9Dpf8MfwyQtPTCYlngt9bSrntn
Qd2rdgyfmawfF5EtQHQvov8pKX1DDqa/FyFjQqGJZU3LzFcnVUEOXiK+nVrXLNGWm7PDChwNtBnf
CU9aesY2xpjU71dRm585Se7UrK5Kd78eWaSjqvxjHu0WTusLPVmA/DviPkaXHMaaglQvRgOxSNDk
BuViDZOYcchfv5Ri6Qz/MD7bRgLI9FKTx1TuvRCg9pDKjpXLWGRTPiFEj9gNeeTBxESin+SmQ8hR
jmFRpvj66EGr+8D7HKZbeJE5FUjWdwZOpzmUXons8YJPFDYbJ+EehdwXT7ZnNCnwsxeBfi8M3VF4
T6vw+5JqqdEDYv5hkdi5R2V8D2vWQvlY643qFr2fUeW2Q9yX+rH194ZCO7WkZ7s0R2Vyk5p1MnX5
HsCev6KiNKOcDP0GVL4y63G/WuOxqGh/qTBJ5bmB7pQxxsvMLOW6wUvhfrcYg45PjaTn+3S2rLC3
17YdyGvHGK/9p/kw8q/bT6B95Xt6SnD6FMC+cyIT74PGZd0D6/iuS256227oW3TFn+aomIiYGmzF
xweG6wG80stn6Dl2JUA1Qxc6/mqxVfwDaW44PLfb7sLSPyLRLkb9d9x3wkyxQQy/xfGeZTG4VChY
d8UVCwO3Fqo9nORkV86D80THdJnPS/EdQfsxnBjxaGr7c7uc+6ELmUikRBvxxFr8vLsHx2BhKT7P
Cc5fgoS7lzw5gbKmnVnTYqyG5kyddS4GwoBA2uD6N2qhxFSh5igsVp5OVj2yj8GYrdiJnDy/yUor
te+Y9c8NOcWclRDLKxh04V47Lg2RM3rgjyT3GrA7yleT/+4uU+VFoSCaOO4Bp5Zskcwmjr9wseqj
K75xuGDeuC+AQUMV3ERZXMmadGQnWFgLOVd+S0KIUt+aFh/moiHHPOssrDeeiuuOuQ7Q3uNp6WaH
NGJlWUG1Qe2uth8iz2jv2D0ccghGT7dZqA8/gdBgrpKVuBvfZgvEP5BTf1J5wL2xzMQtS64CUAD/
ho2dvq++gP0CISnKce5Bq98mZtEy5j5gTrCnzjE3h4yH6FEhXYtQ/GqJySTYGI2+vBRQ5ltV0c73
eBI9HJYntb5yf2MRw21FZ/7szEBZaMRnAkhgDncT4V3Nd/oNqqlaql1M811kZJcshALG04He9h5O
6pU8qODwR8tkxeNiz4u+KZ42zpIp6bkNrZ+1Sk97/kaRSzAtLeDJjvj0v8HsIbtfqGlrp0uozmGH
b5FES3bm7w0AyA1UQqL0YkJ5tRC/4GDxRWmijXrEQ7aTy0jhsrmLzXS5IdJsYCgtWpZik1PgwWLc
vXnGJhev4IdT3KA1Ma6kBk83ssUBMUAE93HkBRtLmzQxx6pbcOSG0RUKGt5Cd0ZYlkRhWNDVOErw
omplOo1OqrKeuje+I2vDRYaLn5Y60b6wz1sznd7CaYmqNAqNjAmFw/LB3XHuEZz22E1BkUOZ1FXk
5SDZNqMZf15rL2/3H3Bq6OVHp8iOnqWbpuUp1B8mQHpkY38k6FljXLNcBJpeSXhkks8+L0gxf/BM
1xK9G707jkPi9Ph7f6808cSHJ+eT0C8ClrUy3bBRksDEuSO8uPLpVF+czQUHpunu5gQAUwkZmV0G
LA0w/kvkhflW+QKYwnGOh/QjJVA8FFaaAbOMnCdH5zlc2+MavV0aAQ6DE2wR19h+lOFc3r6H04m/
epiTNIKVPdon+V8eRHRbvqwaOX6U2W/iMKDZjmy9Sk3giKcFYn8YnHmayxTn3asKNFWUwOK7hRU8
Ji7gnrdm+UrN5QeJQPsh2qXNadHpId/6FbEuJVvMR1WOywb3KUzh9tdnxjwVhiUF5WMcOZIe1i/w
roEgwBRT/++MKeazJAOFh+yvS6MTdCFEN8ZyBc575UXoUws5k/XPcHv1boBWhIX+yhkRz/V4OBxt
zTi6YK4EWF42akVZMHgIeb3yu1mybetcqky7bfnWn51AFz2xXRgmQC2GlkOfN7XXjYiyvDp0Bet6
sUaAmifvoKqEPyGLsQP05P2JwKBPQZqMeahcnNZm77Rla38rTtQZif+RPzWryMPySUncaJZdSy5o
UzSA9FchPX3ay1KXTgEXIzNYd3njs+jiM5oQScY7qX9vAtNsa+sVp7qADUholojDZ24nOrGVCkyb
oLKdSxL+U625Ql05U/dFpVEsoIaZkDq7Jy7Pa2p8Cptv+JcREfHvtM9uP+xLlGiCsIEhCV1G9t/O
WfnX3axxav2FVKgNq/vNsZqqo5HbnKMR/yz+YiM2QSspSOUNEzf9MsMGdXSNQ1qAw6jQyU+UIEL/
obQvfyaLBKmsyfvDi/s9wEF6WsUGt7lQGxd6KBRHyg+FM/1vLzvu8ZVfJKDysiE1U7Zp5Xnp/EFa
9/jmV1cKhaBMuRB5Ekq/VdX/EORO+w5YNfL3P0n7wrMluqUGHhvhsPXRveFBmKPvNGI4CqEB/TVK
+9otlsUzYPR21LLEc+S8fHMyhj3WTBiEfleXzvtweCcqZ4u3lz/+igzUAWVMWHyHxLq/IeDI2jQe
cnDVJxKi6a7SXRhq6jSChEyHfzkqzypDa5AsqLaojlpZH8kDCBHBDWykayQfTymL8E09xaMMLovO
gApzL3lDhHKT01AaKYcp9ZCE/M3mODZiP6h1tQaRhBGpSHgAI45GYAX8+guy3YAeP9IA9aFtwcuA
mv7qygV7EEozsPVv24WomIrB55w9NMNBlObxFOryUduCZ+jwHlIGfzq5SCLsXDfC3s0FqcMiB/K3
I9FG7D0IpUFAtgD1oyYJPVTJ6z9SaehSpCs/40gnrgOTInQECsfkUfcdQRh1YyhkUvgwbZYCFfih
sgpWEXTUDN5XIXRwQyhK7kqyuO5R8kraEvV3gpSs7oMo9/tkgHSJyjHjXeZ1HEQaUmBIrgoNdYPj
aqFm8oovzp7wFAc3LlbLt1zUfgRUjjuC5XAR0y+Hl6e0EqbmE3VH5YVe1Wl+8dhsOHQ51L3SYdvM
jTk2JePTEYuRVQl2KknfXqoQ2Zx13K4BXeNmRZc6uQtzAMBMymB6UZ8AWyXF7DGg1OUHAJCju/Cq
wPRg7uZZzLQTRlqD7QUa00zo1SAwBNoGQvh91Cn/mwpoRErOale8/KneDOfE7r2weJey6Q4JTUo6
e1hLP8u8xGlrn5KItPsApE0UGaPH/qskPneoHxvG7V4pQJU+T9ueQfyUI/EMxDXljb/3yGbsrzEi
EQ8yqI/tQoy0JfqIMPl6Y6/v//czkpxfN9Ge/FnUDVTtlP9CDPxGmz+5zzoOz8YOaTwOD7dfI8WN
yCDovEAXo/jTqdw+4YG31+lvvPXg5E9YuQ/tW4rxQTrIKg+g3cqSuwEBUQEb4wAfOypzJvagIB9w
4MPguAu/etgDrFrehgu8LjEUZephVDjcJwnIDB0VR66IEMuZNHrrFqdacM6v57i/d7Nshq101R9h
IStLsyyPUEE3Sa6swChne02rlsTmE0mWkCZgNmty9oHrxkx+cvoqHXK8XR4u5sHvovtA7RUvblBX
Rw/oOx5FLbrpUyGX8eAsc/7gAGSZ5iqGfIFJ0affb65aNwdlFZwpyfi56vyt9cTLmYeoylgQhcVs
NG+bbsNUQah9mymDtB7is8rPtBSCkYdSiyrKaHx5BcrRH6oO2rRmf0GxChBOsoXX4cZ11lQlAHIg
z+ryhuabCmbObVC5h+0bG6x8pc1paTTHyiSkihkf/ryMeBbhPJBYrnkCcyEG4pDu5ysL0vCBH4Jn
nTg0cdCc8TX9qMumcF35Kg9rcNIrEQdIAqz0vJSqPz4YmxildNpb3ebTVqUQCnMKYnhSBJmZ/bOg
YfIzfNn3ucTub9VA+4B81vP4a7UXMIc73qvUxbYdCqGh9QMnV6XzZZoxycEntx59xT3K3YKwDhnu
wDFhakMOyOI4yNEt4MnRAKdZk1oTSEnnVRBjOyKo1ywWT7q+hscujYkHA3c3WCT27TJzxtG08WvX
+hvO5ROyGZPjOYQLPnq6JjA5GNikaPMyH22SuZ8f7nlxseuuEIbPNV2omoMmvGwbIDlXKhgRI2+B
ct4lZkhggrMf9yj7fs0yYnNNJ+G7SWgrLeRWqoojhhDSPzven6A9OhQICNbFYCFKavxnwd1pK6sA
aELze1VM9+c79EMhyWnlwVjHL67q1JL5v67Xnd/WnnfS9hViOZ6cQwqsHAqAM40+3cGsi1aezTTE
cYYJ7p3UN6/HecFScEywpcTX0myylJR6Dk8m9XPYV6WOqxX9tOOMehNTh/K6VmihnmXynV6Brr/1
j7ALLrIhcIGvB8/tjS3QDmwWMg9T51TsA0K8+SYpdzXQrb329IkCpnxy9tj4N38Yw814eE18dsZc
554MjE/9bb44N/E2v1arT2JuW1zbRnmSgUJaKwTFReysejK2uOaTi8tU2cpweyldAS16WRARdW0Y
du09tzuFOYkB4DV8YtReT9YPduuYi86j4l+GyhaZ77PNRQtV1nJQsYlRW0oNz1/HB0R1Oamxqu/C
H3vB/hB0jcV7m05T1x6h8WtwgTrRUeAu49+wv0AerhVyGtL7B01s1zbqs+xzPHYYqD/qiQRTADXd
zmT2hBzbfCK07wtl290HXMJPiKqz9YZDkIh8GBC9Y/9BTsEtVz06zNkSTphXdeBgM+uW9jlQzius
JHSVSht9BiVS+nDCcNhwEuAZ99xUQ2l6QcXKghR2l2ByztGiKZPPJec1lS919xNXzVRL6XGE+VDX
EGZ9a3PAd5sKz8jTsqk84Mtshu/TAX6X02jXpy0FAGXJLhCWGNQl5M9oVlzyj6F1LrF098rSEk2w
x0HHODLFWAkG+W+54L6igWyMwYi/uMoUkhN3oSnErzef7FKmIHSZUCDpswbM83gOdh/8Pp+uIAZS
ecgv58IQIrQDoHZMtry0S0SaHVPouxD40G4WaDDZKdhQcsrVs7sFSZMUB6Kn4SPFfndTrQFK81YH
2SVlMLyszDpDL44mfEwE9Bq8WOp+CSPIsxVBCYuOMuNgt2+dn0LjkpDXzF4NV53QPcOuhCfPem5O
SMo6P5so49UNCmiRoKUoMf/9UszX5hYlcNZciejMxL2vNuf9fupausUTb8YIAskYjgia71fc03Wc
dU3H0mgKWt1RvYvOrZpxCB1AerfQ/pKo/2k8DZO2fNjj81Vz0y3M+DxwGPBnGhtM3SVxzqUz7W+k
Mw8QIKqbvEHGpBNk2zueby4YNPyIKKbKQRXE9GyUouypaETgSXtoSrE9/+0qRFnLJLfjz8GP62tE
kXN2q3c+nFi/kFZHP2q7Sfw17NkGxMNLrnlLyDf5EHm2xZYRR2kxZ2oceiAK62dX9czl+2mvHmKb
7+UBWjXQsiIYIMLclEK6gNx21+4lk/lF/WBufmigIqHnMSznGXyP0FW41ZH1w0QUENZh8tYkbqUn
OrOZfMpnA0ThMjEBD8brMl/A3aNxDPo4BhdaJgG9ZDGTEgFOowCmT19OSU0Bhi4iLi+lBPGYQRhc
L25/smnemCio/frX+MKNyi1a1BH9WAM+hzwdzTkmUXtQ213MjfCG69x2MuYnAJCOdIq6UosvUP1Z
zxnQy8cf+iJpV/z1swv6HjrGF+g/C6HjtawN1O/i5B6lwSFaU33JuC3b8lJ2c2Oc616cmYINLqL5
Qd88S+nO6b518pVR/IZvN0n6BXGHD5+z0IB8v3rMEIj83t7KH2l3/dYtSR2MlnQKvZGpzlDSmRKP
vmj+pwGfDT2U70PbTgPvpvUcAq90OO+xThL4FNbWQ4B6daLGbuNOUla6w/BOp8asGPfW+5RayR1y
weojmCVWu5HzBF8jYZlR93z1lZAZlpCxYcZxOodDo8c5ItmRhOFmmDro5P+YY18EE4eFnwRGC/Xn
t7RqpXRS1YLLawR436VKY8pzqFKW6jXg3N8ccvBA+Vy1X3O+YiioXBTCs+zPUT6fIMndxsxE38+K
4u00fBJqJdnYQMAWRgwn4H3inYJLmv9R/S1pBTCJMnIRkRgUWAtjZMg1pdH2ujKKayXdxSczHFlZ
ERIVW2eILekI7szjAyTQQaitV5rqv4Vcf47Uc0uGfFPKu88u29+kh3TmFRCt1GaWHbkmVKORn+HL
It2go9nQoir9Zle8mnYvGH6bJ5wTbicN5h38fMf/cwJjYmYiNjmRmSbwJ4YRJCYOYRJhItMIGoZj
y8thvOnlDGWS9voT6pOT7cApGLthd+HHuaircKWX6bNjujumqx12aT9hC1ZmXWMtR9GPmhKCwbvl
bDE1DZGSQ9dWVFGVOkC7jqcjvJ2fcwRqW8auB18Z9NPr/qhWpPPOHfOIrH8L7qhLwWEKVtfke9RX
aPxt0L5hc0/APTwd6eIJkh6vly81aAu09PfVISyECZuvpk4wAkU3mcEIzr9B3WUGCirJkN2pyGyU
bm6mMHTralTPeHI4QZwDjVLvKYHv9Tp18Dv92bB+qqLlhozd6DXAZiL8RRp/dNqU6Ji2N8deWVAG
nKkEKu7UVaMVC2eWBGxUlVwJBEazYu3EmXF11MWJ70ThArJAjNnGaYXFMTzXnmeic1C/6c7WnJKi
i9PFn4aSvSaTe/t5nyJIpjCwNZVc5OzM9yYv/1uQDKdzT61LC8BtE5e/XW5Lvu1gIzn8kNFQB24S
F+dDZcc+porQ+9q5tYs/c1YFm2+l0E9j14wJM34mcgwaNAg9CzNRXvfs3RVFqBpMRnzI6Z7dc+84
3of2E5g/Ksu649sW5EZOQ+ioZHPIK4NeqsNlBhyNQ3qzU2exSsVu9Qi02shvYR3/0K9Pa7lYXEsI
C8jyN+uBsy5zKmMcOCAgi2i8ICzc7MPVGgXbMHK9eBX7/43sSSWyPxdbP3wpGh8ZlNI9vvJ2rRcb
xSpvZ8GBN9UtxwIGxr3SMkn3hBFuDLSCjKj1ITNIL83oPWazEIpMJLw3OOHyipL5fN4/z3JuhyVy
YjsqRP96zHL7OX9N++mUiO/Xa/uNPAFQueteJnXMIUCM368Ea6kE0RuboqcTuahf1txgs3yEIk0g
ykbaciTqYHwk+ipbgce516SpSR/U4ZTHIWCeadDExvXxBjddHX4onZctbwnL8Oj2+DQo233Xnmg6
5wyLmkimoXtacHXPxS9fzAGkYm9lat6A6/JCfvYh65zYuTNsFsIrn4XiRXA7N+yXYm4cAm6a4eVW
Y3Rcg8B5J8lbjSHrqsau0B8uVkj8qKbZjNxgLubQlCELR9gciw0bhVfgX5G5r5ZfiWy35Xo52f7b
7GH/7LxQeNqN5TZfJL0izlfYhK5m9ouLBos1rKMpSg74xXO75jKt5M9DpShBk98ds7ycwINKuBld
Ia6OlKRYRlWhu9QEhY9PVqa7jBvNrV4N9Ame8FiJFi314oAXyGnH03xQEADXlpl/GN4QIWyrD4Uz
eFuIFGt0pCRIANn/N4VWa4NPsqG041Oiz6qgmtGAddhSSxcIn1u/aeyxIQTV3kEpio09jZPkbPM9
RovJgehZhHOUadEXzGwvdUCmBt8vMJyS8s3HivTSqITxlhYwbIpTc73VKhylCmJWfDZCE3OYWvwk
rxBnhGJdrj0dTiB8rFxekNJJrrKIVdJuIA8bayeArEeGVp9BI9ovdoq9LBhuNZSpEhjvJSwW9wXm
zuyUjCWNUNxrJi8nj3s1ezyXuEBJlZY2uyCTWbVW+nI/lU4aTsrcdPA/apwC00+9xqjz1hoA3csz
lPQCw3CtYBf6id1M9I6zC2ZM4fLXZZ6UQ1kVQXdVjE3S4qgtdwz3VGP93COJrgKRcGvSOROyFR4Z
WldnJtWgnavtIcPrjdXH17GoWKXZVvd2HNdq/euUrMnlMEJy16i18HMfI7gh4wv/bS/X2DI9MFxu
Lh+X6ZHi8Ls6p09wmSB6iaxZBjlW61IwWDSM09mqZal1JCix52ffasFu995F2sxTovxvECclzEAO
EL98BH/waKaYUtmC8B77FWWeI6S8AMxqwov6C97fAE+pVn9qVChhoZxjMFm3+lXrZpbXR8jiL7kK
I1NEYbGps7xVH8RVK4UqjZ7PyyGNCvAdEHMR2B791NfEBwLy5A3kmBk/UPylZ+nwP7FcALsJWqT2
grItTZuJE+hQm4E3Mw8ITgetoOxxXSRzjVkqN4BN1tt9KUBpQMaqsMf3gyj8NUEd7aYrjL2q5JEb
UCev1aPp1w4Gikf+vgePJqxI6LHwWSb29GhjpmTdnIiqern6ekdm2TVV6SHietcaeaqLtBXJ7mHI
s+YzCKfWCDhPrlp+7aQZo2euVzBycsZAy6HUwiPFs+lvuZyGKRtbSERPqG9WZyBRyg6SDjp9q/NK
si2deM3ualddWzoQgkWIamDmaRbPnldqosXqw0swEoNzItIJ5js+PKnrMVs/STLdpB6deAiTvY92
B86imu/RVRPtPq6FgxDlfzcVqaSwymkdoJR/G0oyl4SNvocT0m6WAqRUocN4blKWcbLjcLb2Jo5u
RRdsz9G5s/5H3DY/j/T//bHmK1PFzQv1Qiw6obzilEFelE/BC8D9m5CQMupuEUI/tvAu8ay4HFkz
OMQYcfC1MEV7FlZ/CNlI9HoPN7uqMCW1RFv5/fZpEYnT/9+vU7sGZHM0fggG4I8HSrtGdV5tjpF9
6bZXBJLjcp2UQR1QhoQ1M5PMDmAf9JpueHYKX9oDcY0olEQy8bT7oIyR70bQfE6Tcknr7YZ33z1l
Yg8KmTolGxb4NRwFCVdZNVzSVmUwzt7V6quEJapetQH50FTq8uXjEhxQvHN+k2Vil0uYZRDE8K5N
yvZEiSK81jyC8q8BVPYoBiYohIT/NWeR5adRgnkkm948ie6zFmQV4XKtTkLVmLF86Ps+3R6sLlqw
D0NeU030mMB5cXffSMZyVXJh7DT0yV4z86kAx4y0g+Ir9SSiWCkNToOmfVLrFJn+sPJlGZnaPko1
/f2Om7vurot31zvnNs6uAAOPQcj9ZBtXtWNAoZL56Fo4/ENo1mBbPTLfXnWfulbBu643WhUWXsPA
sRslmjZ/N2fhXv4pW+ZLf4cm0yMbZuoADQG4eedRLsJXj81hluDLcXy/lZfgkCei7dJjnyNhniXD
QErKQp3hQcPrEtnOF2D14BgUAhMNSZPHuu8R3+uuldI3HCK18MI2imfLdThiYq18hkh2d5+fRhai
bcfuLfnhQ6MrqEbpJ7YvUR59VTnUUhDgKy4scM2hwMT/1Vmc2pfIauINTkzK9/CTjTQ4JCoUE8cB
a8FpbXXPTGA/dDQMxxGAn9FGplin9eIKnhjNMPnuRidV26hCp4PPf6FMmHTuPEhmVUSCSMgZteT7
hBlJ3AjfSGIJHruHvxkqU8woMvDTO+iCrpXart1El47JdjUdKnD2fyobNHTVMl6Y6H6h9bestn0j
ACnVlhXQ+sPHnMdpTdyuMkKb19yMspJrkede/PuvrSPJS6t8tvXz0Ol+CTnTuIwJS+QF9N3AExTt
z/UOXTiEyWjm1LxA8fFh6bhYLgpBKleEgsEp7LgAVoftPTd9vcQ+LLGPq8DGs/iL2S5jCIqZe49z
9k1sLcCZEhY4x6wOxXnNlqg9IRar0+mVJCWP3SnzaZq1px53AY3HLaOUkq07oPLzzFdj8KpXpl22
cWzIzRgUI9QwXFvoBiVii965jhNJbgsihBs7PUuW283y2dyG8RzxZDaMtVGXaH4JytpYSv1jiHNH
Iw8bCMu1dYlG/cG7fphzMqDQclP3ZDDPk46WR36z4OHC3AqlH0z5IK32WD4wZOz4sXDcppALKLcD
eHKVN7LnbuG9Btb5DqTWlNWdZyolLillo4mWkEQaMhSzWl/YqfsmRNtTosLvNnbEy26VW1N1U/3T
DfuCphnq50Bab2D3DwgJucCjWn5GkcGSKqnpdaUXDdFLty5CkM0vhT4HXcJ9HHEs5bnAePJT6YJy
dLRcOH5t009gSUiVfBmOwGyAQ/16wAlWN2tePtQAu6ogRhjC5uslGLJ0IvutFJGEwNonpdxWq3Fa
z1qzUgUQJHP5yqE5aekIgA6v3BdJRA+aWbc3IanuP1utlJOgnwsXd+cA3PiLGgsdTwUv4FzEgDUJ
ngQGAo/BFJY9FlHfCRkyTJycG81NDpWDkKKqPiQr/0IHsrXQbdWsnwFjd4Q2T785S83rig742LBN
C8QF1M+ngCHjaaVDfmUoA99FQd0qKmgieeOz/Ec9HkC65v75ENomjBvSWAi+Efim8xbAQpvW9QE+
Q3hbdG0u39ZTC4eoKu1MJ3AyzStS4NVwXm9l4fDvVNyl2yjNfunM/S5FVMkvBYsvWj4uXYcOcvUs
K1BiPqLUSI1XBU7F+9E9ug4mgPi60O6c1TCAYZdKKL7X+t7LJu3tZEwILeSKeDmol1q5hPj1ef3F
cwIb2mpNbSh/sQ4BD7PyEA1xtgt5s/Ew6Iz9ThjIOZ6qd2nvKPe++XlnW3lCwICrYR1m2eVYgpk3
H1Gbpd7eoiiefUniCfAGI4znYgY7noUREvoMfz5ctAtOqClVU4DKLYyYRXalNffTf71Og1ARzr+s
btD5UiUI/qvX6+2qMWf7ikqdx2AHNN/INxr06/Ub4SNdjbHMuRGxi484P6Kmh9dIoolpAXgiXF7M
Wfrsg2Uk633xhCXOwrTG5NaQuK+bchEFhW2kRm9qyTz6fA6dD11z4gOsDARDqxgrazOqajP2HwWY
j+AFWOm6/ADomgEy+cWOn/kKzKeRcrYA8l1roAvIzImFM7sRj4oJNFYCeNHWHS/HrcEWcHEc6Ab0
qq8lilu4rnI5i0WRN94ZtgKaCM2hox3BZppHTxKJ4bnzyaI8gg+5Yc3qiDoLHgsqm0vC7YgIexpC
de2vfbi4ZgFi/z7XcynmLMKcprRlkEAhz8h6RSipzrVoRkgsZuObZlgf1QV28W4YX1DKH1nrGeMv
gbArr1megSRoReiN39HP2LZ7cPryI2uiruIh4f1/l20JlnuWn8N/rrYAjydYaXd0olr6F95bXjDp
LK+L1l8ECBRSysLufU1LMYLB/F/r/DsYz7EpufAG4ZFzAwg8OMNE6PQG5LNhkRt6q0VGfuEn8bmL
elwiB/cQWfWw0NCvkIt8QNW6VXKnjgayHsnMpEpUBWheri5x1j/YqdEWWpyTOg8PLKlkVVB4VdCo
Oj4JuJ8SeUi7jZ3N03eLdk+sm3RZFMWBVmB+T3HwBpTStk47ahAUGh3I4DmijpFpTRa7V4JcXyfn
Js659rnVih2q0yIBEhE8rBMiK8HVK3T2zo05Pic9zeVJrsjDRTJcpgGmMVK0iBOCSiW+ySqgaFRm
ByZJ9iJ/YZZ5AkZuuT7fD9Gk7tu/KDGLQ1ot/fFcF0Y4g73iJqepzb0oisSTatURfTgHB+2rcjGG
RUkmNgppXKfM6KowvfdyLFTKIuYT+TkQUQdL1q4JwMq6oZ3MGmSZ7Fg6nwVLrD9QFhaQOTiFNQ/+
MeJLjf7bRc3BL0NXO4A48RxmAPwXVl4Ln9HLfWEDptlcgP7PeXvdB4PF4EWf3WVTaR4PjosU548V
Q0tEDG/2FsQUS6SFOIjVZf2FYSqcIkXlnjfjbHSd/ml78z3yucjjC1Z9WHGHfz5d0spzRyetyjne
b64ZnxOm7PhVMsETDrW9i/Nj0jrUvPs6Hm0xVm0PCZ78GOZ/1ikXrqU0zviN5opW8wzzOFgBGjdz
xhVLWkFs/91Cb7ikBof1+7WLgEUyebQRdOnbqO+GB3xZF8F6FcdcQbwRwohnBFYIg4swBIqUk/2O
r0nOxlx/yNtthRB/cpiVFCIPMvXRDu5OXN0CHl6x9pPmWHI6RVWevXZRNz5I5br8cMh4oCIlEBJc
IIisNcUByOW8cfLVv/Dk+tNhqEk1+41wEcD5E//9z+lkYpHNfiJA58AApYDfbz9/2Cwe0CNLKj5/
X2KF1g3BcvG6zbhSi/Fv7OVP7OpwoCO3iTHUeOqlMoUobqVG4nPott5bkuqh9sAfA65cPr5by4UD
X6iu7nwuvWdxpVIoRhakFPvvkEqqfWhRyx75MoBQ6skOu+OKKKHFpsUIAnjAWU9R6tNJv/kwuIkx
QcT24BpNcRZ+jKt0xMfxnC/yRmm0zISAEql8HWr+n5eycwfIvvOfylRvKf8ljx0EywKeu8lj1u8Y
KG3t2TSZmLnFekXjgShnUAP6lZi6JZCQVXd+ICqL9pX3CmbH24KFjU0/+z0Tvyhq5nvKQgcxYEb7
NMy4bcFh49FR5rtwLBpqqX3DLSX8L9ZdD49rum4hPmi3Gcs+JlOJ/AclT98QI8ImW4CTNmCsjxTn
0pipKtFNoXM/59+WFSdboz/5IMNp5NDEmhqWeE3g8QKFNklZqUNVoc2hYFm5cXRJzZwd7D/csAN7
ZwgSR5w9QQzsDi0PWdHh++CRy9CNHjycCBuXDdhnmq0Ux/2hJqM9wPGzr47Narpw9t4+7gqtGRk+
ARBsLtOcTFCUZIA4CjXZUDXfRsKUDQrQH9aZNzmRinbkowkphavazvyRNDLGt5KCJxaQ22lfpu2d
XymzGj2HclilMBCR1UzwcsE/J9k10oy+rlJxVnUB+NKoLa/YHKOhF7ghusJ1YfcKVYggRbLYrV6h
kw836i7o8ljVCjrc7tyCACVyjeq8HlqBXpchMrEQ/RQwh75sZNIf+SOFUQ/kljdJKDcBbbuOkreA
1z/WabyqGo6f4Ns6O+fE6pjKzXZ+PzaUezLSbIh1k6U0QXLXoXR6oi4uOHf0rjYZtnRAbkVvJUOn
hCA5/MEHXU/LIOYtKhSOZg/YRwG1cfNxLMh+O4kA7nnv1NudcRPTGG50tpCOmmDHQbshv/2szLBB
Vs1gyUef/kpf8Ee5v0AFCHcqGiGYyPp4gM86YpavwFVMuqYagn7oH/A7r2Pwn77TOZNQG15/pIXV
ejuNseq+Vn5u9llTDq0VHgMG4eOd4PZWpB0B5CbLxVP/D+vWOUwibi6Db11WGZxamjrykh3WuSXF
aMTaUXV2C2ZTdUR1fWAbL0BvqBtZ+8FGZ9lAnBI3UZZ1fh877lLKoEUS0ST8/0pVraZW+JNT+aMB
uOeuoxm1TljkaUiVrNpDLI6jNgq7YMkL/PzLYaDIcPPEFa73oiQFF9nAxd9tspLe8zxHzHp3n0Tl
oWIAupSMyvdkLETUYDo/+sEryiCx3HZSd2qDvs46niUjsHSMDtEfsy8f6kvg252Ek946MP8Jy+nH
qui/hdJx0LgLLtT3ZrrQVgA5v/nzuciWrkcvKNd91+E+s44qT0v33T/C9juOfpXy/bMTwZ6TxycF
djM+hm/TtHrZPcK6XhWL+aC5iH1a80z/8mUtavvKRqyb8iogrkmoTH3H6Jt/cT+PBo2rpPf0vYS9
bkDVE13dgAehUTims6VQDCEcWSYyY/yKQB1IlpUipoO+hnuH/UYkGpmzS7d5NrPfYIqSLupcnZwm
bsxqtym97UfHYRP0S4wB3GaB4nu4867UaZMliMnj6GSzPV9efgifisIJL92dhXjM107Hm7vPpfc+
S6LbmUrkPP6Cwi00sfx3eSVdoCSmE7/2Hj/YxahgrUmH/zxGTJLGrbM4Rn+HPDtrHlImLp1AddKe
rBgoWxjO/Xo+H42A/seU9WV67l6mCdQOYRHp/jQk590JiZ3cG2G5TdMIvZU8r+2iiiARzUEdnDD2
6RKp6XuYnPjth7myAbdiztC+Rk6fbUGDy0qPqQh51sE+jNiE0bZDyPyJj/5PKUw+qPWPWrYyhCaU
0te3C/NrboOugUzvsxoNx+j55WXmidhlLdKSJVL2SgyuAKkMH7rGEjkhrlj3O5/aZwx3sC/c+cSe
3qfXKOqAEqI89pDKhW2/Yoepbzw4y/2IvVTthVVA1aoRn3+uSjAdPIz/d9O98zBmZL9LEsJyhJWG
9vw/aKEkdyANq9R2jKxpwj02tg3fnO33w6fmnCsV+6sw2n9KYBNXIcH+cJJFP3stL0bm0cxjJg3r
FXH3ywnhqE4RB38HduBc/Bu6MyJdTOXdvrW5NOLMQZgLc1SjRwbJV87K59t+uZjDlzlroG80CBzc
b5+E7n1inhFXqAIHazuhculFkh5VrkartXSeCw0JeSla7A5JoY2ty+rNlLTwn1wdcluqEr6+8kZW
IE0awleCLSrhh/WKfncJKcNqEiVe6++ueZ/epTSamoJ5nYJjr/0zQapVZlun7qTU0CqWKTqHE+Py
iKRC/jLCtxm1R5jr8nb/XDoBh1nSNRj11K6AUfym7LwO2UoFBDddPFt27kfTwwBk1mzgLJyKjnk+
hnzJcQIVJJkOR06Eidtn2u4gb1RJ8nuJQhspsypo713LiaUfIhMzlLfxNaFsaepJX1f/uCdvXrWf
X5XfXY0t/XvG0YNBjSM3Znxhm4N7XYbs+szvBenlir1OFbiUQyID2EMS57h04GW7IhyjUNia/wIb
VK0ipbI2sD8jx7UkVgjdeVWiSGtud6hxey1HKzbNSFygkTkkRhCRUDfMVg5zv4MvDNEsIp9FOMtg
tNQ5H4/qHkFwbyYD2UiNjCdqXxskkWs4DK08axrvQRlpwljyA4j01CtswYdOKF7UXmoSezIymxsy
uN/wuC0FiMGFdOk1KPvzIcnxMVxP621d8d4qjfNKmQEnOYlDbpXd5Zm2EjKOxKFOk218r7Nw1iqc
rZtZJWLALG47VaNGWCz3TAgEyOdGQcDJoxqgvx7L0h0antVQAI4OBNd7ZQA4aFbE18/pNsu91eFb
199uVmx2a5f3L8voVIEM+P7r9ofWXeqEliTtvoyIA0MCW3Vu9diND8CHG6tTo5HirYKewFfx0HjY
LApznQnxmiLkCzq5vsUIcvRZBQLlGqckuffgbeW2vPmvqjjecRfY5sGGh8wIg3a0jgv0GwwKv4SI
b54+s9aXWn0KHs7lZE0BwwjMAJn/KTt7DtlUmIfw9KbQmh+EUtLue9TOKcr1IC2HkMK2Ku+0K0Y/
I8OgDT4LCd9Hih9nnWFwoJmn7jFxqGNJJ052kngizKWNOd6NyIO7EYsj1n91qU9HQikS+0t0B/7X
A9+5/VZSfjzYfHmqmzAqCce9CQvPdFNNdbMmsHALMszQHcGMq+16zrqJtd1kRPbmAYYEEyNhdCBX
iqtAfayXy+aoTKFQJcaGia9ltQvOf0uBQN0TTadt/bZ9v9HKzcQsVBRXFrWRG58awdjswZ3vQuL2
5aH2CkWWJPpVzy311nXwEWpBHgVb5cLCDe7VIb3jxJ0GadPPlM6gwzkGYdNOaQS2c4ciBNeYO85x
iVbIR+F12dpmgGqYeyTxf3gLuE7iuQO2cpnmPlWxAIgXdNIBKb6eZJNRff1Sz4JyESQDiYHDuU5N
bSsst3/QEAY5LbZf6GUfOU5dUBhx9ErMjx9EUmDKdRsP45RY6+S9gLznncvo4kdm1L0xhgvuvBKc
9zJW9SNFF1ZbPVphnQVvuWEj/96XfGqwtsD8e1tD7q+K/JgiVhEHsVzmUIcigXBadsw70EVxLd4W
+Jff2S2jtp9dF+G8IxD2DVhyV0umTQ4djDMCidUqKKAELCGyklXVwg7GWGM0nND0IKR2Hc2w5V47
5HSUonLSp/62d6/8THarst3j5awllNpU+uEkG6JDs7jWhdjCR3h9AwgktqkFbu5HZiHtH0tyzIBA
8Z6GcnmhEvTtU3/vqcHOWVCxAVPnPG5CWASbztqlFnVoN7Er7Bb44Lxd3CgM1r6sRGCs1Gc4FQ4e
rUS9F5m4qefhtd3Kb4DmZHQjMRlWhc3dQe3vhoWHXvHMZ58oG5rja1Un5PfBqYfQYBpCMMuBvKms
3O9Yu9Q5Hcbqe0VI6L97IEnq2O6E+Lfdr9k5xrHpls90nH0NQp6GikV/e8cisQb/GxR9WcdBamrL
TgRtwJsy98wXVr4GCpJ++01/MFaFcbZg8FKsgnOIglP5InUVick6kzKIN+F/1QmptLa5/qQgChYq
Pws3vCvhpuQHPSce4B+2XAQwSKfUxzOiHK5dBO5DrNszaJgj9bVQZxNMBe0YUT5uyO70naxdfqB4
nZ6KlM0rw6s+jN7ROYsALp648aTgydFvbjd3nZ0inu/xKGzBjQxpDlMaW+izuKqZzjGOu2vzCKwD
cEaPQBV7DaHFlSz+tIlRMYcmJiu8qwyqK+ItS77toH2FRMsIKHyPHfS8NGrfzN6CHEIqornr6Ktr
mm+6uQz+Xu7Hv0Zy//Vt4jcrAknTlVYcZgqEi9tCuIeM0pKw65tZ8eMyM5co1QnYkcIZncWBUVbb
Udax0w8MsINNrx752mpLySIEzfHR7yoIzczVqdKLszRpxZFjLYyG1ysD9Z9GA5bb/6A/kEWSGcL5
58YHKyRYaINa4rKG/8pu2T+992WGj+dN6ryMyuxZuhhEhTWvQHvXoC+L+JJ6IKTPNFxz5+K6xPEv
u6DZ/PkJx4w7aYUhzAuMVrf2KyRSWHn1RZHxftUUOFx+hmVTPgWaXhtPRMWUuaX0TYiOhPlN60bx
mLsmVlc2Bv31cw06Zw8ZQwtHDAIe8rmBmLQYVzXDxdie2aRSppm5pHkeVkzbsYX2k4ouJXd4NH0q
4fIKkwL629pafNAD9Tvoj9/2O8LoHEX/uTNdMuRsCt29ZgrUuuyBRkIGtLXsJpEKzmv5sPFFKq+x
Pl2sEGGE2qg/rJzDxozF/RxpZ9n9Dfe09IJRNg6+YNmvagzO5u33kZDvMsZoC2T5/avKYiVCbAHk
sQ/bVMeusEhGhA4H/rShDyVFYllslI8x1TUpu4ZoRv77rxg41Q6NJY+XfulS9u6+CpiNR0ubr8VE
2Mel6+Ahk5/uFc8E1x4n2qBsGNtIFMd7kuOeHwcgyfO+LNbn5wYgRQLKWwhRh95sDG+wsHZGJkU0
+CvVd451DauVrrX7dn8grS+WMmbQ9Lnc9jnqvmVhR1Me+TgKpDLjzMcLMMvW724aCzYXoveUC2E3
nbPkr9x6i1N/a3lHl6nT/m2axUjAkfzM8PCjn7VHrrcK8KCHYKvGC7KFAy9kgwM9pqcfy06jkMQH
sc9QlUxeG3ir4lWXXzhjnCYj1E0zMQ0LZWOhYV7uFrJRpT/2IjoBUY8W+0MESJORNIi7ax9ku1ib
y80ozU8WjSLQX0BIno0PS0d0s/vnnWfHBuwiRRs/bRSmGYz19le0s+qAiA/g/I1H1rkbEuo94d2u
sJ4kuagwOthp4sdskoZsvg3Iq2ew6DW+w65yX4H57W7ipwH6shC+Beu2inpkXbYEl1qtBS7Yca7I
8ERr5TNUvArJAi3xje12L7+a35eigI3U/guEBmUUIQHgdZcH8Dmh5A+vdamChv7E9o7+jFqf/c98
KNtlICy8xU1AbiG6IVHyP1CdtzmT9yiq1NrR1NifbFkBkoF6b1Uf89GYIG0SKR1dfvsdXLIaWpDg
/eqriYbezMpdZNngiVdb9bMSjf9ffqFBfOMbYBaijucd3K1t3oxGwa/lfKXMwW2FPs+1v9PFAeRg
Yo1CPKHDcAEiyO6fuG6r3BwzkR5WbTONPLpZ+YXCBof8ktJtPCOzBJC8SfSU1rjLtyPl91LLOnUt
aCEx5vMsqWHAuuJQ9l7X047lNGPWeHPz0ijb3S32uBJWYZmSn4vyZZdVuNUCTfD9B4ZpylZlf1NF
KODfcKm6Juhbx9rLps3Gcbu5CVPWwGG/PBEjSC9o54vVS70zQ70kyGol8BGzpXfEKa3aRCcWPwog
XGd34EbSe5+03VDrp+p6Lb0ArKBGYa2dBvxpsqGUTR3JNaUJslczkeAmgQqK5yzNt9eRy7R7uBD2
9EfP232LixG3ievo2Sk0MKdhrwf/VXpCoPeh2F48ip/5sFcpJ9WdR3KISHWAU5RVLEwI2fbJKmuE
ezPA207SNsfNZm1D+Rg3XPtAmzOgsVCprXU3ChoSzRFj7/ZyFdYc1+xn7sQddb2xp/i8YvVjhVpF
F4ZTCYr2qI6roOZxEwaZTzZLKCBF4gbsa+8G/P2/IPMAzWgHOO8zxsSB5Imiq6orLMZvTKvWQ9P0
49ka/ty6SeLz6hv1kmbCE9TQYd2+4jS1JPIfctEolWSI+T9ymygOxWu3vY9MXdCI4HHR5AzlNv4N
6kuRkqYCPvWX/s/NHIB8o5+v4EQ9LZ3u89TUkfYoDoO8kjzoA8wQii9FvhiBpZ9hPDLEMh/mpby8
RA5SqmE/Jo1PMNNtqLU6pHaxy9Eo/USa1G10R4viqfX4xh6QFg5SUPENvQOq0z5/GexC7yz7AGg0
cbuZY4JqlffMBJDUaVpnnwj+PLYMWjwQzZXlPHAqW/0cjOPgaa83wRQOTnP+1/f+wuTdBHnQ+Czg
Qy/fAE2YOSG4trEzlqVsUaUNx3gcf/vB+p3qfD/ETgpuSUro+lGrMiKycH/2gBan1hldUCu4TnVi
wdCi3SrtWwpvTPdv8J0r3Ygsrw3cBizqCbiFubXEs40qdyPZfhRgiVg5wbKaay2Mr79VIEbpkRuZ
6mU1rTpDLEm2CY9vC9DWPv/dgaAmzIb6vJ4Xrn4oGU+NGTHST0G+guhznqb3uAW9p1KpZ7tup+qb
j+5j3kMhm7VQxJFWxPnRMeSzwkA6C9he5GMZ+WZlKwLaatULZxV2WQgT698sZtG2XIK74FKgbmDn
6kdDs2VAtH+P/Tnw73+fJ6luJ1YGDcTlKbyv5Mu4fRXJXQ2ELrYi/W6LtN0j55Xj1HTNZWaQLaLX
dERe9AItj6s2XJ2J+Y2cJsyGgafVaDR02L9vPYv5lSyLMd9JpjEg0pP1wSwPj2laU39GPiDjXFd4
E1U6umXCEkHcOpS57C/xogAEK+GovKsWW/CPigKSafXSKX0ynUqmSsDucBUEqMiya3KdncShWOnv
0jsRwkJulp6DXsNPHVyMaXLlNy+3bJg0OXJ1pu6JmMYscpl0IGbFxkZV1/phBjLKLzm8QeCHbUWk
2/flpgshqonocpkkTQTgJQX/x6yK7K9sElGZXEcbbTQwzAGTsmpt8Eg4rYjCI6qzYu+Z3c7o8fNA
lCD4qIGFJLMfwLw3vFE7m3f05/gxIsOFa2E2cT776n95mCmHm7/pPRJ9YcX41PMwKmOe7EDHCHs5
kKpLr/ZZN+4KYSKcO4smvJVvOn2azVFbNDAEbzWfgi2LQDlsQmrmbohpqG4wnaWxU/y9jpg5qGc9
cMMzrJtgMjel7Atj5cnhhMU+rfh2+HcR1Ps1kB2QXRBgS7OmHM+hvgmnVEbzgZWSaT447XR0VtQD
A8Ee++QN7avPGQVwXqq2Eut/ykCC14wYj3vQdPPEK0cmUrwESkKJzAFpyBHwwC1yc99NAk1S0XIB
oEv1CSSjStp1PIv5QYL6vbDQ1nERZdOyXiURLYLJwmKr4j4MjtzFri5ljpOjVQnOrYG+mzIm7Rt9
TrDzGRiNAB8WSMHiJ06hRUI1xQddroncTEteekxQaFXTS0U9ZGx7p5HAPNQ3xKzq9xdd2co1tcG+
tde2bS1DkDa7L6gNY18jEjQeHGwd2YvpUp3GdsegNb6z/kDFR4M57XAtW8LHAPqpmpfMDpjDTBUk
NzQqtv57zX9wbRZCWRj/jeUM42+qW58Ogz80u1yHMFKvuDU5fCZ361Xwt4DLcUToSdWeaOyrolPQ
9Ra0VsjXaaQ5LefI78QMNobbKVoNsv0h++7yjZnZg4gp8BvbYHRL4LP1RdVIcaDrMTvmZBCU9EBY
k+x8kJeenmqnXUONZHq06kRc85IU+IycW8LlpIz17Sp+kGMOV9RwdpTdKtHAee5jeBuabwwG04yo
H0FnngZi9bwKr8Z5P4OVgQD0oSkbzzaqQmNDmBxpvWXV7eRWEfa03uSLwoWeKmOKfR8OxAkVjKf7
PV/8i/jTGE80juWI9RBXX2MzTi6RAi6pszmhpm64Usz44nd3LJIlY2xMpQNUsqBKIjyV/66g17X6
2LGtZ5FzaQB+MqgtvoIs8ig3KrVutlJRNFWjxvZw+HaJ7Tn8feLNFR6WjowzYl8jNCWOE82gnh8Q
JoScKNigEGiDyOiu0uDwgpL8PfGT5v16QRoQap9nsYB/ZyHITEDnLv+KWqRY5x8D2XN6bYnXMiz+
xFzM7yXIY7urSQaJk/isJ5QFWAeLq1rp4BxVsttYXIB51C0oHQ67sNFmSpkUGaZlcNQMI7Sa7/67
GoivXjrUSCDMsgeDV6SpTpk2MAndMjjAI0CnEBtkaWMJd+/8lxLdH5kMJDeCtwcyFCnmJwv+QAxs
dw0AROqFy/5Xw1Ohpc1Yzk86jjPXQzWLXaXzIFNP0/0KSCpDN47tVl536p21JkuclCutvl49edSm
BgjQ9PiRv0tCwCVFoxgJlGyINowcXeqgWL4e7iwXbMC5VqQfMNn5vIy3Bl+T8l69PGVWWUYDhfkD
5bTS4CfEygaKm/ztioyebUe8yCbYAF48bgE8e8b8zgqXLbGdXCzYdfN7xV/VvvsrGigWJkf0+P5G
8SGBzeRR9IKm+ZUZcPIUMbeJDtq+f6UWcvwtBPhURrlQxLN+oIZ8n6U1w3UY8dDTeQLXi2Jqtuw9
3zSFrMp3CBYlKwSLawmukVhYzSE/Ks6covaKGmIeJbOKUY2sYOZ9Y3AOQJN4jgHLpqtOIiVaMWa3
49jhOfTvLSu4U0V3Ak63tc1giWXR982p5WRiNOvkkU3FcHvu5BPNNUzD1AUjzybVUt4zgMSKR5u5
r+e5VDfHFVp9cSVByJWMioYrMzy46nxsSL8jmDUHT6O/pi47uH/VITZvBivX+ruQfz1mp99K/FFx
cj7L2pvGlNCptpss3aNf8BDgw4r07Tksq8xhiYHZy/iYSLuG9B6A1LPCpcL6Cl09mFTwzt6xVNY7
KG//hF++gJfOKU59xUepGFVvQ3HmAr0CGeLe8/pdyV4aaQuA8lYIzpQ8VwTsZjbjbO5ZXzGOEfiC
KNJ/t+eKP4JjCRWE+QWY4FgsmM9w71WAaI2BOpsCzunvZ8rzY2IhegW98BV0Dz7G36oMfzt9A8cF
ZpaEQM28rT5MPes+puvLXpCcNhoqNRHmq/qENf6ZPQR91ZDOoXxjfu27JXasbfK5w87zzQSFqcbW
W+NibozDiBOAXzDDLF4B9xHubigSUBxc6OaV+j+2EPWhai6GkyiEqqM7UVNfRF8MC3iMrKQYXyDI
kUHpkehCS+1rD4p4Pvzu5M2dD/g9EcTeOe4w9E0NqRhG39wZlpQFi6uwmYP4CK5eW656R2BQ/o4C
ThBna087fmGQXdPfRmoBDDZLoOgdby9PDk1YT8JayF9s7TZOByTiL9DBbvbWLDYXC+J/5CyPQsZv
4/KILhD8LCsewnU98hMfP/Jn5hNjleSD/CYixpYNuddcGIen08xuicOcGA+I9x9XVYhMoGNvta8J
SFotXIGrqsyC7WYKzfjc2F5x2ddxi08KO/xZ4GAwPAkqoYBCMa+Vh04ZJTK8dcYVOkNkhptDl+n/
K7Wf8Rs7ibyGJ4lY9UqnJ3c7X7ghC+cyaIATYeJQFuEmGS09ffRvM48Dfz0YsR0+ytvDeJmxn0GP
6D/qjnz6KAYzSysBJTFBY12dV9BZ4wtDLed78Fa0L8WZC6s13Jy8PQ2cfz4E9zl/1hb2DGRWsARM
V4FnD6am2Q6ibMBSueXwUguGpClGgr7Hw7lQO22ZXT3SMblWOpbHBOmcMl1L9FDawkH5tkCZLHPa
TTWyTGEA4C5cs0cvxtQRWrSfWPC1U7WHyyemTPU5BbW6vqnO9c4jIftuYk4fWVyYr+A96ez/K1nm
Z21waPatmaqPaa8x4V3OhFPDXV1OuHsV3K8RBqoO+tlck/aJiLpUEo9lVoElfQFGQo7sfue7B5YF
CgI5QE+hRaETUh86CFhqA4Z4BF3nbQkWQ+rAGIZfg2eZz84KH3qotlT3NAU0vyk8psNfNij8HbYl
aTEWRGJjM5cazWAOx8ebNt96uAnKj2cpF0GzkHeyoaxdnXCTKnuL10FPCTVm5LIeTDPK5lo6gnSC
TMZ4BKIAQMusltfXZwK69uC9P+4Mrs7cbWsmnWhLlMK1ZrJz39p66l4eSpYHwPzxQFOVUh4MNrBr
dTDVGjumVgZE9XjrYhrXspElU6VhFKVDLnVwMSl72er0CL2VntY5pHvNVWAtjZL/i56wpEqRt/V9
z3Vq+3uJeDQVGHnTxDnZ2C4Iqxi9c4c6gAwWtmHUExwbtFUL0BH/O7bAqqK3SpbAQIs0kU7Qa8Sq
/yGUzljwuKbP6bGDTeIo/LbbwBYci3l92aMwuI/c4r/nUQKN1k6c4HjnJOeAGVc5sd5lwVzTPCwg
dB+wGyDZ60fJa/S92xn05/BYGH4gjh7dsPjtfxRGjK2bI+YSGpxj45oJKdh4wI6ZTXB0wpOUrGnS
2VgaRpkw6+waS+wEn9JZDuzFzI89aMvXsC6NT2nXTRB8WMase6M188/BiT5NrOqsv+KSYHi/aQsT
ZLbuAA2Syxid0TgEB5D78XZJg2qQs2+yv3MqrfHeJouYvKXLHLNlv5cA5ljsv8IzM0aS/yXgbJ5x
EJXwiLNx+BtXXhtlpZK9oaifPxqQjjzBD+WxTrTMncpS3+jYkDiUg5HTW3keBBxaAz2O3NCa4kvl
Eussk2glUnlItV5i31DgoB1v97vW1a08obIYaXsa4I/0k/wlRKztBZWzR7ki1VimNDRsYwqxZNTI
Lgj1OEhqSzlXM5a8VH9jqVcBM2uO2Wy1HOENcQLQK5YPtOjkP0TC3p/3XM5NAATBxp6S24LB+53X
REYuLC7TVyy+apOWZZRuo/R6ANlOgww3wVrD52uLe9Fti2AP7TH/1XoeszxgFt7QbqAe4JzrfRJk
3R7/61IF6C0JuO38wGLqObn7onFK4IdKrgjETQCVmTJsw1jxLsjw3rFALoGfdmi53RrzAIhIjoN/
y9ToTbE0vs9dySx4zosO3l7YYWKiW0yMBLcwrz1AHC1FECsbIT8qbwTHOhMQo3tPYrNTWa7wDbyq
fs0zT0SL1Q0xnQNnWp+klcQbwgLrCtXzsxCXKPzGa2lqTJyLRY/uO1DBV/twNtk6iZvTHCx6fh0p
CZ4XOMlhzT820eT8C7tnrLQVoR/V/c2ZuA1+Dlyxv3/RakiW36DtKSY+GQGYxXMqy0I5do3Bmv1Z
p916FsK/vxi2amwROjaJhk2Im2ev8hcMJUvyLau/t2gb43QFiW+8/CxCvlgTUKTWAW/igrCP9XIZ
7YnF1tfQkSOfv+mnj16PEzo4QbP78a2ylyK9JlFLLEi64AvVcGqdVR2JUSbzKvs2xShKqI6vDiVM
KIxECKV0C+siynil49w+Ho7gMaQECRMf7zmLa0SpI1GAVzL+F/fQgdpKLeEnGH7YU1mwyZl21Sa4
rXLQJvRLfDHvkHqIkEmhI7hwJRLrbU4WULYWp28a+hsdcThfYPrxw2qGejvvg3GgE19Fd8WvMLLU
dRc3RSHQMqB1WqyFqSf4MA0KUNrvdqdigNb/7yQbSYqYXOgLpY8/GiutK1lsV/bbhEFgGiDF0ZsQ
aDv3Nx0Og4TlbQf9xFsfSoUb7YxCUjLcv7RJPzwfDQhw16itTCc0/L6YSVEEkfHbZKixtiQ+psOl
9PCNX+EvkpNWlFh7GgR7tVI8kkNoWJL/aiAORVWO8h/Qac2gx5t0gtY7IhLFQV6BmBwPB49mN0Ch
IoZI55Tkif0n1vHxG3qL/DKS7mww+WdXcIC7IivB9WEuRgXINJAQUGlD7ZXZdpOy9CoDVsT6Wd7/
dPjwoRpQ37ndhigplvmkBEUVJqpKtzMC4DGm4vdnTh6HdQ2nchHRbj7wmJFSchMwqWNE5vTWl+j5
nyoDM1WBVF6RJ4TCTyTKbAjP0/d3nrF+K998knTX3CkbtcDIYtXU5tBl6dftngLFn3AI84w7LiyN
wUhVW0KEftV+y8uvf6cKVE5eivC39d+ZXUxJN70ZjKGKP+5ok0NqfDYpEGBd4zlW5sdPRaV54qZf
qw7tyrzVrWlLEWtSD/tSqhE+bibkf23+YOYFf3c4IslmOs9+dhxObOGG578+qjZkwa0bjeRLqeph
UIPH2CVcGv7s5BFSwdvubcF5H6N+ATbwePFru0NL7BfdxHwDZvgGTaOtmwVJzbiF6pVtOuCihpgp
eTjbfAhqWh09m/evtenxAim+QmRUk0nLQqE9RBNCaHYxewCa62qPH7uq/3AsPae2s67z6kXFIFOe
Qi7F8xwBA/PyR4cXyugKwZvRIN+Cfq5IepyZVfm323WdGwl44IMUr7/LsmXfyVQN+77MoRu6Ch9P
oxYItT04aFpIpzm1mBDMciYaIoOx19XsR73rlRpwLhOx1ISh6fa9yCJI3f0lsrIC8RpEX3G1U3zu
tVxykv+pxugTM08LgG/3zSzizPhNrZo9pC85/SYJYnh2r27xCNuwXlc3igjfuv+bCa/okO7+6sdr
8DE2+WLXxT5mWt9pf5qyyQNYzZmZ8SWtcRKEkSgX9WciBHQKwB1UblJpzhyOMQw0ej4P93YSZ8N/
FnVa1rtghnJzylx+285bu2tOk9ZWoiMuV4iUB/+pyYKY6MW8Mn1rmuGjjD/JLrx536t7ISaDVcnH
5ZkCY/oZjNWssM0a8LXaxQ1z0aaQpYwVoN89g3RzjuK9r3ns2qMd5PylJMeh6mOPLZWRDXwa4xdN
me6o5Lcbo+D0z5yJtdCaU+lMR7VqlNd5kkBhSWrKOSAq1GYrj2c2L9JAKfl8E0I57t2yMrhnyCyG
7XTPj8pqHtXWrc4Qs1IZE6NSNztq6LsXhDsHzmXmZ2n22XxBweTMkr7rcorsDw0Gqt1lOsGJ1Wce
ZdmAyUCiO9P0j03uu0tzQ1acB5OpygLhqaxDy3KqiclrmPsaNEsfijhNutGmQac8BzUNGkfbvAZr
6Yau2R3UE9Fdl4laRgZewscTERdo+1wSVR4z9NDVi1gQ5C30cOdce4iaxsewTfAuC7zq6zNdItdD
YWzxwcjwZhWntmk7NKI2Xn0Bxt9T2L1QSLzH9m9sserswaIb5WUIrF5h3Wc73zFa/cSO4BkUoAsj
Pf3iduBoJ/gESEZfp8koKLNBNUE2S125sDCsv6rBZA9GNYxfaz3XtpEqdcXPxjCLqQ8cRyKILuh0
dSB9gRtPmPYpY5VNcdDdAYa2l8K2DKvnG2JjmsXEOuQmZ+yen2B2n+g3k6XFBNILVbtmhJngL6tt
02+/+f8soAEcVPEcSUBRazIInlgoW822NuFNVuxlnkcfWWQK/d9AEY3OFG7p7qdczLucIlQzYALm
WzK9rqkiwpSk+kB984idFkHJvAkOwKtfTS/M7XcmvjVhoruBRtz/PaxSG282XRPIb8quSVrw76s4
dVHhT0eVA/yzmyDez9lhE0VnEqPwCCoekEIfKLKGFPRwASdqM5tRSokQTJbeX1pRKREQheTmue6R
Y0ULWYyVf2xnqLqX4bXly7YbJ+cmva227VTPkwpWpCejfro2TpBS25aG9ht55b8HvgcFEwCCQIGX
mdEuEjPQ9qvgJVVCdXAXQ+OtWY3vl9Rc2qSDfZFfu42D/k0gOJCCsWv5r6yI8VqZMfKwOaDhn2Yp
fJBFncZGLUkLqr8mboDRCxt/PkramncmKnFRuDU/c+t58RjD3Q4rTqcklLhuYwSnRbcb3QRlfBSH
drz8NEt01yeVV+6NTz3+MNMBw9qKVFJiMJDVY8pni74JGbIHo3KFvaOiEvmpBHcZaPetUZlnR6SP
bnPJ5k/6NSKiy8xiaYmmWBuvuPLGJm2RFTNNpDoWu/+fRb1ztGmYPr2QX4qIYKkrdBnKlw0K2P9b
1MRf3NEFhPvFAL2G4ua2+aQfDOJS0KyJiROhiLAHsSjivnGikcvGHMqsbzeAJE5xmYJisvczfR72
3GFlxI/ZiJooKk184CZAQP4MK/mojkiz1SnhcdSma69o/qrdlnzIPQFVQNamSJKpzaKiT0XB+oY/
N3PZvqjYdLMJtk2B51aFpV/bq+bxr2ftQOzEoIv6BMqzNxWuXP1jYhOuFq+9AyVXps1cKwR9wfca
YBeCfc0yT+IhhB6XmynCbMkSHpAREbRY42ASDk1Wxp5RNPjgWxdxAiuUHiOhB9HdBVKMnZ/8sbt2
LJUka7qKfkK95me97Oe1z9rWFNEA+6Y5VnaVNB8ZBRcOqkyBgUOzlMnGIsjvuOn/0h5nE/byMdxr
TaPccVlvuN07jDV0JFrrFNCjPXNswHWehdHfEQNM/Gbo/kZ9aSPANo6Geb1JdPOBhwyUzOUmjhSc
EKdJXTx4ANV//JCIaVZq30YS3IPvvaoYAWfATzpkxaI39yOMFDjU9ldmp06pdTCMhU41zjUxZVOl
dOFyB8I7dJ1eaogvDAVKQXVcGFGAqbD85VRz4WEgLk8zqyqWf8UNS5A5vrnd7QwjYDqDBAQKpM+C
Lgurg2m8RsaOxYsjbVcnblcAzsO8bvgDQhXx0WhEdGhFNKkYz4H9Q8te0lH0e4ClRcOyauzEuonX
xrI3Lb5on5F47zCsQh4p59+/nv0Ys49CggH5RzssXp0OWw6kWeO6jsHZ7YyHZ32Wxt/W2SfSCCn1
CGwZ8mlexaPWhlQrFyg/YwS+CK0ufpM/rLSVYb/aI7TsGWXQ7IhEquUp5Ut4D4D/TdkfVXwl+5v9
NdGGBkD4x9zafTeRCHTKvW+jX9BO+Wbr8NyLkAhkf6ieifGEI70mwPnMcB9tG8pXCG8Q1jDlbP/z
iQ3/9kCyLeT1easXKC3xnLJjUVKaF+7UQTVLD7JhmdBqgESbE8Ji+sd07ZdyCSLg0fbbU4HI6s79
biSA8srhZ1YPy55XmWG27awf6gR/QHTTXgthMvb8hhyVDzBmJMxJ+XVlXt2r+4Tb8OCglOPs4+q/
psIldHlZPOQ7nh52JPP/HVtzsDH3YRJXnjUzUKvZ4m/tPVSdk5Ib0fdkg/ruvx1BzQM9eY7uS/Cc
w+PHu4jHHAz5SuVKXy8zJGUFy8+JJtSAcA7XUmC3GrsdrumibzKzpIJTJtnGgeUrDgur4+h7GzGl
rkkcEnBjLOq5oQLcsPQ2VfM68xqufj8qvLdcm9rWstcyw4ro4ZxLb3EUttdF7Bl7VWD2GTunBzUa
/hf2aHF2/JhlwujpiTGd74Pqa0fcX1SHfLpNyv9XFU/Xi63jm2OTX1uShA3/k3p/rhc3zwgO00yC
bxQ1XUy+tue3pYYbco0nSqKvxxLnIdZV18LZPUiHMBwFNIlzwk+azcR2VXq7nZtzzKNRDMK1VKF1
neaxlSFjxQYyJShpCH/yGslb9eTrFUAbvxAF1rCBq9lJ/bJBsURFas655r+2YtbUWHI0oLK/DOX3
7XetJ7CtwJ9Dzad9R7NXfgrmzNjw5ai/QjDucfyMEZYfyIU31sb+BsX59C1vHA9M9j8qyvOlhmgl
ymsKX7hQ7hFfj2YXMkXVZXY4xt9YY5bzwk/4CZliitmPgzcLv3kSwnpzMCfRzEb9sA+PNIgtHJwZ
OIABBrfVVnYed322qW1DWV5CY57Un+DFMD50Iak9/Fz0WkjSX2br0je8xXEQF8YzfM9fhiXZYocn
1n8DdSK71IE8DlbF368a72rwFK2Ts55PTM0t7+HXnseCjB9v+1rX+4QPWaA7mSP2tXkgZOBREDHu
0ymtLv54nUc2cMI9ZYytXJq+VbZWKhLeZG867dCn3Umq1kdOgr/MS4lns/AnLJ+98N7CcaP1Nqr2
jYa07AKlzntybnUC+qhXmOnilYqkCzyJWF8LIXJgwOVQ7YWj0rnSOgpujj+idsg6MJEp3FnuBQC5
ImhHYlXtbBq01Sx2TuWA+nyEgqij7dvPMx7AMy/XO+0lKGjrZjZ2ue89uGfxheuZ1FWd2uYlchQu
JRO3WY9SY90kblOlI7dwFFBKB4wlEIVSAK28bAAyljb9qkwSYy1NPbeS63xgrZz/nz7VyBo/xwXe
QMpWzLhSJCUXX/vt2LQEocMTARlourVlzfCjZKxJS5NUyKy8UQ20UvGsZHr7Sl77hN7YLfyHpsY8
YtWRBvc3xHJZ8jyhv3cl5pLI8i75m+zvkezAQ2Db7fqYRL7cCdG+9pwKIQsd5f3A+G5AJWa36JTl
J0ZfW9oQCPNu79Ecr+iiBo0Q9TFpAALTQ2J4uFWGIGm3ynBApR2E0x8oElgxUvo+TQ2UGx0lMJXC
dZ0DfXYa5PCAZwd6S5S3CPQ+T8XJy4dMSQwlsvh7plsDO4HVEUrHBcphXyHWdzBSgC8AeRVs3ucV
oOf7sW53r3CdnyAin+8ZJnrhE3h3eCt5Z59KgoJXlQhVpjznGzsqpE2QdkycEJ8EIEOcpqpUYVZM
lPSOsnP+D5FigiPnBVZySt4PdyZTkT1uvIdiIqgnt0zYprUZrqooZk92m/4lhFCDsbNLoXeOGhkz
3fIsxtsIAatzJHI4KRCyHH4TOGnD2L0c0Pq7AIu1W45L7d17WV/vUOrHRXyiu1iEwA/OHxqG+CLd
wJnZJdJ+zq0YPKotCeB7vrBSu9WMlUGIWcWVvwEGihxDJN6zUxfqGZTpW5IZBgJOg/1Y9S58zgj3
0WkH/edIkbdTyjQQ/7pwIkClNrrNzwn1udvGigNFmYDzKHCY08tM75rkUCTHIjeNaCBeSX2x1OcQ
OGZLioEKuiqbi5U9tB1SOb0mxvr+dQjRYkU/UDoUm/Pocv5Qap96fHziUuGSQ7fXAALOvVmZz6x2
iv/FCJQcGMCACy1Oc/Aytq861RZSO8GZQbsiSiMps54NQpgD07aA4Gch5QgMheDXUv3HgCxLR55u
vIj+zC3DBy1sZOfsdpzTSX9+fA1s2+smil3bxlNENZB+S17i29B46jPRZYzhVjn6GisnIht5RtKI
1ublAJVwo9F90kU0OYN87mJsq1l7Is7yyxABLNLvRzrcDcRFILORzPszDGKbfjbpBBUMp3QJAauL
ZZ31p1ab0hMu15JvFT3ZU72xBd/oNMxmTw60Z+7iHVrgWY97+wFiq9amdKBGIKwyv9fvIpPnYmk3
WOla8RJSh97NXV9it3VZtEeGRmQGGEd7z5UPMn20+q57YBZVdPkBGCi/KOrJt92f5Ukz/flO5Vwv
9lSy6H/OErzIG2/KgkpqMF1+fGl00rvLFEp9M8Vyrgd0XZGzuNf4IhhdR/vxs2Gas3voq+9j3sdD
UZM6nDFFEmlyPcPB/SG0Ko3QRxFVUm64fsge3x+ETZamQdf3HKZrnxoppKuvgNasGIi/MSBRAqvi
ZwclFpyNToYXOeKJP48uUAZ+SnV5f2xSY8eqA+sdUrbP+2l0BBLRbSJUqj7U53rmO006s4UqEtAj
atPh6Cww6pxeVdddyeTcNfyCWsfo8m93U7drw37z/s0XCINj438HmEz1VwwrZhnSMZgOQ4AZDuUC
TnxEcXRRt3a8b2sROe+gd9xM4jOHspWmAVcQlkJxxf8+l6WXNAg+eF2jwnflTkAb/QCuKZz2z0nB
e3JfchWOA+HdBAZ/eVLBUjnUUDANTQOItFqpmxMTb73DPpcbagy1+4zfx0zvQEVZc1kYH9ZeasoP
AcDu8Aygxh8A7jXXPUKBSiEox9hAVMrgHHrJvbGikeQVFYWUx6hrg8eNu40wmES5BxA1Wpf6p5Mx
goC6L8PdAEvjRbsoEfvBav96p7AyRqkXp5YghrKFUhiZqvxjW/mYbYjUgY5/bdrptBbDZfLCwVPP
qcEd0vmIZrIQxYlNV4TQdqhBQxezC1D6S+M5RNJChpMqtHKdMe+OiRlH22KAVQVwK7vq0TPI8T2b
uydAryv5CFqgCyBCTsrKJBgogbl6d3sJ68eX9BgIVS0dEQjsLRw8w0sz+yqo/Hqr8aKeIoooYHqO
VkVyLU3jUFVOcdjPZIu2FCQ+TM6wAgyzj7ebPjbKJU6T4fGnpvu9KSncPEd0Z3yG6m9WLDwHyoDE
UJ8WgRpHCL/5RQoGE1A1l4/+AN2YDPEv4sRLoBVoaP5hHXYhxa43T6nycQLQDH2r+k6JRQvNKitg
2fNTZzhCKCVqvCgYDPixgaJeVBjU6Bh6seC8jpv+s+Erq197fusHlzAM16H8xK4u1ZlL5WGExoW3
GPJQ4/Y0GG/EooUWrBWAHtkDkPZ7X3y2Y3ZUzwZbCyHRxToZGKYMcnt+XmOoqelnEW70UYErU+zQ
Hc+YMrro76DYYm1IUpGvT6Kxb5F7RS06DDxt6v3Bs8Rd7Mq5JL94jiuW38h6yYRXn/LQquu3Y2LQ
uKO+rnjLhl/8d0KYgvRp+AQBIvZtkeDtFpSD1VT20CmYmKWFsY0JxZGi/glwE9hGEfn4plXwpQB/
nT4u4cGYpZFr92qEd36ESiZATimd90Gxxu7TvkfE80ZK7xYBQxUzyHiy7EZ7FAr26sFpFxAhgbNJ
TMPYTnf1koxe/uGEbqVfBlaz+E41KijzNMjs1nJLNE5EVoh35+sGCAjLLHiP24+FX+EeyZYsjV9z
5f7Cxk1apry3jnNWQ2Cn4FQR639+Ucvl/uFjVoC9/LOeIh/BEYXLRzT/KvM88xRMKClzTUmvDbnz
3PSLygIVB5kcUQanQr5m2zRdt0IiDJzE2XwJbqkehheobI7294pD8NFGi22j4BoQ8ibLhctlGqGk
NpLDidfCb19ExU9Ab05GXrxUvVUQ7Bq8refq33ecLbCpWuObzfXubzFFcnVogzVlIZFS86zIkkWq
jrfmiax0dpl/Jvd35cA7mepwSJa5ukaLw0a7SBJ0jfdhirvAYYOJtHZzTzxzkMTVzRxqCq5yoAHs
MDilqyHho8ohWH6z2CpI+mfWOhq5UsDPUMX8fx75uKMRaNwva+okW6Gv5OP8gxbRt/7BnNq9fUWj
vHtfBhQ6mmMflS71VOYKuN6xLW02YBKSwgH18DLzzytlgQ7Gbcm7rI9sBxaus7BAmsCV1D14+l+v
49qKq0Z63X7s4cmByxESxN7gekJabVL3IQBcTs94AsgfwApGveEe/3DHJNuXtJVkeL/EHTArZMys
/ryilm3rQhTgrvIvfXx5hqCDIXRwRkoB+YsKmNSwfbz6h1CNy7cskj/DxwI5XEIOdSiEyUodJ9Or
rZL3sJchWOa31Zyz+yk62ozwHAoNsCNkzfa+/iyvNl/yQFhtwA/qIX9zQyWp0J77/4b9BEhD9ABR
anYRmFot0wBCVksh3QmRksxb5Fhy4439a5zIv3cz344lJw2SKPa9Us/1DLQJs6+aSBC9cXuHeD2Y
PuHSsEqMZPkbuesOnFUn70k5d6RcNV+TLfNm9RmmUd5Kb2csi2YjUsI5mZGW/fECUV6cuwZ4Mhfs
k9yfR1j0WVj9WpvPcWyx6mRfaByNCJZXZjdKz75vQto3xbNU7c/T14aKypIhmiqdvSqyOeUGKTkL
WKYbGZPbyaB1sr1RgbLXuojgZf6cTdBMaQ80771pWDkCkK4s1OXqStmmm91ftdgBLL50YQC9xhKU
u5UuTXlli3swE96+lAXRkeD5Tlr7FVZPHnPCyJbKCpHEq6//LLy761HmE/IzjZJkUlwIgZvDKKpZ
5iQwQx2eQCm+xY0oQ6w9aCkMcCqOYTVitUCNLAdAuFXPYd2G6kxt+q+1zeNSi4/ZwCgWXgWDpnNg
+7q54/k4tZX0RG1yqSSp9FffRUVhHEMPEYTGP+GQ0Aa3+e0sPAuU0wFiVkhbkUT7zw9+pFLBBft6
ry1Ee7sDUoxFPze6XLZA60lP8WgCWrMsVcdgrsD+yHHrxKgFzBPNr3EusNia+RirjtlelsxI7Ny6
JsLFl6igBOQNdEelf5S6tv65RpCcuXLr+K4CGRLKKBqz+DI2hhSdzL/zUjE8biLxuKFJBWl3QcN6
hu9atFa5WgxV1gyNZgflHYHr46Fk9mVqPh7bF7nUoBPd2SGcmdqJ6Nsi73Ivhds8QKD48Ylehbw2
DHS1FDlJmjbtRLbw6KJlSvpjNDQRVAj+vu78zFm+Lb0DBAiRwPKi+wAOiFmd7eqhStU7sWhTNvuP
P/sXqPBAFIrdBlvBP0JQ4ypxIqeS+CPXPTcpx/euH9VyIc6OeVtV3WkOUw1RD4jXhkNX4+ypYDry
p1tbcG5oPJ68WXMITA0U/xwSw2MKsO45XMpUPUGBG513HptUZScz+dKlPBD8X1Q9k97/AnjPImRJ
ZEqSKv42SZXruzfS8gWGK1WhRU0BM9AfnQ3ywidEy0cF7LAC9gOqjrkPftk0ALxI6E2zLD+K8Uwm
CNzgXN+jgEZYDQKfxPPPyHjjf/K0VUDcm8YTq5aMz34LC4gwuAxv9ZoLy9f6X4hvN1vO3FV6vvns
ocIWMKI86fCjH7ssZjfYfCQ5DKA498zrxvTvzuJfccTn5s/UG5YA21pU7+Zd+5qUk0PpuqQBrsXY
68aTOqfp6MrzqeAD793tWm9ya//C4r0Ka3IBVHT42iERiEYNaXlFf2uPZVQTQtvxDiDpKM6iA63w
vmfPSZ/k58lNju8htwwfjoMcYmDctDWn+tQiIrYQiJcWFYuiQmxeZBe9QzJvDwK63+FnWN3EnuH9
YF966bX+oVgMjodlFcfYolY2yB0gWm9o6vAGAOglspep0O8z2Y5AZTyxmsFCa+gXJcDW3Xjxvpqx
PS2GL4hhD3MOnXuFQ0Oiy4rWpdSuAl79PeOa7BdVMQQcFqBLhT3x7MFrbQ62HrjN16+42+p6dN7O
iq1Qpy/Gi9ngNJGWb8PNMfmUCeS4KiJBFgc56ZKD6WbKor0tu+u8uMszUqtd5Stz2VWV2jZJ6pO3
P697VvJD6ohI7NUWaDw3pSlDxNqVQLMnFd+qzX8cIdFPxXeIWXJCDteR8oawBkYlHruCTFC8GmHV
qx6uOJrHb1xxeHSrPYZz0SrVddA2qV8xz8UO8bEz8d8jxoG4pn2+7k1Y3aclHoczs5ZuSj9UnP9o
7HQoxhFRdnarSlYMpQSqtqfZ55D4jN8bBri1Op/PmbfIddx6EcMDPeJZ1ftmuVHbLyEbyWBQntm3
zmu41zMI6bK5Vg4vinyskGKEUqzx459xAG8Q8y40wBJpgs8MuORKDghMZV6OL8bGNyiKS/pFVgVB
1yEdt1F3qTJwkM2FyA2pGjasyDxrUWn5Bzxg06s6y9ubsEcH5RmA7pjm9RPYipox4mf6Hol1zNO9
sp4IhhZyagnh92lQnPH4R/p9nk/En2ygDKaQWc+aRt/c76x8WmdhIyjmDqmO7SLv7WBR6bolMRRp
omtgaFkqQ9edm/nDqbMzfXnZm2uj6FMNGDzfDo7HJjqsZcfQAN4E40pXr6AN7uyhcv94Z9tQ7ZLu
eTNr+nZBWimtdr14RgaGZXvdG1NbplR8EycZ6bIR8Raq7o3WzobOf9uu2GBAh1p3QPOHtgd1QQcy
nFBJifvystw12EUptuDG5bx05u95DLEcu4MxmWJvO4ugbKszCspF5WPBsHs7fgBEIVKI3H7I0HEA
gxLFzWkBGKN66b92ahW2eVhX5xRUynydXP5yJSleB+O6+rPXP0iWUJVpLNbwp9bvi3HLjANEZkka
WQV7owzTPFqenSsOH+3aMslIPkhMkNfG3wwkjjznbaN6W4JcLkMseQDr8ZRA8i4cM+5YfIdscq84
jmRd0cvhhEvhFhd42vpuKT2qhLHvDGJighDWsYGfKy1Ona8QR7bfkgKFCA5VKnmHG0uGp4fu/k/H
baEqJkT2YMts0+ZiWnlkYamEZxZXLDpx+OzEYhyqW4K9PIzDe5SkN6XbSQc6lUqcSHoR3nv1/h7B
NuDf2dhVtMCTRllQCE1v8yX7JkOfjyYYI6bqTHMleBiKGObRKUrL9Jyh4kdwIdX9xEmvpWQnrkZ8
4qBqN1rGYc6xsJWxqcR6Crp/gjIzWxctv/kdagdCaGvdBCDlhhw/DP2H60DYFi2EdZ8/BEpB0rUQ
8pmN90625ea5BJZu96OEM0uHcf74uvywgNmReCMpJq+CrwLhOydTEVkgp6lxNITzKS6laBmJ7KIC
zcYGw/KRtt6DDsqlZUkHD92jcFjEUu0Q2JXEbviYW3hFpQllNwUNr0JUgHRW9Bl6TT/4yYOLCkto
VF7eSkgLodfQhCmAjsWTXom3Jk4nx+1xGOptfa7/nf5GVqLB5UWRllIXI1dtu4V2HKVoKYmkw72A
c7XkfpMvRFzMZc7x6GRtwVOoNTWoWCUlsh1oatmx+wIOeoBgMR2m2iXPRrSevw/+khlVKwejiY9d
QeWyjAwh6N6Q449EJvt+UW5BHdFkHOvxggY/eR2eMA+oy7tpvu4norlXXnP092QBjtxkhB6UmhBt
0oWdUdcfbs22dpFm2iZ5WmvQIxjThUT3TUctpLBueX2gVUKvxLKGvDZp0a4jIZVLygXuzJBajNtU
uF0WeoVxrEqpQ1aHyyhjzeMDzVcdCO5GtXIEbfl8sgyfUGErBvs+gw8npgCj13E91C+yUth21riz
WZ8jj62pn5lajnJ5hOAdz1VLgxNTLRJY7V6VBhWFfGx3rGKcUe3uArYDdzgXgih6/xOq9VRiCW+L
p4H+/WoApspXsbt7veWPD8Uc6JPuuw+U0mcMuLmlv993ngO2eCH+MX/6rNvGM3hwL+6LwteEchng
C1QaxKELgvCQtXICpJ4y+2WbyzqnxjDt4AxUGYD+bcLfmj+X4XmH4m25guhi3FMKbp03PyY6a5uh
EcA1Wr21iKhvS18Y/J8SptWmnq7OfiNkhMDvIHERBEUdvgDCJgF4MzwHBRMCkzP6rJUDJUB9bRyQ
vlDZYVWlGhlu830iQJaJzGSupewdMIRYy4oTse2Ks9ytMqntx4jGtv4OtDN1cK86e/fUimNHLmYc
ulrBl/pFxwnE5Vmm/NenZLX3hTGwDDnLLNrXUYJtAFCbaNU7H+f7SJbTzBXJjjGeZ3ldq4z8b0Zq
VFS8y33zvXtdUHfii6nMJLZFE0loRVZUmGIDdzrU2JGWbhKsSzPXL38BkeCTrAKrRDB4EfQbTgy+
NZN3mr4sR6x1TAreNmtbdNzs5k4/atb+2giVhPA9AuhVOT7C3XQzheT8OSfeigpJmTZdBB9LQkbm
bjsf+yMUzHO3uTtKGiul34+DPd/vpbQqE+ufW7wFr8pxWuc6heHIqW5Wq59sqnivwnpYjBpELC7p
SpGMwaxMX47ASlmtomDztrgO+v82JLt9Xx3Zy92YlAhtCdR5UbHbYT5bfzvi6UfJUH1D3HuAxdzy
MYFMkCjHpn27WGFIyvlSasImHPyY/Tmasp/gGiwU5oN3IsakvXe6e+1pcDPw0guGfX5atRWYs72W
m3FDnMeORB1aQbGSmYboIQ50oCillk8iW01D80WSdEln9gs72MTBPKYP/wwbnsYtweVmf0+INpdW
Gmlmmz8A30bh0tonq++Y4Y32P6CIQv8iB9FP6Eu8E8KHsuyYJ1XTfCjnuficH7KRFWxmjTjE9tHa
RUaYmd8n3btKw1PiQSVXauJNi/C0ghQfWL+kGlpWMoAtKuBIvgXM8BtSd4h+SntxKH+ylO6IgW3m
Bj15KEg5oIU0w5N2q+vRnEJvNiA1n+IsFpz35nFNRWJC2b7xCSerRy7gO1E7aQhY5P2ihjby+3dC
uXbrnozImLwtXylSm/HCXiOJL68dcizJKYPkYvztL/oMPlfsgxFYjWUYMZZL/9f/LFCWTDT1HI8m
+GHW4/ArKauXqn2umE/i81ed8dT6LcD8VmsCNctIihYKc3vG3TaC4hm94oZ40C9nyQgqNcWfmauL
EkyT5Y6uBOTL5FIPGCNengiv+a/thFZBOhme//M1b3sLJwYhLxtq0gCKSfwSU6v9azeggTY8MFbX
Z9erycuTI8dlqvcY2h9CufcTMDfJvagyY4G9f9f6US6uHAiDq1JG0Ay2ptgwsahLPLAzpIbFjYNw
oZMywhu2D8sqfu8rXoKzQRcvIXo4b21pjrqcK9NCKjuYi6alLlo3ELm070UZCMyrAuuoaaCUaJvY
KH5NIH7cikcdR7MLnadPCwxqJ4Jg5vBbM3ahhiPTLd+NsDrBP+qLNXh28F5j1/cXFfll55wF85uN
kW8gGIwVfBaYZM4PT4ViQ+UY3pli5SwI8N2+UUX+tZjnkq/rTQkvU0z3U+uzqMZh44XeFbn/6kr8
85Tyheg6OO1jPNeXv5BJCnje4NBgSZpg//h0SPxtnAbBNQagx/F2t96oLDJ2W0Cth2P2YoZWVXCg
6D/QzZP629aut9na4JT6CWnsbg53XIGH2z+efoIlkulbhK9uKsvWZXCbRG6F96LvhNTuiKc9LuMF
ygGp/hNVLu/0az7eHn7JGvUTDoUnOwiVQp5OQOZPXnz3+k+XtYb3Y3O8gmuLaoGnidtIP3QJ/u8u
imVyu4apVLUriMzUHOzIKP4NOHZXJzg5sD+YhAMmEhvZvvDMnOYYUbdPn7bppyQ2e+4kh0MtZ0+F
CWyxk+Y0wBO8cRHWbxUBirMnetiYJmIofhdMfs17m9L3INauBJ9KVy1mpxhyPl/v1wLVLhyGO5eF
B+OMxpdrGbQTFkYIkUPP6p6L/tfk5/yf4YOqBd54fz15T9uzjhW+ocVjKbbgsL71Y/Q+GZhhJdwI
8T+daD+YR6eRtm7B2dq49J0imGWdFG5BkW0wkrPtolWDnOLMV8EsChiK59efKJs7gWjIdItQqNe3
mis45NPVcNa24udPLrkv1P2cRwQh9GrZy8wjf/oCgkTNC4z2sF39g+OHtllJeasTZDENQSXDxx3D
6Z1et83reyaaWgExTvYMkNEWCm1Pzyut13fT3QR8uDjtCmhYah0a+PZfjak++JDqwitbbf8Ny9TD
2sLYKpf8XIh4LRJS78uzyfPjiSUV42HVtjPcaCLoztk+uc2wDxhcWu/aJTGeCVUa00eE/VRnyBug
S4LBxvov2MPppzHRjuw1najWxvNtxnwWB7FPatUzX+b+LaZYKieTlLRj9WGtOCft8RijpBPPdoQD
mCd596MvjB37V5uTjRBi6bkoYB+QTH090/itU9kvtYBGI5ZXAhomNdeh3fuvGVskenfif0TnD9YX
iq7xxbNPUSnVyM0AMD3i26qdVvJKPYdXHVfD3fKQMGBr2+rE4lBTvTqjRbjdWbmClp4aQdI2B+tU
sVeP4mupVE52A1VccleHAZxZnkihDaPIQWwQGqs4Bs4y5m42lSEy277h6yn0PYkR9UD/NVurvoP9
bovoY9622bYiqFBMB9DW3JEk69eYgWawO6e+XQhRd9SoUkuDW1eSkGSDJzvKNSVdUWQE+RreOZ/O
f8pVJavRPKwGtRf0ElimaicomYbpK8caFF4bHhm+r36481aunIeiHxabSEiDtnSuAtz2B3zV2W5O
HEeshblYfSKn18yd8seka5S6+bSUB04O0obo1CLlDXocmxmZ2kgYp7930PcZCTb/UEaKKeqBmimj
DiO7kMBYDISVZcuVdu6OT3KN+WhyAr1OpHARzS3bbergfJzB+6Gwi7BaRkIVlgVN4o0S4NhByix2
W5uVXrExQETA15kIgWm6S7NSgIDAnKyjrbp7lgj/p8B1eB5EIO8ubWcaS5JQYEWHv+xL+R82t9Fl
LDPDScA2HKWz9qvj4LLdy3mIxcRV75sjicwRuDTiHjyy6YnH1b3ZSBGcsIn8Bq9kP33kF2klENmj
an16UZUAFYMXQUeY5cTzAJzOxGjOjxu5R3+XdlpC9Kok3AveF/fQKGodokTVgEQIsi62uofYC9uh
pVvCMHQLltReTiQTQFdNT3XmrmP+zCLtskHa48ia931VnFz7mkfuItagJ7o3QP+o2UjYVZSo2lZJ
FpsAGdsSItNyvnYKPOdQ/bH6/1T5eNPAQVylBKDQe53pb2CJ3CiR4dQIwE1Y05cwNk0xvUmPChmg
8igIee/rNTpVLRMOht5uGhXQQCcyJk8DBJ3khxiCMV0ZBRalESgwvxRdbQhGSx5t2ArKyui9+lwJ
WuNRcBT5ux+QHGeNcdA6ERfIG36/rb9qKnwLfsDLlxoE3tCyYZdU3+1kWnxyY1uTyHlShISmBtnM
YVI3buTFOvT00I+W0pbGIerrwPVRNRb5MvOKzK95Nm/Ifz1qcVtMyv+XCa+0dXN0oFPJHesJboSr
f3IatglUKQISjx8JYgvL8Q7v6Ue0dnUwu4QonHQf4BQJ2PVotXoxQLS4RkQLpO/d1CpprKv7bFjx
ix6x/DQ7FIOBvXG8z0H+sHlEA2hGVDbQbWeZQ7H9JQKlY6wpvYoIDR5fAQSU4MjEAwwaYZVCKfqu
M3NbSgzGhK9ttTRN9ddXRtsOIcLgfbVCsq0NSF0W5Cn4I9NIpFCJunAuatxLYWtCMdptzKXuDDRX
0kRZTUA6YzABEwmw4pPpbkGNauOF9NPlZWncz3v8EEsJtHisXkrJt6E0nDiNfKoikxKQ9ANoNJjh
1LvDZ2g82jARNPg5uyODvxjwYXmu+efbQcNSNqiQbRuCrQs155RyJRhHQE7k+ldS8rY3ALajCRBl
3rgBAFb60mApDcuLIuFNV+GjLA9W4oFMGv1bWSDyw+SGsls8h7jgnUdPAH4mDBYlcXM3or7o2MGs
GK9yX5O2L2yS5iWzcV3U4S7APGvHBWOVvnTfcC+wi4m18QrgBy0UJ/WcE9INGu7sP12UthRkbcCx
M+0JML3rAZFZ+F2ueB/jklqsewQFl8q8DYuhldhqL6VLomX4Ijax5hDciUVdKHqQIScFbxhnVTPR
9Ao1maFqwY0WT7NuvRQkfWlPvdY0S7mAW/xSLDbxH3RL5CePreGGCEWzOzHK4cD0qaRuuLTX/OmT
lMI/urg9nAAKYJA1hLRz0RtdzS7RZ52txQSxkEClEYYXyNNQkTVlKchguDKNBOPR6qzAuBIy96Ou
CMgwslHg1Jy082rcXCtbXJmFIyp2YZ6BCIb6pLzPM6VIGmapN8kpy5P/KKZxtomkJEWeRwlSMsNN
KxxuZC50wKLI++Ei8SKcES8b5Q4BSTtqtYjFpytRPSueloUaVLh1OhyMGUhn1eYU9JzRVA+CrjWB
WGrTp8FcuFMUmiKM/3XnqeGAA+bix9up11cXcNapAdycnDlqcJG9wM0ZRIOHTj2CIjVWzFoZJYZW
SH59d7RsY9TqymEghnRY0/ojEcaA3pgqFGFMkbWMyvpeGul10IW/sP34wI0XD7UB5L1AZixaov84
nrx5y90vhclzZnuhq/6XXIlZ9iiPn4PyjebQaZWAAGMxQBmCUwVEGufVD75DYTjnhJ9AJ+klycnS
nSWzBzONsrd+tVq0wYcb5XbOBeCo0aqWL0vPk7HWGEkGFQ2ev6t8HJAXFnnh/dTMK35XbGyLOQfQ
P5Zv4CNI179LwjW8cN3rMJlhYpo+bPoUKlQXn/yBklySfPoZjCS5EpGRces+POiE9eyDbbmfoo/9
vIFt8kxZdKcwq9GoF8IXJJBuXggK5LhaZd3QOWK+GnhmKhcc1iiIyBZ00kPCczPq/8Fa+du+3abK
pvlkm+MYKMBtY6nxjoAFnc6s/ub72qCYfnW+nrcXi1EqsSeUP9w+NQHI5eQBPrgar3LPiy9mYV4H
UDYUswMAfhiCFZK/J1Yhs56GSoWxLSTfjApUWCVtAGZfoalekZL9BHnVY9nKAqKMcGHBBqvWP17S
+/mTlZp8rMILhVg4MdsgXtNy8Vg7An49MZAluJJO3uNyMS5I7a9r7V6bYnVRJd9hw25nbNlEtbcn
oYAQQc639SbokTXikRJbm+5jwGN/TtBuYP3VSbOznQ1zYirRiQyc2hNJOhJa27ApNLP0J+jaJuTg
jE0picOuFNgLmLAFp57dExtcv4jkpe/B4EZJnNzMSqyfYEqTxMi4rSDJtv2ubaQMoDoDvCbNfJBx
hc1c968T/D9xg8yS/2wDLAbXhz8JPOofRrRB4FdF9D+YLvXQCu9Bc1HW8I7mF+ixJSdR/QEJydTA
/FzT5OdN0t5vjZpTdAfHZ4d3CqtyCJziENqjwfIJ1iyGyP9mmHTS5NEjiEot9AP8DlIsbGuXNMjp
eWUK6Jhdcr6TZCcCLz2aczIurl16RSU8xliEzZ3oFaIRuJDvQ26gbapPvJCPm4K9osgXsnbz54yn
pDZL5eWpFtNzM3CA/NSt6gPrYM740CpFadOiQKPVgmq3szBDqRWYA9Q1ggD4c1AuQJNZuKrSqeDU
xapyP2L/crl8GbT6KaMpygZybokiNRmpz2s7YAjPBIvIKjGaL6bHucV4AevsP6m8mcG+mw9Zr5ja
+ymvcGjxBm4/ua7+TLeudMaaJagg6WoATcSMBnPWO7B0pQf7toXmlUCvdC/lhqbn+QvGHULSwmo3
aWO6O9/U1beXU3XekjeIk4bfqeo+0CURD9zNcRqp+w90E+SkX7dIv7yJ0KI7wkDcRo1vY0se3I7o
f4YtnQz8Z9IpKj2S4o9YyZKLvmpFlfnUDQvd4ineRQ1e9rqU1PTKjd/fJMujIPMvsZMTfSXdyb7M
IRuAZIsz4GO7akVd9jbdbtti+2j05n8zsPmj0xviVbMeZwC4+jlbRW6nThYcaNYAldIfJQVhb16m
5Uh/PyO2d9bvoOLL8COZCtq+h7nx6Tll6MVe1eJV4WA9GZ7yhGeH4W36WGzSSEQT6l/PaB4NTVct
pQDXBes1lXcxjrXn4YCApgo6nabYSfroJtOXp303kq8bNi6Q1dk3NYZfcCmBXDEetKWU808Fy3Ss
0ZcyJpv+vxwgTh68BGHQ9wNIfP8iJRckM65wwGcg9rD3t3qkGWCWwJgZ1rONk2dpd62UrcPKFuXU
phVHsfSeg3PsX0vR5g+Uo4lhJBlL70X01C/zVF5UvfBDpsVAGMlDKhpXpEJoKOCvp66o8hk650LX
5LeZdJZSvhBSNvKk8uNAuTfdnauiZhp/NeEfknrHmfnpK6i8KTSgpkhEjdFdDLJPzVWUV5WeYszv
BlejjnO+BQPXMtHGg2wmR5m+3fRHdGNEPgz8wyPo12+jCmhRlEi0RWOGv3LkqyjsqKygHcecZhkH
3hfO2bUTfTM5AGTKITdSovadcGek+ZY0GHsnFzvQRtw3o67oX/DNZ+dn608lQtB5eSzXi6nB+uXm
s8w7mv5PytnDI8roncYEWGTHgg7qhbGkAchr+u5G4M4ghF4NrZTApKwY5/cRrZTaBUvzxUjPbIUm
1qho8paoIwCAiAPNwPI4YnJ7VbO4/ZTBidhRxjArQyTsfmXz4gdn/jWv+VkM7nmm4+Ce/uvBQLr6
51wtBMK9gyjvnsIQD14Lb9IJzEUZI92gkPdNwUeJxfOZ7JjHUh6HSyk7BstfjY2o9Txslw5u7fI4
PxpRqu7xiqM5Tv49qYgzVhC6yF76CjLDsmEAamxdQy74ubZSihdSoaT3orWzJA9RgpGj7KH/vyIl
sGbA60DPu9/ifPRBrVS984fG5+KWUeXb+dK4h4GFpQLgPX9NJw2dBJsTm+YoMfjBtzAmSVDzUcaw
JsKcR2G6oVZtDou+cVoquO+z/LRLIiZKDJJ87RUhlx/0jA4Q5GINzOqYN4hbCAifbzykmbk7mycN
4IfS3iCw/M/llQOBLWhP7QfzajMKTBRZi2cPSscilHhqDEHclYdF1jI/2LXwbBdVw0b1V1xtuI01
DZtTyOYw0tDNUx2BvC85gOZZI9dWXspoZFmL8bpUmBapa0q9Xg6iiuOmtimgKDbyT3rXe7DpkJrl
OEt6pPMq90TTm45DdEPQBnmsne/xkODVLms6kSWkUNXJDTVYn8wVuUCD1M5ahJWWFuKWKh66a6rn
ClpS71frTkxjMt0SRQmq+zroMeh+gXD+FR3+rAw3/bC0kjAsP6NykbNBgSfhNdSMG11mfbf6aq9i
7iNdcMz5zhiJ/fJzEeaDYrpjo5ZeiT7SBGi3uRvCquSW7sGl6PMZe77U50YGNkFi28oJFlzfoEHw
7G4uuqxRLcNWjKn0WW4ui5CSM30VliJm8sORguo0Jn1fpeT3T3Ag1WsAFA6aSFPgp1qqYQuhNXQm
dp30RMpvWoh24bUftG3d8FUokEzSEjtvCqDCMI7seL2xP5e9RRLbxLI7Rs3/1JBIJ+Lmuk8UmGLe
SWyY7Aqa344/qOQmoj85kqX8RAVuHYSwYoW3A0lwHgI45hvtY2OAxOnRdXTJRokf0/Vn7mqjiZgv
DKon/Gwwbyly7JY86lDbvU+aXFCX+PiD7NY29fg/xrz7EIQFCaMVd+RezztyfR2OBC2FVS/m6+/m
ZXpPULQtP3FZiARjnWAU1/WyGjbVyeYuagI9ayTo3hQmRhs2nxKqxpb6XbUlgqjBmNPfzXOEpQxz
MagCaGmtqKRd+CsR4A7eCmMdMOcxDafTQTy85yQgPhjEo6EDBI2wvEbT/Xb9+j8x3x4JE6OHPWQP
1se1pm+7xkXNd21tn3UegO1FUkopiFjP4dT9rWbfE97FtGw3eOPzKBMyxOJRnHzlasvuBEbb3hXe
zLDPXCaYvXgnnBDfItyQV5Q9bgZzTjFG7Q/TjkjCd3/AjZDE9ix0ZQvFA6OUP5qokKUnib/4vuX6
qnLG/xAXxJgPhyAew9Tx9lsFNLIg6mqrDIaPy4vgrxE8qGUHQWInUZiRgXeSmrl6ySxxBbXVA0Mi
puqfrgYqn60mkzybvkaZJVZuKgPeJKE6+kLlhbFb6QRUEcVebsOWU7NMSE+M35vOjX3qZtGrWv+V
UeYcTBgkQquKGrLXj2T+5nvQ4n/zkNQu4wOHFPDHOwpd1PVj54NB8GxtdK//G19WqFCnetGgzwcY
mqpEhItqcPBnGSUHKEbJ+n49VqZVZSKeeiseCNY5nXaHkhSuusXHhnjKJZKzUPJH+l6eG/Q2pkWs
AXNGMmMXSF1rQH9bv7LCEpCq87RGiMAOkIQUhDhzjLRZReAz/k/3gWCzR5cpmj0Q2xAoPanbKSs1
QAyg+NhlikBBscdweicQvWGKmpuW0GJHvMSQwuJuflq5XnUBsecW0xsviwaf8nUBa7SKpXaghSfO
D9VCNDKc80ZO3tX5qdaoIM2lBZKNIRdDlJhDaQ1Bawaq/D5N352KnHksXHe302u5sqmQ4ctWRsGs
xGsxcWLKWRZdR4P9we7eGaqsNZWpOEJk8oN4PKlaJ05iIrdKCejVxwdsm2FtShBwlzMpR3csf4BY
BtuAPnDwkbN+exrgzxYODr31JtS0eCtyJwdXilLM8GO0nKIWmIjrmKk5Heoyv+ZnMYtE/pC9UFBZ
Svi0bMuN8/nA9afp5v8JobFPwXtTGgLH3WZJI0fxcJw3kVP62P422LpGc1sdMfATI9AhoaHWrH/H
068aEeVYXELeIk+j92WzERL6Aoq1w3fv5BNWz+kwXcaLXvFNeUmnnw27lyTOnjmJjZF2la+ClSaP
5t3F16A+TnCU8qRM/62kzcjZ9R/RVWyihyCsxSgbRxYSDbt5x5AQ1/zbBQLJBN0cg86dZde8HurH
dUIUPkozKFu+nM3VifIQNGnvyOYvRu5nmrK65B1WtJyq8JN21huFzI4yyxeHlDI1RAunGDHEnp0U
rxu0Mq+iOMZQnIrGb3esypkk1zQaIg5APGI9SkRLhmGG0/mRDFYwkPC38Fc15rraPkBcaaDURfF6
jo/ejHsSYUDDM8sA9tJ3diF1wuyf3cDzDImIZa6TDquuotM7q1RxNTCiejogxJ4kR/D7ApEyM9bu
/cn4Ebd6diiBHFBNwK2jwizhgaxufHRKhnSX1yvx1/lbAwA2Y8HjW8nt4EdahsYj+QM0sX0k3H/G
XGNS7/FAFBXW+J0pljP0+Gh/ns8xOXztBg0iB/MLiZc7QsnEqN/+0dFD6/6LClDEjmeoM/aeGksd
VUt4m7n0S1pzBmyktoHztDfIJkpERRmPt1Jyc4Gq47Q57cb9oDqPQbjHLyNfK76RRHGiE96qP4DA
8ywpH1fLXjpWCm8yDy1fz23Vygrq2EJs62atwh6FS+b+Nrju2mhWJvySK+S5syaTSaKHeTbJ5VLi
asfWW6ff2otcvLYqzuJnDR9stgHWc0JojvhC+ip1X7qU0ttjVSxqAL6YqXcVrtF//DY6+afeZk2t
yJfnG24KyxLwqx93LQBcCr6Rb+9BOQoUa3c6ChEwHd1/aFBlOYKelZGcthaaDCHwpC1HsCT/KqiN
dxW0HHoeTHTp9YTXmf0K9BOmvYHBhGt0zAKGo8xGhz9XcJU8a5SkIiFBllHkOfHcwLtxJhHWET5R
Py0O98L1LlsIkrm0z74XZkFM0b5Rx5+NRBM9NQkEUpTffk20s4sz8Vv++Q33cxnO7zgSGHrSw92S
2ZSr7is2lEFHZ2Q4Yvz/bVKtkqqEH0x2zB669kWr0EMkKqVzbqbreoZ6OcIecuu2Wao0FTkARKto
535PKAM+4b+exQ4HLGH1aLUmqebSUzAcGFYjHSdMlmi49SLPYnv4zto2Vp1XT3f+4aKRu4/QB9UD
tB41R+Laz+B2m8CU9PkScYgENvFf0eX2Obuc4EABOc29JhSH0IEgG3jocqhTGC3W/UY/Vi1UAZ4N
kiFB9puV9/4p3dTJKmB8sN/QzhflpnzXM7tr2BfB/gcURaG3C/LcsU32bKW8os2ZXtrez18yNHaa
P4Fifcquc6EUUnDx53fIAw1SJwtOmt+2mRXbpP1XIk+PnbiithU9zQnCYJ5isU9oeSzC3dmmcakR
obT4Efyh6b4kQgrdDRPo4do6BPu3XDBR/suMGFGyq2PaN4rFHchjQFNiHAdE4iHywFzcv8l3blVO
zoY2ONlggpNdmfd81H3gIwpOkjGAfXXK2o08kfDFkbiU36SCnCly96BO2YIGMlHhS+AbtWrU1NIL
YQiFZOgcSAyrySLmbGI3mwIGlKa4O5UWFB2B0jMIKIuekh2zN6Sdfk9V1ng0MTgh/svaIbXFzUlE
dy4mgG+4f4FKGQEVewsMxAKiHC1Nw0SkoC7GIXRrxJn2Q711UjFuhvZA4mMfPl6KLTAxzscod5+R
XMrWOVbqJDpofZIxcdYuiafLtrZBhRL2FbcALA9hYM6755oIg4NbBve9kNgJc0Efxc1R5+cGLzWf
M7gPphnkHPa13rtBU4zAnqaH3UVwE5RaQY/4f4KyigNhsSU+xe+9CIRNkGe6kmO0IN6nEP+HIUU4
wNUKrwjGV0fXRFXmQ9jBF7TYfJoYTGQf6m37RPBL431xidvhp6KEwQlUyw9lrMv4dkQAI7+0/a2e
rM0O3+ZJGupKOmt3lTo5iR0W144/dcLin6/3Q+wfsqiLbf9O+xOUccHBZvu2v1BHRhF73RrhEFC6
5Wy/GOBGCc9KG4F/v+ExcEcwea45sTqiR39+AzXeT3BokBBdOkmG0BaGU+/jz6x8asRy18bN5uHQ
ox5wJ1sWmsez7yetOR23XmOyucETO97xmq91vpzAhbrV6xXdYhzuxkTz0P5xuGri5kC3xBPku+su
wYFhaRy7xUWMUmSrPmu5vc3Z+oZBC5Em+ryRcUxSXnqFJfoQJT8Idmo68vyO64viACBX9SPyY5QY
xDuu42Z17yOT8YBKxcZEKvZBQV8hjuNPtlvwMKgUidbJ8wJvs0/SmTa7q0F278DrWuZVWYdgbxIs
vMSxxkvKkuuoOe/qopU/oo2rw/1Ih9hJq2zEL1F8mFQHqX9EsQj7hHqxgSznFwNBt/cUr6BFb9d8
IOqUKTgbhhP3Oal4HkA0cL1PlqAqakOEG4Wt8WAVDMLVSCAA+4lUFI6Sa3HpQhYGOL22X5KVFIUT
gOtjrqILMY475B8nS/etn4W8j8vKoZJ2EzJZKw/MCNYO755v0E8O7VzJxrS+XwRAoin3+hEoIAWC
5K9yiC7jjacdBdkdGZP4uNT38AhXka9jgJ+YrKel4dnjyEB1gCrVS5xiESy30XLWLHEiyUDMmwIx
CkTYfcw0uVc2mp1NWsf+r3kCekRGaJyMGuLra4So0BN5LLg00MfqGwsy47gPMl4JIyGpRDtNW6LF
xSHVR4KnkpPWenVQ09ZUnuwUHt91eCOnHJRO6rs7SB7UaOdarqRO2kKBLBTCoks2yttO+UOnGgTO
t6oP0yfhBbcXl/aS6+FuCzWH0CIoEo9vkJ8yhD23qSFBxgOTgs9QuM7RrIvEQLnykPJAy4AWNEIc
R10ebQbSc4vUTWtfoLenbWBJtQerRq9PXP8iPCbjSL7BUVcv+7kPGr1j290TH67LEnXp6yduezWY
L40NfvVNX+G0FX1pbk/smqseg9hlgygrTgiYyUDwvXHT9t0DAbp9N8E9X86ugglhWjU0CT3xDcoc
3WKOHDsJy0LHvrsdbiWteGrcY2sFZxQWIYIMYXPIPkWZWI5+RLes+myajg15CwVT2CF7k9jxiUv2
kxya0JK25X5yk/iZHoRbtR77C+cnRbbIjLtK0rgpSEdbpn8qwhuf8mbhI5cNFI7e2eTdGB20+K1X
+/ziAlvPz+LvXSXiMtH/DXdh4GagOnmXNalLSZ/MxeHP2X5dTmI4AxoYhXYhH95fwdWY3ZJSJQxe
sahWCEup+VO1rS3lRLnvyAAZbRG+/gllLzVkLzXSEajCKlfjCZfTOtU3+NNtjEfOCqxxrJRz1479
02NxTnjUMEG2C4NGsWn0qnIDrR29VfBKtsFK28QrkDo7LBZRHqmdA4xRBhUy9HTfzUrTbR4MpYYF
COLKwKFwZhs2t97bfTP8V8UZVLnN0L3YS98E6vBs8jAbCfRhmQeWpiR/YKny16LSwSldXJYUKVk1
EqqFz0zb5l20QS9tBXYiIcMTEE64iEQwrqRLfI7vtbb+ChZNJ/awMf8vwIFTrCF0iwOQ9h3v5Roe
iMYuKvRFoI/36GhMMULWCCnUbHcJmQ7xoc9fBCKIMiRPmZmchblw2neZaYi5YjqxzAJrKPnmXCaN
Ly93gLWz/6bGdricXmtC97yFkNpvOorWDULSrXFqR3A/3GnACvtQkr6V5ZfgNT7UnvBbVsYYpWOn
comelFbufTPYvESt31pGQ8P1OcQUMG9bwa8S5MiewgXGdyAVmumrGdMPmMcUMLHgW+v8aUF5pSBH
BWmLE/er2WGf0avSGqqw/BU8mLum+GwP1/K8ieoeq0GFZ96St1NdeB57t/pKkN4kVA0Xo75b6NQ3
ztvcNiCLf29lkOHEkxXKSXNMxtMUna1fdvQ9I/egu2D1Y2ugx9AFI0hSV2w3IuRlQufDQ1N73EFV
Y4jrpl1dlR9izrFJa3wtqn8z+qiUgoMBSx3UGl9DC8wqtgrj+Q7jH6iLcnNvhQoOIIhCGLZ63B/V
AzlIA5F0xkHsmGn9qapO3xsy/DTdPLe6XQqjthNTpzZYeyhODBOpu0s4mn8jZ3puSwbD/KnhmY8X
2kfTC/J3zK1GAgsImzkxpNvQPF1uOTVYI+MBEcZb2FmiC41WfVEwbmYgMOjSHM13fBeRfwUxwUKi
Wr5EllbUQpYGL21XDQ2qFM5HncMpasfh20OYR5xJcMBLnN/0V9CJa65hHVSWaTzno9Av1OYhe4IS
jqkQh98xgq5oJTK3Mme31Q82n2qhfoRQWRgAlIIjJ/m4sX/jkZk/+jjt0Xj1zlv7BeXVKULjrOLh
EZyxizIaDqfsmv4mxjsljFLgjtnW1NbgTG0/imcLAoLbOvp71YuKb8xpB5j2sRQRxMU8vJqH6DCH
QVh50hZldKVm57ChvSR+vVmJOIUiuGhDRKXY12UGQxJEPTYWqfRzQT8zEyxQ5+HiaH6Y8ccl+gX/
Yh7SRh65tI0N4whrO6lPVzEQOic5SH4k8Lbkx6xdSWkqCX+ijAXpalSvjq/c/GTnn41J/Py4lCPA
WVCL/6LwdcRBSUsUrigGPo6r/Rjaiz9F0nF6SPtk2KToBWAyd2dBjoGJ8v7vb7QqViaFpUoAdIcV
B/JxoH1R386m/cCthHTNv9QtA8SLPtossCx1R7mLX0b/bxX9QiKuX0eA5Jsg1fp4TMQbbVyEd0Pk
W++OdhTlsOM8++wAg3dPJD12r7/CRN6j/z4BpEAvyUskiZvRmNbYJIxdForkmBPnved6s+jhF5Z+
SDkh/5c0M403HhfcWZWzzKFI+Xr8iETCe+I6lP8FP/sS9A/iyizNRIdgfMurU43e3WKJFQ9X0XxY
wLRji464YkNocokbvdWnVF6YbWP2WuMnLFMxn3cS7aoyLh8jjqZWpLN08WR0o064MIz2MGx2w6KX
2W+apFQvizm93e6YQ0uCCkWXslygSk3dBCv4Brqup+4XOxbPgvEIm236b8qjZWdkUCHKv4UN6zNt
h/q3/PUjRTYKHqu03mE1o54w7/jyr7SGLO/GPEtJV9wpRRKOqsaQiazZZLqE88XwR9E/OHuPE80D
KhYUWbF74x1GAP8VPn/Jmp/vCLWy5+NEAMtbQA/dC07U89hrA3EYWZvVEMrHmoVo97GCghZP1wnc
E0QqJ/mcD6iM0rEgJ/aGyJxBEZrofT+9A9FXdBVqNaTDx9NArVs+1LNrGoQGB2yQA76TRugSlfLq
G1fLKm2YpKiRPWtQ43aSzCOzi/VEXmAaOabLlEmPNjlITRr1lCsi4jAcXfuZRNBxEvK0NoWEvead
OZQ4YPYuOU4p8ZSvQIhxcFsxIlU7Mqboa3sM5UOAn1FTBEp5GnvnSfR+k0OrnDJ1NCkfFAB1fN4P
s0BnuULKLlTxb6pKg8xh7+84DSbdBqjM8PLqDvgX5xP4Bu36GB2n7b1LAU4897dGeP8hfanhgdaF
7QUFkEm2o8/Bjn7rrlQOWTRoURmM55RFVRHjNSTPkAjK62i1rdSxsPo9N1xg6HbyXdUg/c+hInJd
IXPlJ0M8bkGw7R8UR9f8fQ/wbySS4qEWbh9VP+RwLxLcTvYQfPCxuYf06t32xmuwr5YjMSBR2r+N
vMPBxgAOuGYz5jtmuNcaLyKg5aCCXN3gAX0BSNTCD1uadstNYDibdh5yAQQC7YAKu85ihhzTukjT
zIqXenVMrYMTpy5zY88tEq+hctbowL/FvWfPSThxKMLpvJUUtSPyjkgaOo7a0TxfyX44Ha3XwBE7
HwOY1QV3RVae2VLBTsUKkv00GbSZmR16/81WI+yV9B6qxPyfU7jmZY+hYaoQutYnAK2z/WJ7l6gL
IgF45EQ1GwwZZdm0Y3+9rbz9xOXVkAX0x8VC9JxzJXY6li3pCpfh1VQks2oFnAVb9AYv7W9t1HD5
5I/zDLwN867zDm7RKsvBDmjqk4/29VBl6MkiBATLiSrocz76OiGtMvXWT5url4hwF0wrbBG/HxU9
dIczMSH5eSbWPmtzotQXedLbEDPWINIPLfd0U/7e9PlyMbgnf/TMJBBg7YrSx4qatq8zN0h+zz4O
/TaPSYLqEbP2eusC82pmIvzxZ9ARsYgbjXlRdJYHOW0sAV6AivjyLqypRpKc0fZ2vA2XuH90WmAX
mY4IUdN3nEiUw30JtL6Nw5lFxKGfJr7x/M75oKXPptySCVrc2hXj7MAP0xPQRvf4Ln1jFbYMJ9ga
0iD97pavipdl3RdPWViZpL0guAiQV9VsVdiuE1DlmoCbYyy+u0LL1OPIpxd0hBFRwuz3n1oSC0GZ
YLko3zVwHr5asr+wmC8KvnYa7gdbs+v374u8yX9Mt3svrLT5rjBqpo9xWd2Bl2SBznBF1JggnaAq
kFUaVDRVdHXpuS5IWX0Of/i42pgazsgK7zEUu47qPRTDJDboAdonZz/MYf79+0dznfKkrwr+Hxkt
hX7wX7IxusH/8kmoL7CJHGrs++LopThvvJmS/zUIXQr0L4pcwg4JX9Mxcpqn5hedN9KCGf0KHEo8
hSBEGzceRb87CtLhx5IaoNDvfT0mAK2rFfCAQcFAN/Hl2Eg/Z5bVIE011uM7QjFP7PnNj0iuuSKb
/2QRaZEx8si70xStbS3Ieu0slDcyXoo/yVQ7f6FIABFUCkZEKrN74jQ0VAzQst2KUSAy05fht4G+
4cP35/DW6+YFJqBY2FKHfpVV8kRLlGWhnMl3qB0VZvbyVJwqiAO0AogGk1JTtURDfu5QnrS+Fc90
o0TjkamNIT9wYKZSC5RBlX/j+qWuAoxZgAofFDJDCIJfIHecxuCGqXQ7ij0pvV6efboVAzO7Gmix
SaUi6iDjct4OIpp1hq1O7dhtpjWpKnJ0yuRvDRDMcbAuT4Z4bac4ipbBewVbjnILeg1ofCBN4R7n
qpMXxD8x1u6opLa5BXBglUsCtxgQoVMSriPxUyNFvPNvFtvsXZ844mPqlAVawIhPEzjQbbJVtHHA
ixmwTLjEh4TZjxh2Uu7UpqFzOhNnlfjaER3Po415qwcNLG6U6Yp+cSf4QXopJcf8a3jQ5ZBRBfi5
Nl8zcFo0AW9eLMiqI5TLSI04jqfcHAeHe3BGa4wpIz0HD4VTtdI+0tsFargUlufHx0CVDqh9pcWc
QtLSYw2c5i9wnHnLB0hKn6NoJpDn4ejqsuMWmLtzs+trL/UiPhg2h+3s5ZQ7CHwv93vp8XLyacqO
geueUDe5pinKtfvO5NgO8L1PemMXRmqBqYytaBclag7DvLt3B9jNsac+uropUAfWwNvsfMzPcAYj
ubt7MQRPykPcagKyGy2nEQxG9+qO9ZajExuRx5LKL29qA/Ld9OwFTD+TXbp57JsWMDb21/tg5pLw
h6sKGA4HbgXpdP64t/DBYrYkELKDvIPCGYUmirCoMgVqmy8/y0ad7n0Pbanq1e8PebPL4gyBx7jZ
BM2ZrISn9AUrAS6dA9f1aPMoTxGfNp2RtIDuqd97frDCMt69eTlRPA9JGff8QjXLgshHfTAcfnHY
RJ8wcktGqFG9FlAkfehTjgTklBnKNMiA29tkN9xS/FZVbK0UcAuPo34WJOhY49BuGWa5FsAYXXIt
PiiG7AH0tmapGBMOI/XS4kWEkT/eTYCp9sk6piXJk5wVWXBe4g+p4X7tUYsNSitte5BVN8iuqHXw
NyrCeKEcN/vQnWyBdeMLNUql3zSpOawbMgUaP3LCR5Mbx6a5j6KwfQOHj1WoL7znIqEmODmtK6Ga
0hQPmgJqln0c3mPRd9kfj0tqiWVia3jy2hR2avMAiJHpLB9l3gDpbyIpftYdeVDuZVRSTFm9x6yb
TfnnGezOl04NIeCaoKntQv/5QglrmSXKH+Os9YqdNGzQK74yImRix0rtosE+TRQg421j2w/5myCm
t1T6t585PN+Xd1NUdPH8PBiqZ1byz3IQdB8ocjDvfBZR1lENf3OoH7y092g/0bE6pMe4B5hjIZz8
Izs8tGgkeXIA6IiLLs0sr/+Jtzcn9NyDxw/FFck2d0tNKyHWhSwC4s364AVzHv5aI8EoMQ8WZFXB
ILmi0XTPox9JaoTww0UXWr8fnIAEVDEv/fbBpaha9BGygWwTamAPciGtDlCDx+VWz8dKbBRhL28x
m3jsHa23JEr21gDVy8OJ/sT++wUcFIegEiuUqxIpOs8aMFfmafqXRVuGnsapDtDgUqYbJLKk72wn
X9ADBfTA+3ZPMhcRNQOjaO5CBR2g6olynkzOhRrf5YZpYRMbszlk8FlPfalPGO1wSIanLG4XZkmc
kOKnDl0Z0boAh1xLchy32lCV6ltcKNCsNUvavn3ANKUdwnVKgCeGgy5YnS7nHkumNE+T3hfLf6HA
viQu+QqJHtkoyBcoiJW9Bq+W+AoSHFvrI2UjaTutQ1N9iEUTz38U4Xv0J1FD000+fRJQyYObM87I
L0q3E1hghbNJDaBF6lDK9lBuWL7vz3kGuyzhJR9PhZA2bwoBitYdoOa7VD8pMqlLMmD9g1/KNNRP
nY2+LPGEm55+8yWSDfH37n9348O5auAVxutXql7caD6SQg/3TPCg6j1kwao5RB5QKujCP7Dl7BAf
ZdMPpHGsvjerOSci6eGfhkEUMqsDSIlvjnQjtz6HPU5Jiy17L9LfzG2RCAH4527AC5pksGn00Xai
3lh3KrEdLCT0xqfvP9I+iBumrtqDwSLaeOStHbC+KZ6cwJ9DyF+1HXsOt9N829ZdfnhsTk5YlOoO
BGzQkqD0SnObkR3gH3IbLyZBIXRddCdV7JBYy5yicHL04DOJtSM5ribT8bY0Jl/my0L2MXDwz8+i
kGD04iACwYR1MnAcdcUhJv8GXdLL7W35nIAtT83FGbR1r+Y+zSpxAS5y1r7vqdaRVmwiB4dLVJ67
5vsHY9tK3R5JWwSn5LPVMKuAvOihIq64/W4/ZUsWc8Gn1bHZUXtwFnnQXqxdQmmWHzXu4PLQcAKC
w1JbuBOkzfhau3geY/gtfoClZSFV3rkEp0IbnXxQeQIq4SVh8uziiYAacqgXsaoLyseTV3XhfNQd
M5Tt4Rni9Uo8bqlySuuBRQuGxOm3ZPCWbbUYo+mYPPIwXloH+6Y3awxW1AJ6LlMBxdZqVWg4TRAE
XtiM9vURQMcsAHb/1Ibw9mhd4TYkQIiyvo79gNji0RukGGjtSLbDOzAQtszcB3BE2F+gQpUCiO3j
fDrHqT8xP4+hV7kHXc2+OJ05/8aB14GEan7K/dqSPmNwQa/RbNXtcax/EyAo0qco+T60W0WeXr2h
iYKvNfwRxx939FaXWTvcBD1QpoPDMhXLYiPKW/cuUe+oJoWE+995c5qD51ql+eNDgdgOE/D5G8kn
Ip2xaGNW1wFX+FGdz8FmFK2yyCdaFK0ydnu00KAoHViaQTajExW6MXP5u8IW2PgypqW1kJQDDjWu
mefeHZAJU5brwhh16pvTPQQvsPeT7yPqFcRIYkOOtRK8Bq6s300x86PrjyIY514hMPlMEyaClMGq
U9jH8Hq2E20MYw6MXabwsUBdDZ9j66tNE8/CsLHIL5P4gS953qSNP4cDUoX4esiXQPLvVX+qJJti
She7pPzTusf9hO2NLJUPsbUY7yWzCAsdTZtp0EKXeUvjLu/GucOK/CWWnqO7DkFxb7nBhrNLRMIl
B7EVGeJFud8OpayCq/2Z1Wbz7yIaxF7ALF1w/Ijz5VG1GcgD8nx3grQ+UDv1bLKB6/0rPLenzNOf
Y8eG4UL/7Pr4Z2h6Zni/b9SUtZ48KMIIr/eDOF7dUKRLgd9d1nW1gx9tI2UfWWYxgbrBWZI+a53p
xpVSkZJ1SqVlslh7vwxZqFN9oiM+lcFpSp3uGH9DkNno4R4OyB+XQSviBO+QJJnwuH9zc8LwvqGs
eBW6Ep6Y2nbnK8dEM4JFMpIKfNkPa+8vZqpURp7IMn1XYLFgI98Ckr9kXAp+73HSNMUuHtYhARSl
R2QToPHHojfdVIB06x4rzjx+Uy0k1B0/bASrVVsERoczL8QqrL0Gp4RHdirdus6qXRZ3RlG3uhK9
phX4RUoQ+AEN2dPX8iGkCN0GiOgLwZ/kwMcoNepTeeTUQKFeYImzhPDzG/I9NfiajMLWuWrGuuB+
bUIiEDShvD6oy/iiHy+ooCy3B7LRaF7Xm73/ZJNhSgwHlwpW71qe/UO2l9HHuneX9dKvpevmooHO
zl1+26RqQZRGWNS7hE+PTy/nKhMu7bkF8eycP7l3MquEnP6aiG/65Pp0aYIlgOxAUMNBIWVDVhWU
iCMzuo0ovZws7jLWnOAraw+wvG1SjggUzkeP4J04WeTSxaJM7AaKo9GVW3fh/D/Uc6WLQjI0tLOM
ocEJv6w7fGJq5CgjX6XQ41mz3extalfvnH63GiD7Ng4hnDsYD1kbA6Aq7Iuj7ch5qgGRqcXeavsE
uysGu3/KveC6lkUnUUOkl9u7klbyH93hscfFUN8WkuUDiyBzikQXVtl0rSOOMLdH4q81884tYZNh
xz5Fiv5K0ut78vCEDHDHLyUUAbgpRrxvYO+jQpDm01DEeYwgmCCogeI25wyAVhQ8saYikX8WJn3Q
DZqj12vx80Ld1GHfTVHkTKcUyv0vkJOTxkHAQZ/uci2nOKhESbZFhNbsYYom2gm+c3x3TDlNh9yq
j18OsJfN30+ebTyMe/ara8xsrCuL17HvUdi25Ze0lSF9ybv3Nn7taCMm/eRau9P4CMNK7kGJq/cN
Bl9bz0pyojLiiwTpFTKsnECmKg2becUJXgD4WEFzcr+9E6o3uMh2wGXemjxkZtUCZzy+C9O4WX2Y
KADXzUqTmj3kG6keXiKzpxAGupMnf59okQesChB/QXeODaBnONVVrFnu26hY+Z0ylHb0xpG1x/5O
oYQMlDY2EuhUYS5AOpaTvec8ZzBT0eGfbLisKvGH7NaPAoR/CAZaPb6jI/AWl3XkkUDXzzFPqAyB
Yw5g5+T6DtPOJsm+r3Ik32SBP02M848aZPAW87aedIdELJ9FnlTKlQRpEPSFUEyxROb9jc1iShEX
1LXYieJVlLWLfhHEGZ459GztK6Gpdp3VbGQhEa6K8ohc+eYH2fOaPdyUjudiuUOZx4MawbrDBWoT
uJN2Kqu/u+iD7fVIKzbNlJYF2gZIOFeXI/7vPJsLT9Ri9BWj1B3ppLMSY6ERQmm+VzGDuZ4VHUYy
VilgYiqN0/f8ZJcqzrt2eluZMD+7G8GJn3BcJu+35KRrQFQsBAHMXD8CzXlJW9pXr9nXJ27LYQl3
0n/YdzBaVxM98dEsk6wgw/WiGiQ6lkH02Dq0qB77rmLcGq4En+AqmVWBXSFNb3iGfhOIMbZkPi+r
+n/dPdmfsJE4bYPd40UY/P412gn8Bq7lNmpquW5qKQqB+cdOoGLLoVoMfwLwfpW7YWj8kFWZbgio
f6c46vfPbNlqTg51OXFhWnpn7CNMPg+yCm/wodI4RCRtQ9sOHul8H4JZRU0lkHATKSdIyfJynMIC
zGjBTTiKUyXTDElvP3MfZbmdt60De3QKGSpERukLnaRz+ylhy+nXBnPhGabVjlcj2NdXQ/aKnhhc
w9o8yJySSpNixxnwfOrT/JLmgNnqK/HnmXkM7LZ7R7CSdjzsLXd4OWxIt7he/T30hkylj1eCHpLK
nTcdXuIO0bx1zmo6lE0p+z5hsFwjl5+aCNOOOVE+M7J6T2nmZdbFbHLvdVHt4Lk2WUSlDOHEnw6w
Ta8aWhi3jRAf5DcUc6IMqqJNN+9U2WaTAkCQVlmDZrxgB0clFjYfmqlIl4SvqQxYmQr0tbqdGRoc
Z2OBdQprJSaANIz1I8mSOUseIdlctGeC1ehcs+yFlDKrWHddEVFEcQmwirGiI6oHUg4CWHsy6Aod
55CDeHdYwrei2K6TVFxTTKjP4xQ+L4UCSvhZTyeX0DmzxsClGUXv00Z5m+x7f8HOsjJmmAmdUGI8
4Qi4rTxreR/nRXPBYIw/lz9UTfvrw4MCbb+xWc5mMiM01dRaJn2cwPj1/WBFHgRS4SImTjaWadtW
Ei/qnbWondz2QaIDbGR3w5UbJxtbOIIVof8oqOte05mJawedkF1r/NRV7rlrzKr9ZPCNCE+UcSg/
YOxgosEgV6yPPWMwbuOnx0Z8TAJYxKbc02By7c4hsGkwf5ZgcD4v6vMnbik8CjEJP7dySeU6KHfo
wN+YYhja/pohIVhiF9hUaWhc0m6haqHfXIvNaWCDpaw3PJa3CKkTOuVF6tLB0XbTmQ+rnLppg3ZC
G/vAWZK7xBOZ2qITpiOIxwzd3aPoSyX4VdGddF6BC/zjsg8nlTJq3K53WpLOkZ+Wgkg3NIn+w7X3
0mx7rqh0QyC/RfOYkQLw2PHDB8zChvdF2Pnqe3nMKqwo9CzFRNXScw6NVCAnkXiQjE/PopgTHclE
bZUodbjDxLNTHXid872JQboGABV8B6yp634EOcwGi5GKhnoCJ1rZFqGFpHRoGZik3qez0PiCgHC+
6ySEw3EwyCu8xumLRssbMO7CkyWzlnJPeK/Z6w5+gUE9Wk4TwqZjNYZRjZlBFQmwvefARGRW6XI1
oroFcTclbraaVgqUvJSs7u2fMxKTSK3+DLMH0/LpAqHeg5a5AVR3GeY6136LrWPqWp2ctazxmPRc
arWT0OKWeD5XbSqoFfRpLDnHF+KqYBfj2AGoelGn+wg46XMsj5o6IwPZFz3RfT8k0uqXrbkvTrI1
AYprHCe1qKKc4zu4NNyhDHtI8BCs0sB5vcaRvuik+yYYLC7WmCoy0iirLaAaEhKJoyRcq1HJo9cp
BwrKBxKMd6hQAQsD8AkHE4tg/7Hq33gLF4pqS+kPOq0/x+//BdscDwzJWAScVVrhmwjZdX4xs2R1
h1jX1eO3+R9nGyyqz7D3QqaA2JZoturpBQk5twcey5nNWf2OZpP1GIDWqtvEzw2RnxLh3H5+5itA
Gh8ka+vLWPsPaed/I7c5MxraFrTzFBo6Jo8jMmYc9B81Lfv5gop3wAOlzTMWEte1iAUP1d0x/QM2
fI5PfEvjzUGDa4hcjjnnsmgsfsC1qFDHTpFkMqp8PQDGxSPqLkHq0ZWARUE3NDvQTogZLZj25Eh6
eah/3hojvORQ0aY0EgDE8yXABqg0Eyq4gL4VQHeozSrxoOI+dBvmnWFXQHzzRaIg3YoS4PBuVdGa
dGLkVKEM0EI5GFCBX8cxsDF14L6hOX2rR3XJr35ARSGGk9/Pd2Scjpz7tGdRhWXtvBdGZvIAv8/K
8NsJDJJLHeIiR7zexw0k3uK0bz8qYc/x+P6eik5lFbTlDgDFrQy5faqrZmiv1gCT2CIlQ8TtXwz3
N724pPswB9uh5+16L9hiJbWuyLrNdL0D5TjZLpbyBqyiPnOjaOc5VYRgsne/XkDLLWu/mvG44flb
1QFCuboAaWrEH8q+pErXW6JqVuooBWZPnflA96G/x+81ozlrpd+zjfugEZoV68z9RYMLOEO4AvO5
ejDtFRPhtLqM/V1V2g3cSwdbxd0KVAju0Eto8dQwpfjx7AUMl//h5wKNadSqiWy3I1S/r+1AjSfd
e96kURGWH8+IY7rxVJ9UadBEc57SC8n13VS0tYp2FpVY6NpogyCYcliNfHbpht0XMY2bzcxHdpTA
zbMIytT+zdOJ9W5lgcWX7Jl16TZko0jqs5n4YX9snUhHejOCLzLpSzALgIEIP+Q7RfIRamG1yNce
LayhUEHQc6BIqhRecGe5/C1NnkDA1M0T+TUn+Qv9OgWuM3zr08MsMOJZ1ImEsAtTyYkS8NhqCga9
ZcaUnRxkOHfEVEkUwW4ub4/yfWfMOiawz4cQnxmSAbG/7zFEaYO1o4tAnJDN3B28Z7XVCxuD90ha
9JSjcimRoJHxECiLo0WioQZ0blN9mHqffYv+12wIR/aTS+wmyStftGf3n+rzFlzq4olda8gbW3bj
DYn373YaxDgUfWcTt2Hh17UdGy6BpkS9pmfrKpr0fsGRZxTf6Sr6gyVv8LIvuxsAal1ZLm45lZkD
X8dF2/RgrIa2EVU6fLvDR6rcQkI8eZG8Q90I8OwuPqev8HF9IDV8hcdoxqS3m7EVsB8Is6yEHRpQ
G54y7t2x45p3U6L0oqC7fa48+nkJGpsvwrK0lkSe73O8gjhu97E9cBUSgmqWXq9lbnEt8GDXlJwK
lUlGxmPeRQ9l853lYPPs+SEn1L5bcK8qRG1gGcmKH8jIEMiXEGMJvA1cC+7vJ8gOxzanAtXiDqZp
0W1hWFSYdoZIuvDGEtI1nibUki/Cwg33UrxmKD1Eun6PyvdtUbt5vFAD0bPfB4OzHdCI9m0vFSW5
bJ2tbGsGJnqsypoRI8VbbmWotd3RpBxwX1QhfEAW9iuM1FfWpj1nV/w2aODl7qXu0yXL+ZIubWm8
MhSDV0CyJV59mb7xm7nJEX56GpoyqDe4/ScGYjWNQmC+eittm9uIchfxHFWt+HAGTUSCph9uBqk/
gHRM5JDa5+TSKIN+QqKDWiOwaZpufrtjHbaHna4XFz953UX+8mfWN563HxcpMBsXPBRknBl6Kp3d
L8rkLfWDykcsavSfnltvmkMa7qSfCgEz3lrmiQiDIFnNEfiAUpQpk2+IIjuUqKywzs/aoFOFjp1x
xqiUu1pGplsSfhDirdDgFCRnk+YExIgS2Ek2DPStz0tXEa/2msg85nOwOUKiLKxel/D0/XIN789b
RM1ulvKU5YCq7SCCW1apP0H4CMvZZUL97CK7kr/gvYhysW0+GTuNMnNzyUwfPDMSdyJyIK9vLVWb
1e7Bm4evoy/wIOkOqWKEeKN34owgrN0B3+X+D5MvolW4ScgKrBheKAE9TQAQhA8iHHFaEJHwRZgo
806JNNRUgEJ8P+0N6tIdfQVOg1TcoDrG/87xv0Q42vL4Oz6ZlX443ualyYIJ7ETnzzVY3chGTENy
i0q4+RcNhQGYawYa9p6bk9Qmhxwec68dLYMFhAuFensnCMcA3f3BttxT7SpicO9lkcg+n/tmKY/L
xGLq4jaJsIHJRWP06lyMWhbGjZdzUn3F0trh5Zpp1w2DiyGP7D2RlZ8AGTLBiwirC71vZ6TwYm8X
d5VIqozV86V/BTbDnL7mANRRiMAILU8uyJk0CCq+GFJB2umGLTm8SMKf/TfdvMYPwHkNYCY8rUqJ
NE8NtBF0P7NP2zIw5vunEcpqWHHevJ3a1rMIU8ywWWJQqMtEZaJ28UBIsYN8dk0eVlxyBmZwx7tX
rIL/8o2ts6G76uPRjcx/uZ3A5prUAGkeuV99CFBvq1i8+2mxWmNRUNoZavrpzzH+M7rxDqqWEzsW
cBmjCv8ixdaSWndJzTQ6mtvIVwZf6fOM+MZwV0Zs5wsRrKAF6+h8Ii2VSmYE5mVG+kOAvmFzhCMI
WJI1weNkupRX1PKH/Z9qskbwCxrx8NBfA0hBbCneK/IxNBdS3c53DV9LClbVILGC1wVCkjQJhmSx
Yc7uDYn8U9ISiLyAwPnCZLtZPPTvLpZZa43XDqr85+3lGZJqRApv2ZKwfkXalBIfHWzPJ1N7jcvm
JDkdBtP11ty+xe/sNn7WfI4tluOFq0RYMU6SCgxI544aN1Bpb7pRqW0mcVBqUHkVRBmxRNp0rSuR
7NHgn3G/kaN95BZVEnhRbBhHr3XGWHGiE1ihzAaEKBP02DBMPh3NeX333Wpz6NFjCAAPMCVJKd5N
KqlXHT9eSYMkuQP3ILbCuZ8zVhezCKXxdD2ccZjI/V3RuhSQHxd9f9iXuidfHwR93YEac38FIUhy
1b3Itvc/FtVQ0Q6sIkSw4cie6LNlf14nFaS+W7T87WNGHxIWV8tAABICv8obbo7LbV4+OeWJYBl4
3AZd2yH4aaOtFPaFLg/Mv3Eglm0O6AyxljF6eeQoZYaqfGQSOYeH280DWgKo4FQB+fPLy7qSugJz
af58qxk6gvFDCog+gcMAP8le2hXrFGy5ZfCzC7dRlD4LPwoZoz7fRhMxt1RQAjMmsg+D6sVAKqT1
AvOgoP+sizhQyvzXzgs4VMppYfxdgoVXsNPqNZasPwDT2TKKH3Fn4eAwQBSW/kZr/y4HNhipKc5X
4UL1DaCFph01uSzGYKvzhDZzBEwTfieVLEbN5uJ+N8m4m/Zc5D2ObR1u+odkDo+HuUUeHQ7kyqDJ
swMwywr+7Zqb6BImM4rVIWyZebFCL0uVRj4pKOEvVCBa/WSh6xtYCa077946dqZRJ9fh4KqslNNt
KjPqmyUfLHQc9yH8qfoY31P8gpI9g9HXKzzIxmh/N11dp37TnScnKRzQSyWiflh56EhFokj39Sua
dfD3Cf6MDBlCQ0K2dGudxb4SnfmsBYce9WG/xKh5JyjOQfky8KC3gPdtmd3sLUqvtghd1stOWmzn
az/PSOGKQU9e42K5rFl+Y7Gf7B5/Y1wAgxqpTsbpqZ0IY8dQxJirVZqHufkCu/5boYXCPZ30//KA
8/j2FUTUmf9H2uVHHYMhl058aRW5VyNhJWxgm5cS4enZp8vU//KR25q4Bc1dsRl1KqM0DoNr4Puh
hj4RfuiGjslEXwX7fQoV+B3g1AH7FM0FHsLzAcmeoUD8Ox/7cc4Y/sodThMncFfJ/VMhAMkhh1zu
5QhEzH8OxHIC1P325pXjdembSHSo5SGOuDbRa5ragggWwo0CYPLP+8N6HbKHgJJSwPN14XXGR0tv
gZKti5GTkKcHgimNf/jRYJ3l8fbh0NJLwCJ4ChXLPaTPUa8ViwiW/htN5aR6TFeyrZPJsFOlHYyW
FKVzUtZ+94uTdGwywsDCOdXq7gA0pi6bUlBNw3ef/U5PAVqZw1FASp1OYUsRBHPKz2zJcmZiuZB1
JMjI64RuPdl0BXOHz7iJhd68j7pu8ENn6gPyab4Hm9uG0ayvOo09gGrDjIsIf98xtPxlkwzaOMEZ
dj9s3U9Z1Exzt8TZYIp2sBOtdvKOLHRt/tJEwIKuCTx0KpNkD+O1Sf3A72psB0oDPDicaIu4vmuI
QfBg/ORiIsUI8Wz2jpRceXZ4A7MenW3q04dOA7W+alm0JBLJVgsyxOE1BxKi8iak1l3aYHeI5KTs
9smNr/X5LYrwoKGZAs2b0V0LX2KHrq2yBpF+REH0yPU/AeU9pCMdTmZinJfxvcZzVhJyePtaSdJu
HPlRYMME9xPAwU8nR3XWXWxwaeoOQ/bQKq2PXPFl/jgAKH8F8MD5dsvjwvFQF95Z0wzV6yg8AKSG
Gt7doDB+rJGWxMts+Dw7X0UXxIzKrZP14XeZ5cNKXDaa3zSunUH20IyzCDjSABBtJx2c26BSl1sZ
jndVO5Y1BEVmkgJa4RCL/nufDJq2T8ODys9nxaUycCrHPDgYWG/+1WA37h6gxe8IZbCDEStCPPi4
1+rZL7zCBVk8ETnWzGGb1RmUsLYmPT5f0dHI9Hf2w0tGPoKC9/wN4DoI4dA7V6sczJ9CTpE1J3lO
5GAAt4R8j3H8If0afQ1rLiBahgVVIToyLjOUUo/G18RCwjbRsv06cDhmrwUX2mnLrVX3kBB4uUyP
DYW0O0guQCorNeLNGNjQFwLwiKVFww7v4JrN2rm5ndrF1zT5JS5nGUAY5LfpHaTBE3/0tGwexEY7
/l0OvIPLp+BGYZUK4R0MB21o/mF2ysuQ23ABwtw8YZsrk7VRLSzriqumx1a6biIt6oDLGJDslwUS
uXSvnEMZJDsDScqIM3ZutRxdM7zsmymyVlfRB2Ido/+IOpHX5S3COr7m/Ttqj/S3Fbg86fF8eIht
BHYafuGxMIIK2qNPYc++0NFygZszXJKtxRGGMwcPbFEHN7wbRUNvF9RABZsSmzcL8CBamS4RLWJy
zgZX9H0wz9ovH5l+HZHgqiC/m3MPH8eB9L7T0jdg1l2I0DEOm2BHT/IHnMQv6JBvWkcf8aBowGgL
1QCwAjL/7S5B7d5E6W4GMymNKikFOJhRS4qX8bLg6kD0UC+vR+U+o1wc+SQTD73/NCGYceFlq/EF
fNRpnvNzBbJ5qxXnU21xWSLMubhAgt3xYDzIeBoelFiH8qXo25M2Ng6oUBsfdY3Vys1ZpCYfqWLv
DlfJHwe6odhlMPjxuj1frrTzVsDaPVK3oBVJpSBcneSZyjiXIniIjM+iGtlV46+lI4JvBMZChbBo
EWXzlVfby1jUvSOwNAXrENvo+QY2NMsZpDtD8Ho2MztjZ96pi9f9gp+akAimszlDnT3yyAsKU6dT
fnL1n108Xr8xyUTjD5kygqyqcPo4fN/k/Tms1r4KuJOxkWjFdq8Ugg/pCXta/sZyxytlE+jFiD+U
4ii5RFL2SU1Kb0w1XNoyAQzwP0AaoEpoKHIfa+zN2kmz1OTq3xOEshGwRo4R9J7tE8rjZUPo38RV
D85vWAGbe1Aq450pE+9BUAbMxaCTgDvIr1SWRGgxeA9IAqawrTTIHWaizm9rcAd03m7H3svJWC0L
dv/0+B5KlAJhBEPQRtbR9aCYCK1+ZbHrwd7qqbbZlcOgvlCbWdeDZvqRjZjwviu9s6XRtgC7kpRG
RU4xwYcv0Smike6QT183KCKsxIRC9vKeq/KD5WpU2vcfprBhpqNRrUaje4zs3Rn0J7KcBns1aCwL
Ue0J0PrkI+G6Eeo00J8rl9aAESnEWpjBovSJiuRUENz+TXf5lQDq5UnmdIhMP4Gr0RHNkLrG+vWV
RyjDWl8+v2HFljaUfBKyv9bOQyvR1eh/oU4S+zfJ6Yyivn6h4//2XAXGYqWAouS6aGdoR8mXMBsN
/pfsxGdhv2J7nNtAmYA216zNKUQLVu2akYazb4CUfB/ud+liaKup8dkFyCdu4Gf6cNeRUuw26z7y
GV6dM7VlGhiAa/XLtOMTvyJmjT8uObFa/tZZApXRgJVb0axOSi+tgt+W1T6lOe9u+c3xZemqga16
49920lG5raEIduGvpMCLT99U59lBrfJsIG+bTf1Y+hl6w98/H9nioAUTszfSvpVKw/R3APvATV3D
+AmJ5NRgOOVabWb13OR7n1P388EjFCtx8ApELMwz30vLNxFEBtFsBRTmyY8Wy8GOqUl4uTvqysN8
56BCckrktBVQO3fxeMRQJCR9jR34as0+VAw/78U0N+AWqKo9AIF/rUZV724q89daJD8WUv/k14Bo
2XRZs0Nlo/RLlKVkFG+fLfPEP9I9a4ZxojA75dTdvQhhApGta2ciO49YVYD4stgo21UOFliSHFEs
V013JeavxngL+IgTSYkJ55/DL+NFdmCS7kIyy5biOZ7TLpbrYEHXP0EpBj1b2bJ9wdUK413BrXfg
6m/s7CbmtCKSIIURdglqKcA2p+AlRt8eXTUGOwYHJqAz1UnlKjP33ZeHzbGTIyVT8TOdzqDUjpLh
vlqcKFhVxxB8FC77nIh+WzXNY3kiKDFXevQPy25i3dv8dna7Wmgj0FWiYZAuxexQJvcvqEDn0lUI
AM4ZvGB17jw/AZS0qvnH5PVg/ZwJgzP4L3MbZKEmXg8ATA21mWKkubtpgks9Fmc6vZUO6pGPWZ++
mwlAeJyrrzzE+F8fl7iiHtrfToBdkPl8gixkPhpxKYWyne9TUyV6M7ds6/uCdmrHcdr5+szVi7m0
CUVaHarDMqEXAySpQU+Ekr9wwDOmMvDFiWZ7DXh1m2nDYqTxuS9K86kSLO0S0KfsnY83qF4KuH2Y
0FCt/otYueVDMhsZTt6m/XhcxDNiA3t1xlEE73L+TF2og6X00v6M0Y3E/xuS62Ie3DhZXeQGxhpf
H1GcXzFzUfsJLVeOpfz+aL9p1HBMhuv+AA65/LJlQEb/Un40r8iU/CT5HHG5N58g0J4b2N1pErUB
9k+ZJTWK9bGd1t0egrFkhKfqdXzWejG3n6hMw9r//BDZbx13SLhd+UMxr/K+Vbg3yk6ruEobGOgl
KGPSniRBwCVjLviAFCy+htpFR2Jn9aWFdStHn30fzCpwteGQfb2j4zd0yC7CDjG5tNQVsYe3VE/0
Qj60Cpudv4w7ZQAIaDA3tMPN+dLszT7FPMfNeKMTqXIlzpMzF7290Sf7+le/McxzcsvBbyprDDpe
6VPXNKEtIE6oJvvkTibCO0oyBN7PduZVPPM4tZW4Bi4BQJWGVLFp7nh1wbIca5+Cy0m3+653IHKh
kSv/As0sS7hWmdANphbwZzSLpb3TzlxaKNz7Um8oYaiUFP/uqpQEL8gAKE1wwiy7ryPdlztHjnSl
KPq3Qk1Oiodq37D1hZgo/pHmN8T+Dht1jmUgNc4FTKmgfAYYIXgJQtxcCxf+0R25wW7SAsn0pThW
VvcLQCkLo5dcTHL0ZQzy6DRZe9xvKCMXCv6/NLbdXuudaPQs9VK9YdBumSxBmBzvvqsfYRgh+pVG
mTi65de7CcZNidIdYouSGuEt1Q0Y2Pw268sVqwPQGGE3phKX3kWA72r4wDQ1ItmQOT52eZxatIkM
JIpiJzai9xdjCkzSNLrh/5PvFTJge19Edk8VnhKonUBxc3QsuGbfqh0U/U3aEkRE9fUuBdZYYUma
ZsmXBw9I0gHh+yeZZ23KpH8Kn9R7/ODUcdEwDX7/RQ2QgiOS5gfWfZg/GP4Uj3D64XPEOzPzE/MS
ea4NWGsUycR3Wk8jyaEUVWotge+Vur83toWh2kcDkqKY69OW+MfWdKTFe7/63BiDidKNA35LP4Iv
Z8wVuir9AHaUA8Mk2Vhe7C85M1ar8JwxnXeseN5ZP4ziJwmJcVsSXamNNl0geVmWTiVJ+BBrpfTe
jZt27nH07HQ5YB60SFtI1dSMW4ur1l8b9nxtp7D7C7tSt4I7Vuw5mYGXEFzT/09PMqmKnF9T0Tc/
SIGV00TFpzEw7hlOOUsxrSY3LCcXdXQhAQrMG5Sk0a37bLzVY52BcDYmNZLGr6/w61zXW3GUo+3s
okKE85MSWn7xmS7AujnyH/otT07tdUCYcbQzMcrBBC6dfnonNsZ4yFdyreUXlMPzzldzSfrlgai6
1ng+a8kXsMbfe6nP0MTncdwLpuvYFnj2XHVkUuiqy5havhiDI3Syjw2whiVAnaodt9t7D5urRgdH
J18MhiJXEgzKgx9dpVmZW0n/XLhV2i0WRrr/bTvYyd5lXq0tRVbB9Kf3dT2sex+lZVhOTvTkFFEH
0vBqdba36MwzRNGyJrONwsqS24cPto6C9rGaE26NJPlYLfCZU4jy7Y4U+wyjQOq9zdRZSzyHYSV+
sg5zbMHYg60sbO+mesmHHRDlrpEhjiHBObQVDxdjQkbaDRlZN7+ixx1iS8PydxXQNSRla5NwHOor
9Z18LAeLSkq4ra/mXJCGTL7lKhzS7cAZIqSeJiUERqVOENCmrdRDxNcDqN+fHNgFqhG/wNVdGQsy
4cbF0DiJpszeS9Viptt3jKj8WE331lKbN6BMADga75QXk+sDoPss+acWcpTUrFwQdATRyyi3pkRI
QXXbG67dJJtOX0PR5TOL1EQVWILy8ejEjzQMoWswEP6u2YZXS466isSc+L6ucN9egf0ui8Kl+/MO
XUkLsMO4PuPT3eHBgQc7aIMTHU6HEdEtOAHucJWZ9K2zFW3jk8r/9D8mDxsBNkcwu665ZB+nbk1B
LiIXWHqfV4P+I4cIQcQh+N5apz8tw90hejQPwwvRhLXBgbgK2r3GTQp8+qPFPXzAhFceLim+1ZtT
VVExtwB2FleAhisiWE+X+Hnf9bnASDtqy2VOeWR7CwsNeFVLRyjYMoX/i2md/BacRLafoyGvqvbq
11UNKdd/2J3WVj0T3SW5mKvhIGwGWbChpdZvFEHLZRmpBsZtxkHCG3mmFhet+V4rJ484lQ8MSPnT
VQEd1O4GZHX3C18KJ1lEcwe8te/oz+j10umIJu4ZU/GZ+kenCnfoW0uaERYip2L6W3jsgU85DH+h
l5YPHk3iPdsBvDEtmCBN7273VWOlKrRJJuqSRI+W5pEGyTWdgVqC+LRVtNBuyJ3kMsVrz3hTQUtv
ZSJy1QTe5ybJsmpd9B4iE0Y7wDhkhaifHLMYSUfn8OPrk7dOOnmjC6JQbK2T+unOVtDKB7XvJNyz
j7Yim0H9XyPqmm4aEWapdZUzf2OUftGhG3tiowMreMsFtkfcyyomETvyemr6FBUocQ7fzo9CudvC
Ps7RcSRxnjmtVKQwl42N66eHJLlmSYjH0VAF3zxolJJmAmFdbMUpR2pN6JaXFb2EzUdFzv+voHDe
PDejPKPYiXqzcjtHm3Pyl0N2ZfQbX/WUHMglTSjCm6xeBT41Yjg1h1rcMvmwpvyt+BnzUBIka5/S
2X3RZr4ruWdvapjEV4qpUt4IqtAt9aESsugslXCcm2EX4C9XnlbEflzAXJYhr8rySyU0d5mvCypG
2HN0VUL3/Us/RTBUXKvn37Wik4nxahO/7HoM9VRHn419inyGDdUMuCzydghL2Bbbe2xWB0/Ki+NJ
uCKiFiEpk5M43ZZ7f/PDzB9QkdsXd6JaW4qCCIVhAHBeYX9BnbzK61q6t87dk83/AvW3XoD/aVXu
FHjc18bnvJIaQk/pwlkqEQjLEYGDAkdqlC27FYi9l3GdNE72qoqNs8L/uZFfRX4WKhg3j5xO6n12
UOYQ7nxp+vEdJVCui3qb7goUayrDsMvul7zhzORYHKYfDo0ng4vK21Q3lHW/hRnJGi01Z2gcb/4t
EM4S+8NAJNfAPVmnAHfz7q3+Jitq2KHEbB9JZOzKtepXytRMVv95as3XbxagI1ycw/K9FobaiVve
uA1SiB58S+UxiuZUTAxf48wVW9hf+jLkLAeNNIM/gapfdmf6HG6LkjAYG564ILfPwL5qtf57QbOu
Byt8KRJaSb1HEZgfWhW87CxiNamQrCWtFcbHy0WfWCaWeVQoa0cwGtuihofzqOSXtkQOkqpplmzb
WvElkqrRLQRgkYCu3ppbwpr7v0lUCKrXlZPcAxemr0dz5uXwa7ktooy7tzuIBlwgO4xTlqTSojgc
XStV7W/2l053a1s4TN/HCjdTLCE3CIVuWdx55Pt0gaFp9NgJcRDW2gRJjZoemPJXOeaHVFW9JiEf
zaHiTeKLLvbRc0F4RCxwddpyJ+UtrSRCC8OWLQ/S/Gz1Nkb/OXrOiEoHM9ZMYyEMvVeBh8dsC5UO
dh/iK4tvMcm0Dn7V6DUdnTDKuoASCXs8tiWmuGycZJ3OcXNaNbRUwPUgHVnoi4rSG/B4wb7LrmUj
YIUZfdgADxpw3ttNHlUed5+1chujr7oad9r7fNHClI43fS84xQyPJmR2cBJKsiGrZspzXqMyrNvO
tkG9KA/flKA4f9k+RvkPeOmOGcP9OE1o/NUTSfgVoYKwMbTrTiyA9AvwouU/gv8zKnGa0T9NMEIX
2jBXr0Y98sp39G1Mr9tI86fwkXc2mPVo1f8gGHpp83AvBqOjdbQwdWYmM4k8/V7bpUpJCDL+fd6f
yqaZ6Njl+RueQimzuJNnq0CMyeIG9MpKZ2jGrzSyctbbN+wKuX0gF8CN1Aam5y1O+mzJhzPtIfqb
r6RD3xHvC3lBsyJ81Yko2K1AkqQSMoY+/JhaqDm6lprG/9IWoG650VFbwZszovvA6SAk2Fj7pe3n
L5ji8ZW2DN63LG1dYKw9xzeHkaK1Sv0LosMX+o10y4QHYBWuILUq/vhn4e2Je3hYrzaUS+SzxWoB
gpzMEC3VkPu2+5uOyo4cRAGzNtZvaRuuVVgUHG/pFfkBqiP44PwX5QtIoNxRyoVx6bW9cPT9lNPX
tALtAiHLg/vd0+YfAtnIH4U1MWyjMQrD8gGhq2snuKHi96Sfkce5p4ZDEJnVKdKlELqhudqexiia
3zroqpWSYxpnBkQ6tEGYtrtVzSJ+YgNcxQOJVFuhFRqqM7c2CUIJz5l+JOzBk3vT3MvhZNVo8xBC
d7+TT9f/MU6ZJfAyGFDsU+FICp0JwOdZZ7Dr25h1bqr1vsdrl7Knv2gVc2RW2Nzd833eshUDl1XB
5X6koAgc5SBR1o8grevkKwCMEcLsI4LPGkYn9vJFkccuVMlK0M6eW98xAUXEbWoH1rXaxmY0VhYK
mcogeL0FpX1byyCbl/qabqFCs3gFjQiBvzpbox8TJsQ3bVcefCKOSS6OMib3a16jr22KqVe2F3h2
7PcvYNn/s7j/bTkDCItjSapRNkdogX3ZHpIQffn6bRBh4tEPqm5BhCnnrdgVHF/oxjnkEXgDBTAO
amUcq3SFDG0YDX0NaORZYqGC/aTPIuHFny2hZMpls5br0rMBlHBcnXEADqe/3FAEuPE69amEVeam
hnGBJsvcu7w/4zmEmzEQVjd9w5/0tr8meGJjDJjpnTJaobnega3uK4Xp1wLWtvy8ofOTrmxNFGrp
nP3KT5yzEzmV2Yn/M2xDeBUfB5JiUgJcGHWFpvvfeyAOT3y6ncUkXHmlN9mzhW0DJ8ZfFRKbQqcQ
T+H14750FffzJ6auQ53wWLY4UukwkQWYV0J5BVlG50OEbKh4yDB7LI0pkp3pB4SdfGwUunCq1VB1
HWwYTsfS297eBrWlEjZwHIrhFC77aw2I8fQlrZ5Vzx3mCxBj85gY4kY5aT5+5pDHmGpEPuAmS2V9
kWt+q6CX1aMDi+NbKG+j2MsQnGZDHr3flJL7LUrtfvFpYpcuk3RicW9kXjl8JLLUQC7GuRDDvuKb
A7eipM9YkecRcqH6pCUFtURD0uhqlwG6kwRzHVljMV572w6XUbjDGuzJlmtxJADxV28QCgRUIdAc
U5QoOgEwWKIvPNBR2TXDzXgCRsMaXbATUnD0Bs7rpug3J3fCa0Cfe2Am3BymsSJkZWvevQqJFG69
DoFIbTKyistfbYg7ES3/ZOxFORs2C3kPNRjim2rMztuffsEvBL3r5yHXybFxsDkXen/z9JcnsrJy
0u6SWVBYT+seoDUdj/8aGzZBVB6B/uftjqIVlnaGb7w1zDbwA0XCAa7+WYiYTZtu/Lvb4DCOjrqw
4BfRFrntVO+UiWIDuivNsss+O56dX/uW7/xV2aj7uFW1hlMxdjZuRUcPjdS51dikGSELXbx7zYoX
6k3r9Mc9l43uqxA5h9xqDszeXAd/7U9LRv3MVInInZGNdZyi4ibx5Og4HBKidtII2FiloMFddsTZ
9YQmICG4NN1fgyfZ8JCa7knsH7HCzbD9qJNX06izv9oCcv2FvJcs3jFbez/sNXdDGmtf0AFM6DNa
zyBajFJdHYnMW+38H6FSi3jsewwttDgqvNZbamIrfYE4dJan5QmpfqDN89MnODR2Wcg89LIajL9Y
gyed2YFYbAaRgYM1AlUEMoTHyV88g3JMa1E20nsLwG8d2UoKj6qHLsQfDQ6jiMG2UogdibnFIOIe
jM6/IS/NVk5Cw1OG5/HtC45exIw4p8YCJN5z22/E4dMz8f72jiRnUf/3FN0Cd2fS5ge3tX5G52Pg
KSTME9saCpRK1GT+Vd9U9YaZfTdr0RLePICnYh+qgLUHyS6RZ9PHtChHUJ8jnJJpgK+AYdsC41s4
hB6u1zLe0pxUQDy9pPhxjssxiQN2mrRmnFs34uNiHW12HyXa9/w/QclUjjrczPEvDKQgUUfsjvWV
ZN+DcO0NqtC7v2huEQD+so6GjBly0Iq1UK+muI+lj9GzEZb0L+wyA7WS19+mVE4kjOkZD/Fwo3M7
DjCLhtNLRzl3ZOXJm4ETP6SVhtq0RfyPLvooixqXpKaEmTM8UP4d+QOo6lPnHfjFelZxPGmyWCYb
BJtZ7o2ogc/3Pbwm5qZjIZyUSX/qOT/957Phzek1YEAaw3oIzMkgy7EJRlUgDKv3eLnKsSTeBj+6
WXB/bDuVqeI5l9ncoOSYdC9NDnV7OwFlKwm29vQErhZQl46oXzZGj40ji7gUZOY/dvXlxAp8nC3C
MXNo/lUWHfuH9kv9IssXSn8bRWB6ji0J9uZn+aHTRSjHc5KpBHtdtNL5Oom4TicMQ9Pqsk+Y3+Yl
EYaCeJFjR2tcEY2fXXB6XiZbLdMwBd+vPrY6U1MMcxz9J/rLJ3UFlF45SUkAeKQEJWiLKoeqFP03
aLxag+A3CcM2DWxKTgrvRU7wRvQYWYx29K2rUPlgjmMdQ2jv9Vebak9EEZ+koTmfBOE8S/3dr3Ee
Qyx0MkIaDeShRPi4VhEPVLnAZS5fgvpszIeASLUQLGQMcmdj1cMJlalPfzhymv0R1uayGctjfo6F
yMOR80R4QamcxgIfaEFRtlBHBlDFEGBaCLtwY9AxjeaWrFhpUqd9Kzx5afPR85F8YoAjNNf3hNpf
V5JDp8RAUVspHZXurdSohhbgVo4xCBDa4C6tVmSx5IilXjyjgSz0SSCIxxzL59bDpbrA7amhl++y
8V9qDgVzFlqDDY1bLtqef6hCZfTJAa1W14vGSjPYBZMyTfoG5lpCjMgc/8y78iMBo0p248pnQr+7
qKe8DhBb6JVtZmfyO3UGPz6ykYejnsBXQVMg9INT99MfhkmOmjniQUl43QzujUn/v7EgRLwxM6O1
OLI5ZEy5zT3ITz5AEqzDRPQ2lCarvcTHEHl9/zK0PzEF9V3pZN7QA5Gk4hYYWx8zLPMWFTMTWEcz
lQQf16lCyzsHkFk+gjgHYZ1W2mu6oJaJW85dxKM6yTkUR5lamoO2D9hDYm9DjiSEGx/MPj0a6gLT
ugipGmVErauaLrJI0Pv+GCN3psr37Jmoz8P4PRqZ+UIvOQrOuBHhqeZVOUK9mGS8/ldCXXnVW+xM
fQHGsb6j58FiSvMoCoayKm3iP7lfNsIg8ziPWRY3gU54fMHRthbbCcpa0RSiloDtIqIuBKN04HMK
0oLsxvcwI6C2amu0GsF+ZsILLQXhubIYQQ/VR5vrqb0XVpSjP02gId+Aujx7JTlcoS+GgaM4CM1H
ltZULCfW2uSlUPJjZBRooejHRddOItSq2T1YUDGKbn0nkLNW0cZe9aFxVDghcxkGoytx+1Cg19YB
C3uZpglXoMKiwKihp1k7ZYtyC/F3ARDJO7mxpFIoGO77pEz07g871Eg6gvxZ79eRJJasRkdQE1vI
HiLT/qb9FVvKkBEksVHXFAhy5Iy/ZTz/iYqIcVDu1Y0RCmPzlipJiO9HxPAP9EJHH1Iq8ty9NWVU
1ffVrwpdIv+Ue13+QLKkdTpYcSdK7PwX8AOPfNs0H7A8gpY8ja9f+H+psbAK//mUFnEraMg4GrMo
rvbIGFh0E+nGLyF3qGsC6rpeZgfkYwOI6DHifw8dxdCKUFUX/yeLQSMG1YT5E36CL638fB+LZumB
qFBUSHcya+AXXpfPcOB32U2ulyPhlm/vxSMPLO/HIdJfttn2jTmp/+JATiLSsijJwfJlWJRnQQpN
FFgCHRGkoqT5L3H6lM53fE5nUbHlCmGcB58m8GCq2SM3xOzr4pnkpCV4MofORqow1z4jhq6aP3Wm
fPjw3BdAnHIkZIaaLuhgcyH3MlU7Q5Z9c2nzLDba7IykqiJL4rtsn08vKaGL6dC+yhdOdKILhA8P
U3JMeJtbcLPFzl8E6RYLuwcTcQBba80hXg0r0i33fvwOn+sUQytrmPCGSI+ADAit1txkb4w80W+B
1FLwoZizdWfQZXOdCxQoK4tYJwWlzk+yafdpPrKNEtfcwXyIH9maVX9G1UaucOjH7oIOBz/N+Ao5
V4zqShzRJdRTGky3bjlV8BoeKaG7SBaq9S3YAn8go7ojGNLFJkfzAYBIDrx/mxkU8qKfEmKWFF4l
ogn6KvA/Pp0o84z/NHBy8qbbksacQdx3NQvivanHlFIfkHkpFx04nBYPxkFBi8CS7wLcmDzBrmh8
YukPdScj58S7qUI2G0H454eqG68x1CLUMF09U373/7pH0mtgo9bfOhfq3sj6JJpQC4mySsPx+EAD
1RD0K2JEVQR9SFGUkla2mH2stCg2VllNVJPKM53SRVWwafmsddxQPM55vMnGFzfMt91Sh4SpfdDv
vTNVdDzaGv6aVT4oLa0p5b8Fwtki9hZ+l8HBQL0lWVea0zuKIIKoLmhtv8o4IbI7yhotYvjwRZ0U
Y4yZNxOsnTPN7wGP5fObdK1pzhpU83qlHEPx2r3iy2DPq+ZJZWIY/egjK62jiRplG6SBnhxoh6b7
RHGDXcPuaX/YkBQmoYYdl9BB6XcJb1E6UteYZQUBahAZ6I52OSshwJSFbkp33yCXXyeAbrYlUf4N
eoZ5hi608WnttKtN21LfoF++s+DE7VNlD2pU7qLWN6c5Qdv84KQNDegPimxyJGqlhU+yyQ0lOzpS
YM57ZqOgdwdR+aPq6UN/rUD+Ld+lUF1MWJOi15arJDZWhGInh41de4vkBSoNZcMJB/gBBTCZhwrk
5vOyumMUBcARnRxqCYLlcUxI/F9kCvfcU5vZ+2jNZVVbvawTHnL3864tcnteTBwgwcTzEPpkmJkR
Q1A9kfiWy4Z0IRgKHWtIjDaHxq6karWz1vBw3gwd2BqaAHseZKvYeWn12Ns7FiTptGfF/Elgzl7m
/2cXNzDXHWFn6OlzaSbq2yFvgMeUab/lajIN6inmSyWyHvjbzTXB5nJ5mSjxDD2HT1shgivTFt8u
J8HjG5Ruvo2CM3yDGj91pCL3Oo/Fddt6Q8HfI0QTofOQfurxwZPzBXiMy+Ye9ii1L6C+oGimi9O4
suQxM3u8mGIL8Zt6DzN0Gmpx/zuezk9JUdLLqDvc2HjqdIW6OmH3k8bd4T1aC9FH9EA+OrcG8WbB
UACG+ezhIwuKaZFBzWmeYCcIGBxk2PoYg72YIZGMV+Ljpsqa4YFRdWzWerm8VHqKNe9VKSCr9T2c
FKN9CF3jlp67Dyf5c9yBV5ReAQPj6sTabyJkKMQ5SlzmdHRxca8iI+OoMHQ3SH2z4y3ViMH+Spqs
huHy9GyHoF+YLKccjttZE0MZ8Rn3T8iR8P4bGTBZw1JV8CBzdCRtbm0EBv5YzynFtNgCKtSo5GKS
P6q5X6UsHEqYKHhlOoA4/07NDUD3Z9NunlEVzqvYcEhpi0A8UlGd4NMB5AGf1ZhqUWAxyzClckmn
l5emrQPwsicrxSvXm1Xh0m7M6dd/V8Y1kFvbHw6NOjY+5jbgz0LdELYxFUvUtN7MdXP+/3S7UiOI
FfQuxxUf+Wh0OPZxFVEmN1MsEgxvL6TAuXuB6dU3+PkRcWSf+9gQePBb1AfKu7uCr04iDNLNjXr1
q9u6ZZBzOHcqaodu4mzwhu9pHKGEqOIN3GuaL2GCCw44Hd99H6o0fUS6OGVGyWdAlE8H4PrtHYbd
Xkg3oww/2UAsIwUDnhaj4BMSdxn41//RSadY8Um9vRZvpl/vIuIRvgkjgh6ahwJV+afwF5enKbnW
++hdmE6KZy0s7SXSToAzgyDeruiiOFPNDigf6U4P1mCvxOoQ5tK7Rz8hluM6yB1GjmvAjHUS5JHh
sKcTnS/6D3Yczdy3qPK1pjPmpBltEmJtMYdIGK4Vh+fZ9iXLbAiCF9BkcsedhlQOuj5Dr3dTzSse
RfHri1dLO6LMmT57/fohdO5UgNJmjVRvWms1wexBQd5f5De/oGBdRhJ/ZTtf06LoDzj3yhPrq+13
V8PTDBVpaLF4cdWaXXw3+zweVucz2YW0gEj2oCBiIQgdcqUwLZwXdDwLF4A6r0PY027Nxrl0nZBM
+zgPRN24Sokh94WIFZw8i3yret7Dov/n0YbUkct25Pkgy5Yee594JGralkYT9nIpDET1DPod027Y
tVDIC31WDuaDD8xZO+gZMKJN3GOTNo1j7FBTkhYuSYRKYTRBs8qJYNEB1Qm7KPm5OQFjeI5Z9Hs1
hs3O9/RvfF8fKw65b+kCUJhJ21qIrzQmhq3px/ySdZs9bZvUTmRZxRzZBPWFoh/USNO3qAw6vzb9
KKlfFWG62DhEQxQ+4X8GX6tXX5emRCs2Wauk6/SE013lpuMnkyAqRw+uGWgjNmlBwG5MdXoGCJ8w
Yii8c/FD/kF1d2TJE3q/1OQ6/72aZxo0y1LXepSeLpc4QXVyx9XmLnCO71shhPMog7UIOx/j+BUr
TLt8fX/SpxR86cEo0tl6kk4FOzfpvT5IX2+CWsyDfC3JGgmPQ6azdFtAipDnPTWJJuK1xIkOCrWU
xkPS5kIRNsl7xsXI2l6MwAq+op50HIgvktgdlRD5cbkuzD00CxLOyppIPbN2X/KHfRzZrkaMlM+P
0t7L0NC6Hv+czdrTR5bg8OnMWlAR5qgzue1DuE+I6ZTpoqmgZ7tvTlc1kMbPtpoHW6JQmL9a8t59
c3urvL4MeQqROCRHabFUbD50Tz7R7yhpu/2gpZ22Yb3AtpgCtz4BtFFSlMwkkw2uXvicTlE8rf8Q
OvZ45Ny6GnOkcqGAaObbNpS0yaBBDcGKz7hsjpFPUBjLXUvSkOxDff97nSCF2AyBEGTEk3VskWiS
MzVIouhYpCLlQzuowaeAVvHKLDJLR+RhHocJ3hG5FkMieuGp7jBGriXFhN5BBlzqJvQQLNEsHyxH
6u1ZXuPEkX8eFQnWt4IQ96Pc56hk1kmPDZBX93M1IEGnfFFEqFfKNzhG4l1ln+oTpa7tY8RLn9KS
pLcxIIKb0Zq2kjv/rJCQluRi93nQip0khsSpgw/H6ouSgYkq8ORNz/hLHEsujHECY7CMjnBUgSOw
0xREv9OK/PERk/AAVVdBzgmEjuSeW6HGcO2iAZAUIXcp5EFLGhHVKFeBz7LazgiZ9oCteSVU8RA7
yoBViYIIplBA1s91Zy8nRkLUcSGrzvsJD5/CFQ2sj+95XsGPyfkgVrmEeLZoAGhuPaV12UJiEUUm
hWrUnZRMclM+R3YA2ffzhZc1uQBmwGck7uX1MoRLl+5Ic4OgLTzrK4ZaGlfjSQddjzo1QilsEylI
g75Xh7JBmE7Qc9Dbp9UWBRJNEUNBD4lkKVMED24wsaCQhWzCsy4KxcF3f2kXJK25JyMx4yUpyJCh
r9xvJji9q5fF+Cv4bC0gY4ZMP1fWPKCC2BVJyAcJeLfyUq4oK7Dn2hjw+sXJHRGuX7t/iu/WmtnG
SzRmRxlJHyzGRPhxIsnTdxMqBGoRlLLOv7GUhorLM4EV89xZ0bOOb2Rl5i1+rmjHyvRndL43ZSsB
eyGGx/rl+SUfReoXte7kX96vr2EPtcrEjAyAOf3x5mHXTohLUOKz+bW3fCtAGC2MK/0B+oRpOKff
IJRFH/hwX9hIv63n5KfEjQchpoYBP4Mgj6j158VRB3pSLk/SnJMrleKLd5Owgk4b8TLe6kYokUHQ
T/6je5JJd6ONvP/q4+ms9FMdkS5jM/1KlkJXcf6dsPPR1d+huqhuOYQLUrtO3wjRUkk51RPxkMFZ
7l8F/tHb8IB/AWgI6h/MJqrosBUCQqLoI+HLEvGj3lZBCrgQv4vdULJ91746+PXhaJ55RGUcPHMv
FRmTbLSCX5LSSDdIfR1r2qQOG0ecYhXfh4TlhBOuu7omcxQ2eFcpAnMpiMZliGMTmfAFIrBBdN1v
wfyPqTPhMYJpWkzt3Runa8jAGyYCa0UvSFq3eYYpTedbuRpIsgXiJtej/AFljxj6epUL6sEgXFg2
lDPZv4y5Wk1mBvi17D7k6ccpS9WaUhqfOEqa1/WXI8AjFAQCyLrR0CJwv9m2fQPFb6VH2AiNTuTd
yh5BbJTA4/5undSj7G8i7RQC2mrTIDWj840dTB8QG0Rsj6FlEnckYO7l+bwuA3auLCiQdTYs/uMx
sA25iH2SNzwQXjxQJXLeFxxMKezBWurM6CQl3Ew30pp8Kq8HCwp4QwvxF+r3/8/Br8ydXJvzSh2y
QA241vRynlMbSXPtdPg8z9nbe5UxA1qWkKd7MZjWzSr+VsMSA3p6LTobmmEv4j58Squmdrm3BXud
sgGTI0PeCF2mrWzY0PQ4SFc1pl1kHwfYnx1ZUcX1GRORBKCacHwsx0jVbwXJFY/qTIYBQK+O8aHe
5VRwN1c83A/LKSvf6qy6BgUro62xNmOwNS2E5borX8KclKFdwSFTmkBvU8gZBssfz/u6mzfVWMoo
tkGTbpAt8kG6rW2+hvaRXQi6L+ggRRgO4QEF+gPPU1koMVVjbO2MMyFtQPGYPGYLSdTFXZln2237
Hza0XlTgVwP0bRcWoAmqj5ZoljmhnQWCQtbD6NlPPkMR/91Ft7Yh/Qi50ORjiwR2xELLSOlYWTKs
yEiEKzA8Q4w1sju4t4ebvADH1ZMLV+c8FlDF369d0odt4hY0FgkZP5D8Yi1mmcws/hdjmGUpycgL
vm96MmmuV7R6RFd6xVSOpX8S1Kw4t3C4XI5BJbYkVeP0pPqQeuxB3w9eZLZ93MBnrG2jDGoFG/NN
MtXUjWkQDjm1nDCxr/eaD7CSJMUj8NUULDpyrbI8q6telfTupLlkSJ5KTIw3fD9mMfvQu9NgLnqJ
W9PbnChApflO70rw8z64W8iuTGYmZIOtjvNOEksDqayj86X/xfcBkHVr32LVKIazL3PNo/aixUpA
Q0sjbq1QK2L95d5CLXfxJS9FWntMbKQOCMuRQnuK6aynRVsiIwu6hQUY+IVlv4wHVjbJBnibXGME
qzNatfvJMM3dvwsv0mM4AZ4x1+H+oT2bGeG+CEdzkSuvpaOBXRv0OB0CGOk/C/W4weLdv7G61UTW
DoENLqIoMcUjSNqTPcPmLeSDa8GGH54KPr3g0s0PnU1XcuJvQ3xf8Qr6kkwQ3r/K6SG4Bdzewem0
8+uUahCCEqjgBhoFBTOteprYZJi5DkAMMh5ipOnX326qd4pMR0/O1SJBdOd8RLI2Fw4RImZ7na2u
82sPvlz97w2KQg5xjjP6oFcwoMhAQLfN/X4DrLDD4dRpAoVuM4wM40m9PvYYzB4rciVwTrSSRoh5
lJiIW2o8jVgg5EoZ2bWg0YsoByLtY/qzUQ5qFm8tw84zhVjOGRfyvqKPT/E6VW0/4cd5bgiz/RyP
XDdjmJIFl8rLJtA8PcUxeN3tPHjTtzxCxaD31PAety0NOG1FO7eD272mQSM9DKfhwpsFipR3LuSq
SRDDHkgYmfAMBFlkXbx0VJYZ1LXWpgvp7gl3Zk3ku9AxDSmZmHhRgMN7dwGqx8hKKN5kTiToNU/q
mktxeg38M6613u3QXzFJ+VEBpdRgTvcXDZVOTzhDwS8YIqaTN+Zqi84gc9+2MY+UbcdvhZAhp1EI
4HvERF7rP2eR7rMO08CkIDMsOviaETnSLzVyrisM6XIluaHkViAo7aZpOFXh/b8mgE5dyMyX5Wpq
cRRJqYZmuXZX/LDLqEpqieKcRhLX+f4XCqrHZbLDejuNM9zz0Okynk2Ku+oolm4903E8ieKPnuQC
34KQpAwwehON05YktHTw9vIYrR76m9Uhgh+kJ40Ukub58MMyLVLvKNrHcO+zai7mwzjvaZZhT8Fz
yD95Ohk0dGWUVQzUunysx3vnwydHr3f9Lm0CxZv0goylEte6FmqTYSRcNmlOdiUnb4LbuS+Su1jR
9C2pFbc1d8LnonPTnlZTD8QbVGZuG4oVaKm4+M2Y7UQNeyf+EFpi9kSZeufra9qcdoNGOJ7aqQxy
9a3CKhdrIXbtlkpDZ8U58+HJ/v5RXDoZs7vCuGKaDjYTdnJdM9BEROyEXGLYSo1zPQ30WYHI9vrD
i1jw0pASyRcpbHA8jDhC5Ie8x0S3K1j9trRdS/V/H9h3xA+fytsJQ6nZwXEnSbwFAj5fDhSFbZ8S
AT53NwookXMP0nYreOtgQzffMWzSBgzG2vMlIXsfSsFGJ/28tBH5lryzCas5/3L+icUWeW4OhS0m
VI37csZPtMCHVKojKdGAwb+E5RREsVXsdkpsz+VlAPoFWXon722OUPihWvdALrZ358CtVxFBBiFP
Ex6b9VGJcy//izLHa41+UgoJj1a93lpQIzDynhKlBLLWrQRgPLCw2GUYEANu6ugfAsj+nHAdWH9+
zNZIR3qrLkhFfqN8JbrqMMOhJ+Vw+Pv89lsOs9eNYrr/AGuYelEKoVoQDFTeI8SgI/jYs/nVrcwU
GaSGvWVok02LUscMRuNVmOzB2Ybp6ffK4XZUaMmmKLoneGNSneWHoRWB4MkbfdkFNJAohrDXKTSI
vaHeE1Xr/+NLbw+Sc4AmLiFliVKRJojJSYclJshNI3GaUsihdTsQWc9rC9LFvcxSj3DXxKG0OeXK
LcNyb1tVnjWUGeBIKvgZjfXoCWHN9xwWDmo+uCA3ESAYNpD2KApl2fnh0sh9RSKjU0QkjvosQNNF
PrGfscUyQ84GDwtjfSs4t6t7OgvwIM3xhQEWw9Hi+4PIYNUCDDEeg4RfcyUvghJGUC6WeuIZjR/R
6jDPAGPvqnxP+hdfzRleHPouCPxT2iLNr6DP4FDalX7GgNSeZ9gy/icdVmmH4ePpsBJRnx21CuJF
ZfFOMFUeELO4aKrs21aK8xS2VRMgfbWRzZWWrY+8Gk5HYl+BzsRwlNhNOg1oZ0e0Q18ze3vqEi3T
W0n6ixrcJu5ldprbFDT+ly2dfkActvZLkJIQ55juX4wuNtoqYHVwyJQGOqsHJNmvrPgu/u578i66
R3ZNLtkkS5z/4sU1VxuQWnVdBKTDFVfjIQwODSVdY1lyjXEN47obFdrzw/4uQjEuDz2Tcnm6e1Pi
aL0fxIrTlqZofaC5/WBlNGuOGkmDnDaIFerErpDhH6j+Chq62RSvGaSXzDFJ7jyAxV2kwob3SpEd
MFSfuNRIMAgKl/hYFfGnph9R522um5k8uSuzanOcmmH95+KD6+8z8rssoT77V3FH4IKHArKwsj8Y
n2d93HpY1zwlim057whxrsKd5U8YDyXcEoogA/wHbCyxpeQPxtCMKOY/Ys4A4pwju/osPZoyqTLk
ZMC26ME+HqLQLSG984VjbHflLNez7FESRPKkBs5C4H7A8/PfPI6lZerq12xsSCPhD7yixyjB0YA6
QHc34yUZZpiTCdNKIckgbMN9IUmj3kNo1KO2H+ybcLoPj1uUsSw0H9ByxQlpTkFWsj8/2z82SPX0
B4EGcU3bA48DgZa92HT58DV8KXDLaMHWmjGhhgvki3iNqx1sUlBSg/WZpY3GVfaWiMvbCdrqh5XU
MGdOo3rgQ2xW1iTBkRRySxtJbBHX16U5ts1lf7meJCOxkiSVAQRGKW5SW7yz8DqATnUWsK57fWaF
esUSDYqgLpkZ3lDKWWylsg/BX5Pb/V5jeoY/pI6t9EO+N5dYqF1HVIKlyvn/x4Sub30nBN4OpHFY
4uMK9m74VIIAl3LOG3EB44vdXFwYP2NOVSnMjkMJ18y/7WH2FpPuorSX0K1CvP4aut83pp0sWoAi
LKzRThvm5UkXXI3+TnKhxWDZ92kR5uBTU1rV4+0VwbiWLpKPmVQmJRyrC8uOk1UEggusF0KEFbpU
4/l8igPc4tDcUAvoZ+FjIhZy9KftGL/WgbODgXdTpB0XSFq5oxOb4gbYnnPJ00OJ8sWw4sui+21E
lw6iUzK1MoXluzhn5TZY/L07/m9q+VgyP5diYwmcxj6ICr/7Qpgd4HfRBYAqqRni2D8AaqnEuDBd
4CsIbFTtVWVb6PgKXLznU6Fpumo8odfb0i99SSoHgpOS4vpOeuv1Smk+R90Dx4bQpkrW55N6XNHn
pH0SsAXube+U3Ot4YxScWfnAMX655/mDaDEcYn+SasloYLFTTlCQEt8A/ELsq0gvE45asy65qrh4
N+AOwLBoQwzhxKJrXAJ3CyCwkicyYHetvjl/x5WWW09s7fbs8iHYdyf/e5p9YFeZ/LLwS53xMFC6
crfW/IC4XLekbLF5UmZRfSZjsaMlhVocXQEUCEsZ1YjifYUxTJqT67yjVZ+KfpFfkVtqS1wTgbrs
AUcqz2YvsY+v4Afzios86hSYmYWSUJlXM2M0ypwePkkDNezFCIReMUIXQ4S4V/MFhJkOFQLEFYKL
MCmTpOK7okjwDTQlr0G1iayGJ9u58mCVXpY3HZb8J6gt8F3hVnoKPjEHy35rnZSmYFNxPRkSHyjv
/KUEoeB0RCfs+bn7/eeVpIxEMWOSAaTmv0eXwwQpDVCiqhuGvb+4FRZ9gGy/js1cZratswor0E6N
Ma9kXI/Kx901pvJjDW1cKDe/vEzfuaJr/k6+zfsCFORE/R29cCEoV/lIltwr1PaRyCEeOsW2Uudd
wWeAfcC0veq9uoyZ1wuijqhzeIYXP87IM7jqMQAxgn028KIm/YmvZAkMxbnZv4sJ548wpC2608+S
2yTGNpat3+h3OOx8Uwf2irGXnGZMusEqsvzf1c+gmynGYlwD/r7AjyUs0ymNc5Kl6DGxeLUrxGZi
7TJcneRgcAj2Wmr4R+YGhRBKgjA0NfoAzGsWItMGntUiAEbJVQFMkAe+q8V/9MgZZAQykTSGYVba
wfuZh4qWc8FwcJqWcgOKyX1XxcL3z37DOhMlbwB5qLsHc9xx0O0fvNHCLLfm7WTvDbRWRskSy0cu
zCeBqWdaX/RHwEnGpboF1m5Ti+S7fnm4dwAMzNZnXcQ45YgKMHGQzZRmzkV+/LzovcZstiPRakW4
xWg5YfJNZoAjkThqu4NhN0c9A8RiYm/6z5Ix1RD/lO7nBJtTo9fPbBxLDcsX6Q+7qJmyHszkfbn7
34z11ZXJ5uCPLwWdTwFXx7bH4Cf+HPe0tX8J7z0pBUh4eAypPKabzFv2i12I1odBInC4/ROozzsC
iTRU65PXHS060TgZjSGEmh3FQ46G+kRluBKqO3Gzaniz8EqOxUSXUunmuBZa8Og/gfrj27zRTe2K
sQXTjxMWAzfimocho6z+4KgfMNBfTESv0lHOesEbcL7prollfTpAI9SsmfA6S+e54On8dgnpY5tE
6lY/2lbVhg0+6vzrEcKxA7Vqz89SMIRjM0HXcDE0Y8bNABXRScT08iRCQs7uMdawj9qsRvXEMmsP
h4GzLIZ7uSGPl3D2bXWSV9ZIWipc2JVSTmx6MQCLVXeqtLcqf5bFsYQmPQNJbJhVgeIbsFTKgC2U
9PiHHAOzsERIVPDXQCG5nJVsJarLMlzh3KoQ2EBVcoeh7YrCm7+EoOBRvfq3Dou7kVaIXC+8x+Ln
tojr66TCOdGCDwYSpmOkzW1CQc4rlJ7cUmrtMUk3NOKHv6PPmCf01zjI7yvTWS0HYfSoNMvCkUub
PjS4Pnvmk1G3vdRwRp1Wy2YqtFWL5KWqJmahR0fVQU9GMFVq9Vck3hkGJ9htnjqP2kNO8PyYwmWN
gIP+akGBdhe3ELIqj9h4cspxr5CzzfKV9E4WelihPcaOyP9savgmKUdAQVoQZmjc+GHyYGn2dhyv
2d6ULsyFC9LZJMsZjgXGOWX+PqkSrI+TpB5xwxfeVBvPHqO6FV6KDxOxEOi003yw6cfXvWpAAALc
aH8On+aiXOkUXd7F1zB/C74Uhwzn3FUZjQldMwWc83IloRjX5SOhG9gzLKMEHWuwY/muRp+DT38+
uit/TzqfGgm3Tp3HNCWbExevZ4dAyBM/RV/kNyMjDxgKbAKCNvzYaE4gHHecNwyO2C7flAhogRcB
Q9fp5e6P79VPQRSj6fJ2UY4UOKq60UVVUoXrCuncUmcGE0CrC//Slr4KZxtPok0PgyA0ksDYhZSR
0dkzL2thnyJZ0mgXHJX11pOj643JvQAD7+IQaMT/Lme76OuoYzaFMmrJlBhqax/l3NWjTahCJbIo
QQAui7cSG1GJ9DbMWaTS9BayNCl6uRNAAAZ4JMxjSpDIzo3u/GTbukwjta1iUmx4r/c8FdtxO+1m
JvCFnl8ZIrrVQVqY8Y7EDIbDnUTHUqTKo4/hBZQZw7SkW1IrxvpuviRaI1IVbLRX0TngLLfPgnW+
9WgNSwwBx1i8Vylt5TKVKvp6vD2vDna+x6SZ5E/sfFb3Cgv4OUTb2ItatCaMgaUYx0SRcvnq13Ty
sYsaV0bG+VA3t2LQ8Iwpb8avnfdZdRKIN0v+1/4JahBtoyGlsOTQEstyklPgszTme46PQGi5Rfms
qXY6+6QejT+QsS1gbVgLCby+HbmN1VCOvzgxCodHLYsrwUGKU/en40XLVHtAcTrD3fy/Xo2BG7V1
W+4FiiMXy3tI0O7C5XmdVLNPET18TTtGJAJEmuGRU/mxISgzA8Kzxt455Jkg78q3T83p+MkR/UkP
JaPKVJvOPEAOZ5aSMacr11HC/QCAq4QmFtNdxsGHBcnN5W9dquQoj6+6J1WGhykY/GYZG7iu2jfH
AW33kcaq3Ynerv+tz18xDleig9oAp4XqpzvUmeSIzq98AkeMZn1eJE3ONxPbgnHfDE8WR1KxcbgQ
XgzBQbqgQKewAavHUXdA8JDDgdzMCSMRLkG/lrxg5Uv/GFhzOhQxtleYHOJ6ZuljCEe+JHKRoNXe
2dbTtNXxv7gVlbFOB4jjx071HhmL6Rp4qHNDBohOUIPD8W1ihpzCNfyEYfpT3Dq9yFyEz1hR7fhu
9NvscThBLp8ANCPd8lUqM0LQTwIKjaLKjllEb6Ywaqeu1F89I1VkCPZGqCwcHQRmjc91IC8Qu6Wj
1F/8AsjioXFV1hT6qXIdGijcGwKSm0ddVtDuPYSZIHAkHnHhz7FYM+Saq1laSeMlhme7uJl65ODe
XJeDyfuAwhWv0eE41tHEUXsRXvHFB5xlTsMgcFt0Gt+3fi/UBLzwCyrXuwIXqkNOprLSQqkcA3th
cFcnAuUVA2YHp0OjLIOCnT4HA7eFGvXYmd572pOwcMz9T4DZTh6U0SmdlMCNpdmA+9eIodnDkOE6
sMH2u9mDve1yPXZXNZuLlpCYg4hpUB7Uy85y+cyDeQnwN+oEh/N4ufPv7rCE0tCdkg6tz0Lbwo01
+IFHEft1P6F9MKaLZ7VuylZYAQDVtap2H9VmXp4Xb6pfoG/rcsYo1D3Amlf5WuBONwTkGtx4wP0O
+jvsCwU9kmUuLczx+0uI+3XVDQ5wgWM9ZyyQ7fQx0WNHhovSg67ud6D06n8Ygde7/wCQHUN0UVaR
Sg61eG2U1Wda92fZIx9nVZhwi3tPQzGCys0VPmi7x//Ltg7DKfsvKqqxNHUQibXDajRDrz5eNdmG
H4wOwRHG+9JXUGoMIqdpR9Pdmf/zWJB0A+UMaYTbSRuwAhggHVNNLx1FarEzBu+qhKK267CEbOFO
D1X/IS3kGyOUxyzm0+4eVQr8qj0UgYSbIgRGG5CWEHAhaOGm6amKfxn/tx/h66628YgeHgxERCHP
1uxrwaXjdnxcCnxCs6+jkX6cXDP5TLEFrmprRb5xna+PYeInFQIsLZK9Ng1RhrVebh9iOvRV2gzX
MCkgdtZYMJBo0a7KzioqOLiPm4naZur8+YoY5U0aD24p98rpHBI1yzxsXk+eICIuNQJoDUiveUFR
r8z0vVum/C3IaQx/DLaFEzXRmbFNdIercoI2J9zo/3Nmytq0fCqsZvEwNRFZbyPzJK/BtgBLw+Nj
bffzMyLJvAshI3SWoawSiA8mgSYaDcAK3FOMLlApHgfLHtOa0KdRLqdTwkOpBlqeL9t23nMW4M/O
oj49/fmg3nQrsiuNxvEO/DT60MABXWXN7L3YNKODdvhqxzTHXXr/OODciLVUm/7DFTdIgFzllP8S
mLtLXomRhZ5q/GvoLi6215yN/eFK+cZDGcrJ3JnpUb/9VW+sIWF4iuMYA++5fn2sklE9Zl2UEXoz
DFaA99oB/zBJbe/d36LGEoomeJiNq6yjsDKOfSx2vZhgF/Uz5sSr6Nq0Ul3QbInmXp6HqmUBYeJ8
d3YS6qU79U6OK+29f3I3qpsRa1hEMR1D7y8LYWbp1joOXQt4uuCkeI0LQnPFBBQ2fnW4RpAOYWdr
b/mvlncsOYmuF+b7iy4fzhSnAz1DoviKttBc4y/9jogbn25GPXBDTogp1uoqTmNsZBqVSaVE+Xxz
4X+TtBWHFDbuJw8orWQS9rWSDU0S/5J3K6t8PGoosOVAskAbKK/w9xWaUL8fLcquHTExhVVZN7nN
HvBXqIwDNReiFB8hNgcuCBQK0troJljYOwT/JcWXNOrDYpx9dHPRV6hgeL0GP7O3E0M8aqLW9ijP
g9lwk1KQV/TDJ7EodhB0i3XSIvQq8TJWBRwFwwpvgT2Y52JMBHkIrl50HmKGhzQg+NtHWZhg0buN
e+CRg5UT0sXe4u/WcXD9lwVmiB2OEymMG26FKDEiHln4QH3JNb1NPV4crK4q64pA7+CEZbB1GukV
TXDX9NJbaNYNX4zyS7FBrQqvbqkx2FxZ6wqH8uJBaLdqklbJkDfYox8BoMSomXXn94VZKx1mYMWt
2APFMUpdAoSOTEnopxEUVs6Ox6ZZ+8HQQZEzJflzrjBt4BBOMr8mDjBFLnivrJ3PbOSaph+jiotG
rPuRWW2J1um18cIagx6hsewNJFY7jalWN+sFsgk/TJHVOe92XzTxpOC+p1Iztrs9USATBeTIdgTI
rvBmv4DrwV795/ljelIp+1daqVN+s5dW2rEoS4QCfaAzFT+xVFwcii/1Mk8YyYEeP+eYF1uMOPJc
deILTRJwXrWgW2DZf452/+25YDUCWRwxccb/d31j9vmQpeZXKIil8wlU9UHNkAefvuYUghXO53pC
C9q+VfmzRzKRN1U7HuyQS1sQS58Ra2ymvfvENNGw9064qbNL6t9jt6uN9Z+ksQsTho+BCc8e8Pni
CsMen3Vo9z/xtA18TG8Iop5iPDW7jUFEATk7n1lRSm9omVh1YUiByKeXSxGkkqgmTLuXr5U4KIue
0X8pwAjS39F7/2xB/rP7VBu6gGXnzrNteu1RT/CjLZKSJkK3+mw5igQ0vxi2VhH2GYX9xfHIddgD
dhegZ4B85zC6atV3xRZK97ujIePKEEqlYBxEZckZYQzFtKBJdnhEvEqesRLfgT/0fTAtJBlqYqQd
sCwjdhroil9J5TCLiJ/hdefWE68CuwI8JdNIGuJZTvRKLv5Izv/IuImPXeXuVSLZB603VfsVfFsZ
2yMpAEjQ95UuE84nWNUgS1hACyKLthQxeYO6wlG78Pt7my0ZXYcILg+2BHdEaS73MbiUGN0Z0LtU
8qwsZuja70ipkouhTotW9Rp1eIe452XUjfsq2NubYZlG6jJbfBH2yVbCLBdrD5hZoiYAdcLSLyAr
C+aLe5MA/2CL2sbQ2WdtWWZoQAihOc/0d9CSQ7tb0K2bQp6c0tKPT9mKY/hsE4VoNy7eFG81js7u
NewVNRHA/DWKNfuoGtf+qcxZ2g22iq/sAkiu/o5+VWDQyFCiPlp/rDuaQGqZGqq/rS5mQEl5D7rF
5bRRXEdTWs8ZD+RerXcTH1s2g9tfU8htSFXW2CHZvWpo8w76lxfFETHSuD/kUNCXAUPXizousvtV
YM0yu8WNdLLNrPhmumm0REU1V0EOvveI25PpKofzfchX/vGluWd9klJ2VWXOPK7PxlrTiTZlDhCs
GzAod+UwUQrJ26ouSI2Y9M3EWIMSldaQHiMXaeMEs2uBLPkpt9COjgU595RoN6oXAwK1pFWBglVx
N+C+2C/u2LvWVSsnfEWAs5sSyNcyGP/krhhLZJLV9KMxUUBDDxh9gmiitvtSXEwrLMbnYq841+eu
cGjID5TJMPhKKu4kRFHrtaFgOOZiHSVm5vcug4q1z5ujDX5Xu1p2bfO2En9XEZDyOv/zpFgHQQLR
zQJWgR/VYGWsGrRpDL+lyKBge2zRjp6iKlIOuNOHRbPFuNOUH3A2Qnkbssyl0+RwxoSuu9CXr8IO
6OxE9g5KG2QzYL1Ln6mTFbwH2bgm4Brcpw2FA896e8jIrRPMe0x6qEOlfxg9fwLAqza/i4nPaMCZ
Sv3ne3UnEBEt2EhWyukh1PsIayi08wmZSUVrXw5eagvdhaqtt+veUx1AwnUWEDE5RDC26fpoRksN
BFxVQ44CwvXciWjmczq94MMr0t2wEmsV2Ui6C2rbgu849AcOxQbOKn7fSKEVRtB1wt/cx3baoPwd
fHFRwCLBW0i7G0YQ47bXMgZK5edpoxqNrJ8vNvvoxiY4hpo64n+xs8bXsAvho9xabBBW/dWrm8rd
PrRQP9DlSwIkOEaCDNuxexkfGH7HoF7UzL38v99t3JZH3smwiDCbvn0vCRRccLEGx4+Z8o+oMR97
mLRvEZep1XaIpuMSYeMD4LyJ6xfNjcLqBfwIo7a/RYkKxgZHRUDOJYMAhMgXwEckuKnRcvqx8FQt
qaUsShRzcVKrfej5Khm+pkvpNKT1mSjH+8wkMgCFR06z8l9WvalOhZQEJyTZbFK1Z3bjTNgwyVQI
fhhCxtZovKTnPfByqHCp89a9ZFP6OhJLc03omZLUyeucZCFJtWMyGY+2aXJ6mFa6npzdZwQ+gbpR
1FtFVMaHbZHttCaWLUF+WirMeaxML1A93uMG65R5+v4gZRNrANzA3LVBx8YlA1QKwpom/+EdQ4rm
JXy/TI8UdMPJAQKJAiZJBkUJ22+tY3UAV07c5qQRnnzIl1ODBknL5E6RuwxKWD4pp5PhhohKWPMF
JcEdHId6fHkkRimU5QdTPRtGHizSBCdmgoZaudLLJbiEH8G7p6fmtUEvUA4KTAr5cvacHUA4QH0K
gP37P/nhs9MUhGhtX0mXmjO5zrzEHB6sXgJO5AIP4wp0pFE5zlUqKM3MMuRl8FbaTUQ36VtGBfzk
0+QUrpcuay1rtlrIPLpAIFnavGF+OcZMj8SHcjkX9S6kQr4vGeiEWVH1Ke0Sn6c+Y0qugqRjd7pv
6mDvKrfEz1DcwC94r/dC526x0gXRZ0nBfcQ1zDeAA12gz0ZPDra+u0wjM6AEpTA0revUUSpvJByq
tFyo/iKsAE7gcN/9V/zcB5sBWFW6uiXB8T7m3tDXq+DV/8vP0MXGJrtf9lfCMAijbBvLZ352UUZp
ALHrs8oaUp7pbFrwBu5kGJtsoyIFEC5ZD0NG+hzeWwlKQ+FLalYnGH+oDLNhU7yV2CucWDyNCCIA
RPIZs+3HlUBZt5O8m3wePJx61Also89N3KI9F3w0VIaMTIFxw5NPb8pOJ2k43dfpP6SrTCx3TZoh
ugD6ZU+0ayt7qTCNv78G2T92mgcXjuGASIt5ZMZ3Ojn8pi/kJyfuB1V5x4hSel0qRpdw+0cpoZv2
aY6spEx02lQOyd5GwuhDGoj5cQgKcfQtK6Zo0ILjRwdnMY2j4pLZ5KHLOZY7JPKzpcikHb8MERvj
Awk5/V5VDzTyJZ9zJz309TJ4fu8YU08mkfETL/yJQzX3vUK6GPovsVGkt2ygiuWT28wkQFFQcVsy
mvw4fiE+Y6GrixwyHcfnaeb5U1gVeH2u/6Dph0oJrkKoL5zuizguoxQTd15pjfXShsrWQjW6GZR6
pd+A8GHkY8KrhGKeaPwF1ygX5fMFcnHq/5Zdq+EScfWedbQsPuINUy6VgipT2CncggMJVLI3DMUg
cEqIbqF2Wra5w/6ybTgXH3fVNYHR8EhGetvm7UXj2H8UQnBIsvUdtGrqA3eOzmDeOuIADYDS0wws
gO25WQA73koRToAGO5i3UefhZ0bUQdK3ZK6MNkLCL8WY+RwdBMB/O4C12JYPOdwLk3J+3b/bzzph
Onb9TLYM8js/tpLjDM/vUfNhrZMciTKsvbpbe+3KTdLlnvm1vd6ZP7VjEK/KPZlxTp784OM8d5xh
pJ3D41HJdFe0K01043rdoeFhEgie+Lv0ZI/79bXxGEMMCOIzH08+vDGNz0PBNIyWQ9fyhTyA8IrO
Z+wTMH4gmY8yQ5qXPfwkkxg4OLT8whtJJecVdNzyCQNRtJEQ8peVTtt+SHymiX+ARHJ08zLNkMPA
tPCk9u8uglHalng3r2r8nVBLwOTYDCyR8rq3X4oRzmhZT97JCZIFSWN5mKsSZefE8+eYB8/mujPs
SWN4YaKVh8fBTv7gC/Ll83noIig7u6zqlrqUjulCWMXKIUGIkhamRqifGdP2iFkvMzH77ShmWtsN
GbHZ7Gx24e22g9SQumzGe6X6F0daM7NUk1RZ/b3/1aRBVyy8BaHnL6jTENXR1VY5y2HQQ8nhz3wL
yjEcuCLRg7IM8QB2Tii2SdxSB6BrJjxvnlVORWSRW8m3nm4mranIxYN4jcNtpYT+y8kdEV+U0fiX
fcHk8E8I+ToN63fnSIrOXvoAdiaKTO6obOnMZpwZSmJCFqjZgalhSzMbt8vDK583BBRuOk/vOvNl
ijjiuBdsTv/69Z8Q6o9bN+ky7dUbbU5a/ldMrwmKMab3MlWL9YTl81jZvp1ock9w8T9Ef4flybZQ
YMiTP4DTcEkXjRyVopBfGMa8tOZkw61bpsnu+x8sGSDZ+1DRLymlBD8CWzDIBJ8aKzHQXR40EVMe
wyqKI9ulpMff9Zn3SLahcx+gzGRvUHhlIk3U4Mr0L/oam3fApAnl1dDoNO1IR2ERgsmRuIi1C7Av
FIJElEKgciEWDjSx9NZD+hTZotMUldvzoLuhJWZ6snC6FHUy7CEvH5bkDLtfUGhmKctBUpMV+G7+
MT01iWaStpX/d8K2OvxarJXUYdF032k3C9FuIR3DSRJAhQv2TZ5iGIZWw9rex67qdgLmjB+vJ9tr
OmEgi/n/ZFqHnl59dUhMk+PWf/nMY6j3AW2x9HoNVZBxZPkSDk1cgfor1Xt654TViljDgFSVvcSq
RxOpk5V7lbQlxYvGQ9f4hTrK5Ho1CcaoaBkzyd08eyYae+7s4vDXKq0Ut0dNi+EjfOnylSi6Uwow
GkNGinp1jHXKCYANWBizgF2FwvGS6Ed9XYkLBhdquvxh7J6wzPXTSzE8uN63Oz2HAbZyL7NzV4Ml
ifYeEVKwTyiBwbm+ZUrqZhbvDYiNfMIv8zrrjlbqw/XBMW/N8gyLOF1LS6BzJ1Evy4Syf/yZHFR1
wp+XlSleMFHMAR0Qxr8ua8kpP+ww0rZ7M3ZIWxG02nV/vQqtqDM9wkQyb13A8ZWL9BGf3LCBqOFQ
RbbgmUnGa5iFHLpEZbLIvg/FYbVrCRl4D6zhVhj7HwL2T5mhYH3guOY91CSy7pkNP70z/LR6WGZj
PlMNOM2sYJO6NamsyT6mbPieuld4FFZQiMXxuC3Qn2mciGJyH0Ju7AILTyp4F7HSe4q1rW1Q1Xb8
YmdsefRhxf+jG1YJdTfM0TGhd2To5O+e8AeRwlexP5+nIMGoC9kfvlV1kdYxWZ2Uort5ddjxOaFc
YB1/l87woFvFMPWqFL8HIT6DuVgpc7tzNYBZZBM3Y4xEToTPrGR8XBNCJien+g/pAvH/ltMAK4Kr
PUKpIk5Icz6O0DVadeY1Z6r/7e4yDVJZvjphbF71JOpBulGrzKG+6aFbrUQ1PqPyGpjvHRweKPTX
I/CWLEQVc1Zetl7bCjwjz16yWgK9SaYELzIEAjVLdqT5YUunEJq8Mmv6UvqWWZcRa1xeTospvZD3
WgKRxD7MAaEE8w0BFsVy+d4W6hfNchzvpjUtjsBPNogAEJHRxDkqT7T5kl9QRV4kD1a4uhdL7l2v
vq39HFnv34UoRyb750cZqzn8YY4nxWSBPjvCnTBNTlP82dbqZexFed3aPRtz+8avMYCQw9Zuq6C7
7A6II972XXJ1GvLFCDOViWcE3gade9Ml+zc00CQWeWnBECGEK7BcS9rX57kKFblOTCWXFrfHL4Fy
/dE5hIKq3nX1unObUneLSCkvaEYFYoyJmpH5YocmcdhuIRwuNdHkxUqY8ynUnhy9nSCdlgL5zcNZ
y2z3v6tMbJWXhsBNC8SyWfehmvLB2EM+kRqkJAz5l4/7u53cUIeeDM6mciOqYLSrZzYmdwbAwLTI
96nE1jrk9FrttMLndQahUO86mC1OwlnJENeHe5qP2mUC6E2ydY/NwStw5X7tNARijnYFCOAOw6U+
PAQEP/65SnCNHP9tzAMGxCJpeweBOABSZ9S5etSEu3ZJqz0F2WA3G9LCot6Zpkg2kZtBiQJVgeyv
dLH+g2nvN01I72j5ODhg8huYDO/d1A7cJ6Oyx96Wb5EhHs36f4KjcjifkDJGS2Rl7fmJHmDJqbF1
7qz2XHEA24ZT1UV+DcrzmXYGbSs4ZcecJ1TnEa9CUidw+Xn1zhBlSSKcpB7oeQz2NE+/c3kff0XY
KRnGmVUc9e4FpCTikEIbN8fHSxZmfbTAM3cQN2WUPIVlVT/vJXMsqabxRSO2dhAJNRmTXYQTQpuX
uCn2eE8wmmBbV7rhAI+hcGzlCYgxYfct70J7rg4ZS+hRROM4v2qCIvp4daYy0j+h0POMAnYmB6tJ
MHLDXsPWe8lnltQ4egBQP7tUbwqGfuDdO6VbbYqV6tCM3I0nyUujW3QDsIC7yw5i82FdTE+ZY1Xu
Iri0fHxT6WjnReRnKhECigWWow8SecWfPjxUvbRy6YQD/UqwVuaOUKeJkS5pfzYKnNCXwZC+LrOh
Vm1Gfr7ECw5QQmb83EwreImPJNrX0fIEGxnCHbeit5M42jYOMGDvyes3XuRG5FYqHPvVUXfN0k04
v0CSCgNHxki59f/fI66LFQlYzWyhIEzeeTHDuP3TV1EwbcqYBQ0tIEwjPFP5WCWivYzRSFIOBcVb
ezXkLiq21uN2vStumBe0h5PSWeFpkoC+h3Acao0195IJrbmOBUxpiRDNd3ABSZT5Oi+b9vT1VIt3
XaWCwXxXyK04gvAt5HjHPJttkHjKfSeuRLLzG4A/v9E9Xw0kZhdejCT5hA5wxv8BHJrAMJQSa8Dz
9txrhYz+9rJTPUq03jt3IVAY9aH6kTvWHWLEIuaKKu55FJdCuDy4oG7wPfeDaKxRgmu5gzsKvE/y
PrJXHvPndUH7eiG2s0vStFV70swRIHGpcC216ZyDzs2Q1pZUgf3jmlqnC8kQfefTtDP7xeueoG7/
I7Yngpi6dXEjGT2NwRJc96mVdO/ToQuRP7bC1dUrRa8NAnPm8LvPabQmjQ0q96jmSYVbJHhBoLWi
wbMIjWGcJz9XouwEJcOwNOUHHXZBH2qCcekawej2qCuhLcWxXSnr7dlbOwRy2FEl6YSm79B7Mk3y
LvLbfkNa1zl5Uid72lsY77G8STW3cv6MqUssXMnIB98Z3G7PR7+K84QCD5edDnwD685fTFo+3pRz
nFztiG5f1vYz59Mm3PWxVdaeFilJb9qkrKTiG9J0NL7C5lhiQioE8LYqAOhiBFEK1fnn9mCu9HU7
/xbl603Q0XkuJ+XOZJNYJ/omhs+ilryhhVCY7AqOHuCStwLPi5CvrybKxhFuV71t+Vp7kVefniuw
/v8sSKQ0/I98hUA5eRl0E3IBud7iKT7b6X/Bjbz5O1JhpuXKrbJxLMzYgZ4H4P/4NcwzH1Ak50q4
Icnd3tjbc9L5ZTyWHW2xn/nd9QhtXPV8nz3fkTYJp2iy7FQHyHCjAC5rVt7AM8b/CBf17e90LAWF
4D+Zd5eCRtp3XD3kmO9RLa0NA6GCaCii/mrAOXxlVy5Xkxl15jExDBvJIN7hdTAowkCEeJtjx82A
100Px6326UrMPH/M1WBvqvU0W7lIJIBKGrAG/GiFEPHRxrTuxR5HyIp4F+sWvNblVGLHdofu4DCk
fDFDHnj9zMX89K5y5HYaFLgSxF6Km6ZkKqF0oh8jdouLtrAfpEogQBQwuBiUUHh9mdIL5kP4rGAg
PaZNWN4trrWFt7eUF+xg5t9c+1SzdbawHXL1hJDps4s3Lnfv8hb1ACbtAvNirH8BGpeGPnSEnVJi
Zi3F1V3EK9it4gv+0IQIT/SHlDiS7m3HxxwncWEgKC+BdvN0prjdlHEubobLrt5GO/7NquyfN3qW
TWrOSScmWdd0t/nU+tmbZyJj62+8QL7rFgYhGQ5lUEgSqnUt//Z2OJbmwD5Ci8VkVG2g1bsC63lC
RFm06u2VGAVmYXtd/rJQoXU1fq2o3Ev5jWpJvdSpMjSGqtXtFcCObbYR11bA4/h3DZtDgC24JFRf
BSa+4gYs6wJhOo/J0YmOmajUXTSazcfr1/jCYc976LFeNyireebsxjlpIDI9UnfOcXWdktC04bBu
Nfv1ylB8DIDF4CIe2fMqzKG8Q98nYtlfS2SkipPQm2ZQ2DBc0nYqVw0ubNf/kgZxrCoO7tqiFbRc
gpGhDWecOeDoV/U9rIAT+9/pY733i+kgTmUZ+WY+BAV/ivud6c4gIIReaJM7yuPOTLZ/JuhLbMYO
0ctbM/yrHzvwe3z1bP8MOTJrUhesRAFZchLONIXWvxsoFOiA5VMVmZ7ZhfHyhgOm6VKF4BVTtsZP
16Vk5ikOWaoK3Qf06yrTGHr39KrBOoDmh9xrdsQdcdubbKWsf/qyofoJhBOkNHU5kj66FQXriGSp
jBb7fdyWNrJk5nnzv5z1ofoYt0HBxIZIc8Bpu9KsNyNL1vm6czQL/wkLKMTqCxX4etD00W2j+Mlm
gPGrNRnmTFqOJrKgIGHpXjDCd/7pofT3dwTPOn/t0GpWm4boWEL+GONxPCu3ubMPJH4fW/h/Vgn0
bUu+XHQ6ANLrVzLJs+xXAJfGloxBW/w1rii8YGz1tobJu1iNeq+CKuXhRlo3QQ2B41UDMinL19RZ
FCyXcyBRc0Hto/wvn9OE1uG18S9/raeRj96HFnR/tjxusfWgVSTsUsdUZxmksPnJnr19ZeR+hktc
9JJUCTz9cMw26eGgeZ3/bAGpnVum3qkOREMLdwl/6cOTkm+zpnLc7fs0yUtflBlIqwUTxvIKJTBs
ZMpmCQgILuuQxYG30Ogsnf7nsdfJdpu9at6nHtGoLEX2yOcOwEeQMb0dVLt4JIoI50wIvsrebLzJ
kXv5r4kTUHGFp1fM73SD1ztBPDFoz+JektA7vTuoaLxkU0hWKxd+mXoeLk/l1NaULGvTsRcY7Kzr
eJ+1Yya7bS4uUbUER8pWBgOhl66Bo7YdR+R54/VXE5ms3Kz7Yq9YUosVyGUy5IWVy8IxKb5dt17H
MPtQ6gNBKSSFo7m4NOPX+gHpGqdfq9E08u9veAxwL65Xwm1mfnzVvqP4V8vASh13gPI1osnqWxyu
TQuw5mbWSrHOWYlGMnXGwP6jlUFaub+PkIxJ0Bh4rEGfSlMFRHgReanH7OAWigW6L5cJUm8a2Mfc
iyEXWE/60FQBWPVy8CviQ95A9aumF/BB3y62KPYbkr4zyF3hL9F56Q+RCEWgP9F7irlz86jbtF/6
ym3fBKMcdYRMqtsS1BtOM081/j64AR2vAvocYVJsH9j+IH38tcyuL8Bxd9nIGTnwpoeOfc5fDB3E
Ab48V1Yfqj/7AiUz9a58xDawhdCXJo9FujRqHT5tHAKkCt1RdRNjDimXlingffPLEldU3Hvtab6T
hNS6Wmf2p6JAq8ySFG01p96sY0pnB/kEveGpMyvzlRNRWivSFKHHabWV0Mkio/3TEMcJFNHIR25W
4DCNHipizExgIxvL8mptQiR0p26Re/ZDStsnj3MDaBg2p8xHt286jZHiAE9KUtZgLBVy3Pa4LCwd
SvPBtNtL4vI6ySiKLzvCZ2KloYu16zG+dDf3bLAAiukhycyH0SEFNylVbL6fgu12yErHoF870xhm
TY4DLPaATaMJA3bRBrz+8aH58IX17Yt1Xq9HIBCewMkSM0TeRfbnecxdRVQB3mjpOjulwVoKsgux
OVc+cGSPFEX7Muh5C9SuceJaub3hVbMKHuBG6PDjnvT52XkJmjLEdDAOIl5hlxQ1EyGhH5Ypkj4p
EuGedKMlUHHhDXqylTXQkxm1CVFDOF7cQKRZNj5Cq781yXGoGpsaJCDcSzqUcpCxfi9JAl2J9/iJ
6erKlH4A3gD2U0BpMcZWyueHvY1HqvZdTGzZTWhNCRV/sJ8VIODAZMRpEryMaytFI5kBccSZ6NzZ
6pCusb6WrA+axM7PAg3cTns5DhSToMJbMVdFnN0qRENwHz1JWteN2fdYtaQA8/s1khfVmUxO9ryW
Lyp7cTGFL47UBI+Z746W1HYsw+PZTDjHMbckrMIGQSMryTUjO+VlX6xd7IXpqykGhMCPJippp2Cz
Y5HFgxGcZG+Hw1ybdiLxzcSkoWAauNbkxVJ5mhwTbM9DBF83ddQqzSmf2zcHR/VVUSm9I3YSdfS9
DeA2sq19ynB6QBIh+UG2ooynB7YN4R5Ttp/+etZa3dKLQJ7/kkIFZVfsor8m6w7sV/r/yQyd5arT
+0SHRr7oGbijAOSZb6mwSmHZhsr8PRMqlVQXc0fWJxR2f3j8krG3r7cUU8a57vnlLyLsY40Yl/P+
rPKlLi6qp56JUYmSBOA5xKdZGNgkgUCpsVL30Y0DDrn+0vuBklf1yyfSy0lyRHPP/DY3MsAWBC3l
xN2yepvwM6vMNgy+4r79oWSAHl8okzxt08S9lvzq04yIFN23NL5ZCUssvb1wKzggdvAuFeB/8XwX
ufSCHcuwpO8QGHFQAObguOpPofvLS94XzBjwyKkOj4hXhjWjtL74VD9DDPD4IVTcfigmOLcJHgQX
s+CfTvG+TqtPuyI+ygZ/O+ZePrzBSxFWXvSjhcAdVqhD8YlQ+W2WtCyrsSt5PZ+RVGPUSZkRnBPv
DLzEhTEEESnxWcZd7rbxV1UJW9UsU3Dr52rTZ2wfg0bbLmBhe2BBwz0/AdEYdca2wHKXBvyXE0D+
ZVpqduvkVGlveFNhgooTHiuGOWJAxNdlrIbGuwPugXlbMYlcgnu7GzIyt0kXM/O9whssjjFuXz0y
0rW3imrbOzJaP8ugt2KPh4jXsc6bUs1KYBMRtlAkBqTxpDp7uV8ZnQRLVu8Kw8zkvrj9RR6eJ+Ro
EzvH9wzpAbG54BfiW6nB2t76u+sm5N6swcfX+bxALtNWw7H04ofz9SiDnf+WBNcTLU+Tk1YTd/vy
fLf6b57mzQIEHk/kgYPIXjZfzvy/Quoh6ybKMkep0zoGzP/oHmNX3e5DB/255Hb4ErW8FHCbJjoM
yqTMPlo+x3ZxwobNTHeEswt51bImV7udH+1HLCv+mmkevVdMgWIc/zKX+WqLF4Ep8bL7zfwfAjBY
zeHaeXYWBBmfTJDLiXGS6qfwvtSkqyPmHXLfUnpYoNiAEPOmO6C7pOLFT8CHN82ornQkHCfTlPyp
C+NshD7WEb1pR7eFnKaHnAsdgDMc/LqayitE6+EAjJAi6+A3+GkJZDA9Oh7IyqkEj0bzLxcqS7LO
jm9MPHc4WHKcL77uxe1dnbg74r0zN02878lPfRxkrrJy2Q9lB33BoF0ac3YR8t+r3GN7Zrw/xz2s
cdh0jTvv86/s5+hFexIyeOHxDkTenjZOs/c+uZCwQLfVLAZhbrefQGVPbTxWt2mu6eZCcxVZP1bG
BiOfRStPs35H45TLdmOk4fnvLs9Mplv1A0pnBkp2sR/tjv0M/GWIgILoIrgebW0i1nBoha7dTp8m
0eTtjwR/7HE6VTnrvYGa4qMdP/SA+pvx7sjK/kWTNgNUs70nYN+la492kxk1n1uM7/NkRGG6y25m
ioEdTBgpTffX2Fhj15w8RbrIMSWfVhsjKvl3O/j86fpaFilYhnF82t/VVV6z7kdXevtVOnuDI1Cd
8faYSsXDkOA/S+KlscqkzNcILTn5ZIPl41nKtn+sa2bVkyd7JhKhLcbwxwfrocbeYm8OGt8fHgkA
wAeNFv7/b5GVZ5EQAuhg/uTCe6gjgIhujeA/M59FC/ib+FZaM9/+2HE5g6sj21+zqx+cGXer1OC0
cuSip6mzqcp8bFNZqiw63TDdxca23FW6i65deTYaePAjiMjQX6khya/KGXRyQnYjDW7TLzXaVexD
dVO/CAVi0uxIQbFAUEzKWnhXjQ1kkJG/b5FkvL36lnH0B2sU2dVpEJFv5CgcVujVHihwX7Z/jY+J
0kXH9dj0RFy3WDv6Jg7wCwIvnyjIiQ+6jBpGwoP/HOelLvZgj/qcDBmbn8Ky/RGS7M1DcnPsf1Cc
dUGFDFeul8+smKGiS/vMZueW4R0Ufh1hUIMyv6kR9tbESodoy8490M8ojSmyBPNhEq26yXDnz+pU
vpKiFyAsBTjXpRYaii25DjtV7yU1jQbqqEJ7R5qgnWNGSY40ObxGtnfLU7BAcPRoBtkWHOHS3Nlt
WDrMSuiU3Lsn3tWxn86LOEUhaB+YaeIgKrY/gDwAMiceZsuL9uW6yUKlbe5nlEC3Yq0nPmkIitIf
ignf0oW56vtAJGq1bZxYVTc2oKbhFTckqPqFMjNVpNFRoCt5npvrYqAOANlgkGVXHmIVCeJaUww9
fyaLZRAItQVAJm9D4OvwCnY0dMD0njCvkkx4BsrrTBarae5WdaOSCyhDyaYhIAJ9wTX7PxPRzsGO
yaUD9oQFLEMAWja8S7GmWXGKlKD1NUl7vhaktLfQtBW23isQrGfEDClon06WpqIMY/Qa7GqGypoU
xCbX2QFgwa9Hv7LB1mOAGo/amosvNM7mND3Pf7KdREUfE2wiaHHCLBMHMG9//OmkjCCXdmKJsZkj
3XI6+pQgJc1RSaL/LxoIXcF10MFUAag2Wq1MBO3Rdp9CD6xgiGfY1VE9OQQZQxgje5z8+DfbabAf
5mxBxubv0F8fE1tina1jwa16VpjGS0qNlMLMCMqiVksxKekbqt4d728y/RmtoY5KzEbw73T6uCn6
AUM2JR1WU1UovnSJaY7y4oj/MkHEhvzHRysa7Q+9FmlxL11a+6hXAUVrBi3QveNDf+fM1VVtsgoM
ykUXWC05D2dY1ANZ/e9sPtcPx74Hl9OwTqkPp0HakitosRXGUNyVR0U5C7PJbkAt012jOsU1F5t5
KtgIJ2y741cwlK4cByMJKLop0LXRU18Kg+9HcZJBl/+/c5HwdCVjsDNt1qIMJKBSyTIMkB+6mzE4
JT+wzYYX8aWPXkYs01E35kbtmPHQE8+obirwUp8B9J4wwqr4P8EU7fmPtLYF1mmqR0zuTVMqcOFS
tG4U3XdM81HYJ1L2I9xMMZ+u68UEwMWLfGDUsfvmNRUIoh0hkQMI6krRQLG8AKUbpjqljn+R53ew
w148EJ4qInV86fcuirdmXTcPAvbj1NQ3I0f5UQbzAj50Q2L1gD+6ODxhet9tQpgFc3i7UaXOT+/y
iBzIpe6k6I02+QDN5J49uapGclRJRRKxS0Sd3IkwPoEr7msPxWd0KyDqx211g2lNEkgwE6qAe8ww
mvGtpZi243yEU1zE0W7ODtoiZqZIwKgxlgxa2Fr/kjwr6lVxWybAFOZZg2fUIEoZnqJlZVuUtH6p
3kiTot0e1Se3clU5RJaSRm3TzdmP1cEAYeVZIebxHMpgznbK6jtQhkmztrLZ5paxUzxlJfVXXtT/
eFveDzhS9CEDV0044Rw09bcHWvnX/Gbbb5oBhab9qbAqTbbtBAbO3so84aabc+Du213Yuf2b5t83
0SW4VVRuVi4AltyHDPSEW1PaMQ45UvC8f94hmRpwlKlX6OUf4hDWj5smMXEaGVuiewChuVD5Y62c
mEqS6IL4SuyY//4QnKf7VQtHL6a2lEekMNL3hHFiHDQkvpHdA5pl7UoKMEoDpwr5PKtsGGW41qXM
2e1NZyEDUNAD4Pd3UZfcA3xXyxXSXkbopCT4V73OwYjkWvBSMaIbR3WjDy34gaQpkrtqtmAQr1R6
/WNb2vGIC7zExAPfNUDZOO7yF7G7fejSezFwtIhQsJCMHP7IPHWpRTbamIZFFf610f9P+gnX1owa
4EO6vtHDKGXzi8jXXZ4I9NXLXSsbTULzh7tqg1Z9N7pb2NdsfM5fpA+P4tP5U8X0t+cNI8QTfU0/
ZB6cs4WTDqJz8BOKN1N72XiTK3n7KRaej1M/yMhumKgWXC3a2FceNwBZvUJbD+8eiyA+KueFkPx7
o4g4SiRrG4sD8/rQJCBEvq8D3ps2Cb1Ey7lFV1g7szg9jrsR7W+A8jvOQQo1MNuZMSV0GSPnhvzZ
3GLZmOrYtM3pris0OdXH8VEgmsG2WOr41lDvK2SUa/eRNeoUO3DHA0SsOF7zOZsfRVY3t9Jr9aKO
IH6u0XIQxnjMyl4dJZSJJ8okHkO+7+IVobV4DHqYtIBUje7dMJeVVyllRcKxzFmIRXZ/HJjxGnms
NbOxRJo1TT3sbV23sGv7SmZE+kfbBXEzzmMfJIdblIzkmfmKoRdZPVYDh+YvsG3xK5jk9mfd4ayz
qIxMv/zQBNlmbhaRtaFscw0a21TBW2Ec6Hrl88ppMoJ+7btVl6IaDhP8HLFhcsrQ4CbTfQi+CxOi
CX/ngM67ipwviNwBDksQJnd+bUdbnzzAqmueszfyhrQ4WeK/gtXo71PoA1EZAlapvo5nXOtlUJFg
1G/hn+fXrx8U6zKkmLSX8TGrf49mNi78kvO4mXd23mb1a90Ay5N2KcBoT2prGtcBt3p25B5IkqpB
IBRUH8Gr5DNUFlGzBOf6xdhhgLQBrw9hfqQ4Q/81bq/e676pLJTNjZC6e4MyaltbMxaRn1SZZWLh
9thfbh0hO/vC4fa2vA4fJi9xVKvsyTsmm9OfM6fatmkBvttX3rhiHqMm4Rh0mXgfCMpIPYb96sLQ
xgOTfN0Ai36VNLFGJrZl42gMAjnghQkA7IznFn04zzPaITAkigU2IoWRQx3bC7OGlcrK29Qoifxm
zJcv5zZfFUYpvBr0hCAOwWSlnBZlm1+XkIhgtU8p+BDDgHNjn8ptlrEz3U6nMdNdU1eq0OFfPgrW
Jo4KxpMV2J8b1ba8K/GdYzPI/VXvi1wXsGwBuLV007oiPnEVeL4aP1xnJ7mVmQUmewByK4pVlCvF
XovVZXKXFbnNorNGvYGouuBUX9NAgPpQIIn4P16uoaoLd/cRFWIqb8XOwN2jJ5+3K9KGvncW+nWA
NhvYttWosoVMltClGDA6Xvil5kdgRoDD7TkzJo72C5ZTYeutd7xOvILg7qj/0SHKMJ08qzKdZUYs
35xp8K9MFrtEh7YHOXtnOBNSIzcfax7ysV6E0iIUV97xLtFO3IhcmhUv3g7oMRvpJMOL1rPRwgNm
6d9oF9IKYU5PcWF3Uz0rgrnzdeN+ZkQrrwVzx2Gij5WSQ05MEFH3XtIfBMtXlCOtd2FTze5TP/4k
xRq/3ZvTkycy0hVapomDO+HjsUt4WKm4BnDrIk4Dth09VEbNw2UC01fuaRhjMpFCDqVXx+uNAJz7
xagIJbI9PvrO4P+hqHVx3LZaLJD1zWdoSetTBJJ9prpYcDjDBUDj6zE90wRFpkI3XP13M6WEWteR
3lAO7desjQcEPNb08NELHyseLDH8jMnNeKQEzCuUJ7AQmQwqHJeMLgT8x0oYgrOvB4DTOB6vIopn
57d3/kD6mmhk7asSMpe96GyUiZ/z505wQ5gqqSbymREi0tqojOPV++i0IN/CbJVl6RLfB80Ldk3J
UI+Kdca+s+Xewin6XTO65y9LYvFXziFXWB0NUldbwp64myK0hJqeRpUaBiKlbENjA3VU51t+ocUa
Zh8W2QJ3+vo6rjnT452AuUCFIBFwGaLDQpLqdSJsFwDXJ35fA6rE4pYJ0jXwCphGT+A/MdRKE+d/
XnYzrKFqOBB3fmNRij23CLaU0EFIQGinYk5+QLp8dDagki8PFvd/c/ZTeIDFS4sS9Fqj1x/FAKhv
Sic9nmXvrK0mtVnvlIjkkY4t0Vv4vrJWROOx8J3MqXu+4T5fe8aHFPyYLdU2IzeMzf2U0onqWvkk
ROXqs8zkAzIy5QoXjOn7nENNXQA1Oki23CZ46k+M+X7Cz9kgkpjkT0Zv2xwaz+NJH21gEpw30XM0
8mjZDiEcUkYUV+omUC5UEHAtxIGK9qo1eY5YtYw4BJARMChomsOD2mL4wg7RqBMSu28UO9/+/ccV
ekbEURSFk99U+XhEOacuUXVLASJwHawPdy+YM83kN9CtNz4LHnCNyFavW4ygWSdxORoBEMfdV5n/
nENuSbsU9PpAzgWiPwk+ZIh0NE25uWvo1WReyhxLdg5WZJBiDBU0p8Wnn8xHNbxaixo7YjVGLuAV
hXEwN6Xx1OV1sIIXoZRpGvT7RTj2A5kvfcAFFDd5G+VXy+feLHb8PO0jO8gVTbsjnAKHzo3IkJDg
2voEWTPZDCg+F0jBbbx4h8GqGVF3heBEo2LATJ+vJ7odh4B6aIOtI3gV/PX30z7sNT59DhljnQsZ
7k0Q634VEA6SjQ6T1PIqzpO1Owm/P9lr93YiACQjCjVHMeSDT06FxHMGF+AnlxltyIoWooW4KSfF
Gp5bzdo4GV91ysrmbYVuRGub86+Ym0IdvL2fIm8V74CrNytyRUx7faGu/8tjo7j8zNF69JDMjYCM
0zPu8ecOwSAB2+QZ4ZcxWgZ+l9beXff7rmjDvk4RSrcdT2e9KF1HXZgmmYBN5Ps1k+61Gs6Bs8e9
Rv6nhE4pe6npKfcCVlp59U1fBZEnlYTH3OTPetQNLR7/+sW576jkd83DPQ5HwyU/dVehXlvDo/BQ
uKvmwRSNY3/2lvh1oOa8UY+0murm+d2Hb8wFXn9H5200Laz+XyutUJkEI/x8bHEtGPrltQmpeW7U
t88Ng9y5VD3mFM/Xmu9dRX8DVKEWjXOo9QmuzbvnLsmRb2TvZG1s61dbv7UFgvGTB1B9v67EmliS
o0mlsvBom74Cn3iDKbjhtHLA0E2DJfjTnDvGOXJKduv1pTwLcbhyMoKiEq+A5FJa28HQahpV4kWu
k6NgBp3XJEWbbZviC6THz/m3CQJdZX2N6+46NqszJrgBOLSWK2MEwM3ZkIRRLJJe09Atazp9b+/z
yRyMgD+jEjtgMXuIt/JXXuD0DC2lJnPj/h9imX/Vq1NvXYdU/hjL16zOBQMRUrNokcE2hhld0B4t
AWKXCBsGeNMz+Vaa6Pp3fkHkamp0GIF8IF5Wmas8aPi0WbFhi9T3flZrXUuXgzTfJ+D5nqcp5JO/
b9e9BGc4VoRWFqxgTf9nG8H5BT/7/0XRzuX1S1yw9GDnjK0KbjHJ9dr8hls6pcS7ljjb9YBSvm9c
35s84XnqvFGDEAJ+UfqH4heY3NuFI6sCgWOUo0/VN+i9Io0HxHB/ChrRg3QvBxLUCQkIIPrdrsKF
k4zf4CvwCiGXyvpzFC/nXBSCyQGyr01YHwrXizdtYtS5kQED1vO+3Tgg11E4xdI8GcIcyIsHfzxS
sgOW8BBeQC/o8eJoyw9oSB9Nv67FGeTB4J/OdlU9kCAhcNeKK9sqYP4Tn8tIF9wPa3MwdPiyfgTI
co3bSPbraTvXAxCH00KLcpMH3CAVXn5j0cewNMmu4B+rUNECKx6A+X2RqhxczxCPQ1gHK/rG9KYE
czUFaxuGnhjDP6TWU7sprNvxTw9ZS+VfG8OLwyhv6FaAYpGpEfsbwX9tyXrBOJx1jp88rIzOFtLu
14H6elYLHiWhMHfST89mCfn+CkoVko1P66A6EWjrA9gYplozROljzf9eLjjHFzcWk5uQvd3DUcM7
wY9EJT766iB+R77jV0nIYMXrca6Chi45ZFFSkHsbA/ZLclpEa2wNu4oIApkIKSuGqZtJg40fZNbd
/d1Bz7iwIT1BWrnI7Gd+K9Q2e5NHl3n0mIKnq4XHA0m73A/SBG9sX8r3gBhkzH2If0zxkmdnZLQL
U+0YlB/LIx/Qd9BeDPL6m6cUjClG9S7VNALtqsuRjmu5/I4tjNYq6CjgpjNgxTrhVdV3UN2S/wPr
dcuJf+pYTkt5pJTRwDn4KaosI7p9MExDLkmPK7AWR99SdIMQO8pC8zcvI0KT5hQ6nkY0/A5lGsWS
Co3i3ETKenJvyl9ZVO8tqZ6QjJQnNUtHD6h7PvQ6Hn/QWv9jw4YBdp8ockOtBI39jj50xVQLvwAm
qvsr2sUvSjLqf1o4kVlakAamzq9lLdLLdka5SySgjWCsJrPJ1n65VQ6yLYEY6oJ5SwCFu2Gu/Q40
Rl5BzFB2rvA7QotZH1IexTYQksRqMzk8Jj1h/xveABw7YKw5tVpdIDrSLFs6FU8p7te1aoVqDi0A
iSo12iNEbYxTpkKgTBjGsN82KQsR34sPKKDp9ncKKDQh2vZjczRCYDY7loik0m4heq+tGqih50xs
mc44JMaU6fQ74R+jeVDxUdTw0aIzb5pCctWNss79PjIWgJGzzS/lgt7UfOSxArzppJm3pwdkWFrb
Jt7TpGqvXPSByjRRwof9GAl45PoJwa3X75GZuYp4QB7S4sc8B2c1M74WQio7pnlp+zBjg6jU4f0c
xAbE/MtadSjICumXNCbb/7pbPjkOhCRiPxjBsl+nlTDWL3FDQmf7hPU6lNdOi3B3u+9cKaTGMhPi
sFpDdrkIOQFLr//s9PWyilb2gVK6U6yc5viOCRf3LHNfO9RmETNIU6eMDFeJZm+y2KEPY4iKPU2Y
O3TUT7KRDGjBu4UMJVEbmChbmM8lqRAXH9FnJyXoGf/AJO81rHeV6BkyLXF7jPNo+VTtkQLnrFUC
SLQNPFHza76FPBgaapUOECdvKUNqBpui4A2RjOUa8Me5cFXOu8wKQZQkE8PEA/cWVSfTztV0Ben+
QT7cq4hO8rHk9pL6oEgPpvLVXH7Pm36MlxHeI4CaYftbSxGLcJSrWbu526nnvrEpNnKgP13GIsSQ
sgCKErCbpPb6WtzEi2cH59D7eGQdfm7OzAR0ts5aVNTceW2IN7oRXROQ0Bei7vsOToasfj4srbGu
h8xpwMoZ3RXTREfZZyzIhmbIP6MTBm1ro+2Y2kMcjlKl9srXSNi2gRqbomgQbktptneuJ5Txgy5y
gb3dI1eaxLTY+t1xlNfJ4hV8hBjIEN73vdEP8nDlbEnPms7eEKFFzd8F2Tb7LkWcshMz+AVzEJ+x
jYCvDbjcEMBzMiKB4RzCaoT4YRVU/KWYzsd9ukqH0wZ9VQM4vZA/vX9xXs5O+j+pIUrcUSjMjpjB
LTa07ZnVPE1FgBDD0Lw93S+Ss8p90ThnTgYxWFAumIji1i12X5b3YWwKo2Gw/MAK7BNzbAUvchIp
Z/MIY2u6/mqONdFHOI/gLS6uDUDAhlS1ng+tz+Qn/Bm+WB0anPMUBQnO9UIf9JCxkCvVZekhGSwK
w4eBpzbC53yULMNw0c+MgMCNJBCVMvlywyombRPgrUV4f5R3XerizUNYVlc1dBiHPOwpVcJgj6EZ
CfKeh2exEpANWqxRFgs0aXieVlHKRDFBdlXwePjRXPP83F5BnAY5JNzMQ9b6bkdcFqeEQ60lfre2
hEYEp+jGSayH7Fh7DHym7fgJ+HBmtPkZr+Xc1Gfl3LWc7RMgEGsOzK05MBIOPuvnctqKRQmyFbKO
Qr+jmChYiUf1Jtvzx35LeN/DLWKYEfioWfCfeMZL9guhdH0S446qin3SMIne5vRKzHLQsJI6fvEB
JVXzXzUtbas3hqexbkPkilFBRog+pLymdtz5MtgA9L3/pCDL/u1XKXsRHgygBTUC7uZHlV6AfaEx
oWFfNBy1mqQlUp/sl/vToXKVJrT6Lu3TQJ2DSAj89INb2Vp+GFbhvzKrexIpMSeaCdd7JMKHaYAn
9LKoT00Ye1fHhAMSO95d7iWOXqIQtdZ9+ow1vOfCWFGYyj3151klkqM9H7aI7S9WgJ34vlsJhHkI
hy/0LI3WhqEAHnuOI/TrLZlxIDfYWnSRJz5cTteE2+6346ubsJojAHGb6QjjfXlgsixkAmATJCMG
cyQzcDi3aPO92vVxEEotSRJuPtIGKq49eX1AabEodCCgW/skyx7OaenCskZ2bRimKhADY9jX9sjE
HYHF75mFi96JmPHUCnQrP1EduLaaoNysN1eiCju6rLZCz7fcnpO3k0SjX6FJ8m6mfjICHJiECWl+
Y21qLT6EwvONJdmJEmGyCXFMrhV/sQBlqME8ngTVGemvDcPPWwkfkOrHTjibdOfMqRnNV/LQFM0O
KfnS5E/6PTyb2PeXWRi0qPrDpoN7s7RenVM88CQKWmin+rl+SX9AXoBrF9xb5lGb6ivSf4L2R+NA
dTMkKuJSLunYDw+qZ2mUDL2Ie2dzpn5Pk/eWS+bZIaoR+v9e2gPVT/yOzZO/tYudQSMbESNJXQsH
6qJCuRRkzvM5UreY0JXHrW7S3onJYvFkHbK1fRb3hYBwK8219x4W1KQ8BkXmSaVcOSbNZgT92uhg
dkukWlku518agQzC/1/rNA4VZCLb3jiCQYgjvToEv67sTBLAK5l32jV8d41yH1M5XUjHPCi2XesZ
cE2yBPPlVeH0wpLofR8wWX4tSOVFIeDMHAwrjvHOfD6J4MIHaudZJ8CazPiUD9pl97By+AM8JRrA
y8r3nmVZpIMuX2ftTnuK1fRGGBskmRCzngvhrUW9USxtH/JOekVIF3r8XMZC+Z//4MGRVg1+W2JY
WksMkA7CNf31qX/FzNsIYP1oDfuimcqVsaxzmsSY5SYrHmMNEDNmOpTD1aGvFDC755bHmPCWi4cR
JJLzi6kW/PMMUpxwymwP3BZVA1s+E4gCLyb+iSVdCHV5gdJm6k5zOW/WWfbR1HbIY4Iw5+Fwiluk
mWO7YDMdTNYwh4NfAMWawm4ND8+pXlV3Sbjx4o20Rm6xUdQDRHB7BjfY7fPv0zmMPxjUGGqQg/lW
W0FgNVwMN0FD4yi8+0kFUC6jHz86OsFEiN+U9mVXHizjd6yXR0vmA8DS/yVS5H1Pr53ocxR+oaFq
dbWj9q4LCFyHc5UNux2Ot0q7AG24sw+gpCf/soRP77Gea3Pd4uvxvG/AhNIQ1uc2LH8wzGIOGH38
FCFbWs4g3wnubot/XM/BbAT/vmkGYkVL2sqKaxJ8gMyl7eBR2SeNNXq6rP/j0GrMah+dKR672qhi
xmlUUsmqutsnrXWJg8i/26KL213b4hwC2KlE2JaNx9ney9Bku+tQMo/Kn2+MT98lPWQNPOYEgibK
Q83Y3SDqrXJu9x0L6RP3GyW5MXlITZ+vRpEzGfDv04o91cq5Oa9vsWWzhIs2lHzkkbqWW27FESmy
6l2GvVoBUuVqC5WcLz0taso0KHrZLYZZ3dhQQAI/9+lKODKqmxUYjrmXHSs53bYxSPXiHoKqN/vj
K4qoWMClY0zK6oOFaTth0wbgMB9oWo1FO0Mz9KPU5Bgbqmpjo+5CQXy24bUUm5yR5biBOXf/vR1H
3Kqym2XQotr1jGaKCdZ7478MOuE2Ia+Z4Z+A/9okx074gQWkWRrPTyC+Ra83+fx1U4VOZY5dniTB
qIM2JEN+qCGB3RvNieQyWSmuWjoBEgXeUa4aXUY/5yZ9DeEIWWkBFKaadwrODkwH4o5yR0lC7+9v
b+9gGxW/NxXSx3D1x+ESXeLu/VOOy2/hy93BHSyewupX9eFasTkS6eMUBQkF0OzgPpwji2gjO9I+
l3PnTn3XuUnXj3okqRAeJm43X1xLE8iEndmh0be21+vyK7zM/f+ThWuAkMqfcEqNB1rFcPX/iF9j
KOz4+BGELZSbtp5Jp1mkEPfhVnzVd3lvV4xz1Dc7sZglxyyhP2olGTbpni3WNGTVzDmF9VvAq9FD
UrTm0Tby4iX9z3soUttfEKf7N+go3S7NUigQ+5iw8x1xHEBFIPOzGOlMdHm8/Bf2KntZSwGbJAJ3
Q+J8G5N9fjGOPvRu1HYknZ/YNu8PlmpIJbcyGKAKzUq2TFIQJlU/9efeYOfk/NB8/8+TUTCKVEJH
pXe0eXGCjkl4BmIigbM/Cz66iUVvKao+Gj4Rk5CePqA20KgriGpOxr6hX0bIYMP3knjruNoL4TGD
VLWDaTR0K+h56/A+51LOu4dr5el5JL82yWPSaIUjfmDa8u9roWGF2EM3yQWjA1rZ/XwlnK8iJii2
4Tp1JwIkb9eGR8ectU6wgusJr35lVTYK9bjG1duLbmV1W/BtIFskNf/m+SJ56tpPd/aRKOgglXpX
ZSKdSEO9ZsTxY8XrWZMh8LEnL7nBvrEN7oWgp9qDmmRCj0AhidVOvyDAiotETtc4WSPsSHP9VNUE
cm+hcQ7hNJs2/I2RIRL7QMZQz0cNg9GH96FJW1wL/wt1o9YhNOyZ974+2bnQsV17I6kszZowt31C
/9NZlFm/ITPjO4FeW2Zas59uEjTYhUb//KwVoGVi5JHqDfrkncExo1M9WR8rHxMHdKVM7w6Dj8Oi
ykvOZ2qZXNmJH6yLa2mXxSwEFKJBW3Fr0AxI6i3tlXKFJ+ClAOEWe3gBehTn5ORvSEdqyan99h/B
+9SdvUtSxRsdYECkvv4zJHsw9hZh0NEN8LxDeWr6xgS8iKZeYltXKw5EuWLixP4LLVSRWnJ/OGxc
l67EQZp488799xSPoc8yToSvkUG4VhrpMEPkY5IKbgd+Xzh9cRIIgM6febOHgYuGCbCYrPrWc4nd
1xkXTpvL0pelcFexp+ZAK4BeS0lV6FMR1n2Nh6f2qeaJpt0DflxB7QjCmLc05pQ2izNOiPY9Jckp
Z+L2zzx6478oulWmLJJTx/S+xyDJ5bOwJF3gYFJKx7zB9FrS7KUygUn3D+KshYrDRrdmHirIuf2v
r4NzAr23y2m69pGqxQm5scCN0U/a0Auwf/77NYBuxLEwdqmDJ1nnCQQsKNFTAdMnB5N6F02CHbJX
hePCwYgahci4z5yZtEQ3RM3RWxvB+KI84v/E+s33aC7Fb6l4np8Rs8KpQyudrrbGznEwrcFxZrm+
hXQlrH0KgCz7IBdu8ME9VH4NV+q56Anbi0HN2qrAyO9lXrqwBEK6o0Jw78Gxw3Ud3zA+Mtmx+cIq
E9RFzfexQFZsc1Jb8Pr1G7Qi6BN0VS71/e8uwVM9tPE6nUYJSJcJ4hVRZOnvnNb3h7/Cj1MwhMFD
0l7bXjtMKi1U/KbElzJ49XxLmYyFvQ00FxY4U+eC7OChY0FODo2dgjb8g4k3JmhVjql/mAavV77K
fjVHwAxOn0tsUbGVroDlo4DC8IUh2GYE6zKCVtrNNKTXqFQuT7c+ElS2tLX7TGv8O1ede0dX78c1
dk8bF5R0GcXL0gYv0EN9fpL0sb6d9a5QeVPpejvsN+QVr6K2F+X7wCzXT8tGAKKXxJT9MxitZhng
3jZcufN+L/E5G1REM4Vf4iW5gPHoofKHJx9KTX/DfSd5XAZg45gGENnhQ31WTBViD9p4TLb19iYn
TwdmlDydiZeeBA7lMYA5KGxsETQ+IxlMw2z7yo8uvyhEcZKz5s/7THp+Yylvbb+dMD/QK1Rzx99u
my2cGZK+ME7CIFlD59Qmsc1XHZSsAQESiBQSOt4Y+XUJunCaw3bsDh94t0eK+9Z1a0eajSYt1iXX
w0IQOIMKT/tIKtGEsnYOFmwiUYcWOQwcy40b1b98M6WW1eKsUDvR/MurEpk3NF9gXWDj/XXl4yeg
xdzhaE+qIJbP6xi3YdLlHGSPD9H+VKSlRo7XaMocmmk1uerxNbhNr/OSasDteqtuscuhld41//vy
S7pqQmvFVUX/qxjFSI+9IfNksQDmaM+4rpWIm+4BocQI6SV/4wE0nLX2s5+SfGcBvp4F9cyZywbo
avAW4ADfjJ428ufZYJ90XhqNA0Y3y3uO21otNn4mzFiPxCy1bAOLEnUOKM8a0upUpsfKYqSo5dcE
jGsQH8lOdafPjITcc80wSIHIlE9Pm/xYKsKR5HVTiL5dR6/EzCYrTPn3v0SDdG5axCGHxvZsr6fO
p6Ap6uZsCSxfmIM1bIo1bBsjxkNTNMiwF1TlqO/g53kxibii3mz5VmqgTBgsNgj4fLcEf0OiVsMX
RfJP2iggNMi4gYdtRtGCMKwBLJXGbyMWwKz22awwucV7F1EAcgTTZt47iX+QGs3PLO1ci8PYpJLe
jTZFb7VnF2CEKIN7vXh7XQdumg58MMvc+DkA0caJ1X6Nk1gTvvTQX3ewj0sAfEns9cMg/9GKVoXw
lDiMCK6Ypn8XD3NGWNZZz2AIAMDbvKHS0OoiC5HbKMzNfESgA8/vWbHt+YbHqFNyPazh1CRfpiBZ
tpEsRCpts7ZbW2zDH3xJKXtkfMEy9YRSD66K5iK5Fms7gOr9753R/cSjWp9NzryFpCWt85wQtguu
hLmNxq4hTd9+K8jsAElFociX3PYsJw0QH0o6VpHyLDcSYvd9XUKytdddL8KuRjIBvZFRF4VeRJGw
sn3SBerrpDPm/8F1ZFDV3dQIc9uaIS56ABuZkTPjeBkWIwiVAmBAU1Rt0AN21W1TVeIEkEL22SPx
yJYGDPlMpJY5U40gfBcIQDgoJcWAf4RB/jykGNpF6Nu44p9Z04ujPksW4N7KhOLSf98GUD+nx0Gn
9BwVR5BVyToEz399xy+k+0TUrMKXZfai3WgTKVsRx/8VTmUdrikJTOiN4ULTTNMwQRFnih0lOWAi
ZXrTA/5ObpvUR9JL4KbwfFCM1W92DJSXIIysB8P+qUf85SrtxUxpmXQC4fPweAQ5GyPuJObtnutT
+DfCHGwl7l4VWMxwDWol+V5OM8bj2eXYeUHg1X1E3TmyVMO0tRtMInqUzkqgzQC5qedPHuersN34
D9GZZzwz5Dm7XvNfyV24jqS1XLRMW5IePW5djxqZ99v3zV8T9u6YYNvNKtZARCwXc1IyHWHAaXPi
RZkMBjRUmKyjfElh8bTWbOkQbbkcmsyq7KUJDeadN17UeSMQ3NEBfSnBkcg4JKJ0HRhUK1ITT63b
oSwV2Oo89Ot0xc9airsI2QIJxXPqunMKJnMMTx70NgwQW4C7d5DPXyYRQOQfeqLXlyLHjKHQl4oV
x9dLJD2vskPs1KA4TBqx61TVy4rl96/Uqsm06DJd/9Mh6L/ZWw8i/ugehMzFcI4yqo8idJL6/3Od
FpCnddOKy3+0diTvuEuSrT4+i2SFL8ki+sevg19u9ElZYaqCMfCBakKUsY3V1bi3iZgW1bb5JcRv
rG/jO+gk4T9ry87QeAh7p65nxm5PUtXdkttBhUF/W3w8GT7yqi4LdT7tD4zOjpAr32c3rU7HUxzA
7IaPpHYjmxCiAi6Ik+YSERyNQyUrND0abeygXNnfGBjSA+fwGOjE1y93O7p+ogkKYbyZ7xTIiHPK
bNV6eoXmapqupPtx9uLbBQ9KPYsBbPXZOV7BEtOJXXTIrwKacVoJMsxv2VD83fj3IrYUL2mgFPOp
u9ZTmhp0SddEN1E58787EA3ctdpxKFXdXuuu1HBSAqH2FGAnHv1wFf9bx5okCSvibH6MSpggNxL2
TpbBS45mvMcpyYp2Qqs52w29XL8ojgH0BaxGQosMYggvmKuCew4YaO6vo37EW0NC55Ibd+wnwt79
NLJkY61AbsdEUb7JFkmC0P7FI7RSei1+wQCjG/0cjkMEP/icCaL9FDX+QWT1pTfilOjVDsjc7Mix
/0NXdihQwNATCspvwr/Q00Y0cH9l3IphSze1KmkKCnKyYOmcA2wdvNJd9UUEji02EO/yuhL+SFNa
DEmt8U8w2s5Um1Li0pdFANmXXgd8r5BLHdQCmi5RHdFH6OeQuMPX8R4KbOYnNUy4pzjvwzcbSrgz
IztXYFpBwJH2gAusrPfsctfvMYb3sxDKabKdsFoZWJ/YfGTphnHy+Zb9Cjx+oehKg7BJZJ/t7sWL
0vfAogMsnuFS0bLzc+4Iv9t4FfRJguL+91/5ozrFosiTwij2zV71P8KI2AegafPLTuYv6wj8qqhN
hZEzQOuw7+WL2+iMlo/3WAFqlOtUjRPkaUDM1c7HGTm3lOdi+Yem/3jPpv/DsUst1L487s52CquV
h90Wa5uXQa5wJ/kTORsSi597M8ciyCLTQzq2hhamv11sEi2EBdlNHvsGwAcjDYbj22BArlOsg/UV
b3RzU57Nq5t+ptGztQ2NdquvowNtis6cGntzRTYvAHAzLJw2yAIPZjO0NSauDcUGviy8HjRhhNXt
hnbAujRG9kSHQr3T3IZ/opobtEFX2TAwT4YxT4q4Nt73itlcxpWCLPz3SJAXXNY54cE320EOZNq5
vxgT1m5hr4BcTCyv/qfcD5zpVXNM1zuSNiBa4alFUNOLkqw9uoofPrwgS1NSnahq46uyhV8pDJjQ
/kPh163id3CYlEjO2Tadgkn2ziBZUAnibinjyk7IBjwjceIM0yUVB3qGeBeDjNFmBK4bHY5AQrVz
ue4spiUEJ5KFTeRq7FHFU1I2OeKLORUu+dlqJ4aqE/6JV9n+4swBwcC7yTtXnu/wQKJl3sYRixuD
GK6SK/6Wr5diRUiLD2iL2UJkeRDiRNFzB1PXBHno8QhvWOVRQx69f3yhYUjq8fwN4++FrQ2lM7xH
WXZ1LRtq/zbi+QOvmGc5SNg/WBqc4ljjmgFaV/DU3TDJYG9fq8LnBA0UTtl59WE+jVi9OR+xKTUA
7iIgCHQ8Z9gkJ/t2XHAMp+4Rh5UoD1p5WcystBFaNO/DM/qkOP56qvBJpak+Ixrusl+bWgoaCcmp
/hlQss2SaZTRBus8yVbQOJrb0UFm0YLq4auHtzlGb90PdXtmf1T0BnAKyrFzyncAM8j+pMoMgDFC
COUUAQawYa82gxsPlafSRJjBA6P+ACEzo64eczelRbVNzHn4HQWJ9TJQEo0k5hfV16i0Q+pSc+YN
aD5gFid4+pKXVRinOW4mHhMvGF5RpqGdXBbl+su9fB5F+ZGM2J5aZVGExiMkSMXyE4M1Rq5lrbSF
8F8O5LGA6AgFU/e1uxzQQqz8MFh2IdF2P8D3AEvk+TcW5Wmrw/eLSVethmpcZxCeYFlH9VPZ7jQP
t4zuS3d2CIvXepCNrHATvleHHNOzr8NMO5Ns0AGWE75e/Wmqc6x/uDtK436IekRxVf/pIDuJdeJQ
OMZoUnSVG2k5skkch5wlQ4s4otOUUV78wmk9A/VVTm2lRAB6GBMvHREA2hxHR2eVouXKtkEPaOST
5GWPM3Hp7nLG4LZyF5yBn1CUl6vaRbLk+JfE/+lHm2odXkTsBg7RAPkN5duf3UEpBtxOLlKX1MRH
BFR7jM2oagMgHVlrTZFPb+MreGaNZiqzOFidFA6lpoHjViHPPcRDNO0ACnj5SI/ZpT5Ldxng0wt0
oSgKG3tV4bW6v6OMkctKkz023Oyw/QTc/xwLmQiJMk+8kQe+KEuMVew2wgBRJ7S71KWgE8QxJR0V
urzl/BHRdGeRdXER6azigFYYusBtDiXHZ5htuV322+uIJr/+2pHDHvkBDgjWKGRv0d8JyDaKLdgq
+iGMsX5KVrd/dMruX1epPGy75kl+HoATI4xOJP1zuDrbQRPKivKUYrkliWgRS/7s2itYIbhXIyQ7
QcLwMNBOHal4/xsOr4S3i+AFQxzLz+Chi6gwJItHmt7CM9xVFSDXZVFZPyww/uZGBonTpkUU0Dd7
62ukeyyixeU9rr/TAdKKj2q1/ZZzUVZwzBqrcqRsovE4fc1wNoq2o5FVHsXbhLByBGzEoX6s7a3p
rdpFwrTa65XqTvZ8zLP33dHBFpNqc04NA1k/rGCWe/ZVaZ6UXSH7UpUiqgfy9ElghOXS/MOonaqp
sfM0oVH4oSqpJDe42xmk3BU8ut1uE4po8uBxrZkeWUk0BXmxIFs62xsPYR7/Ab/CwZBQKd84fEIs
bCRmpirFyntwGI1iOPAfRlB9PsWCF3x38TYAqQ+Tz0RMtynGBV7jlGsZNZHcsedLcju04u31r8ev
LPwH8vNV2ypcPstQelPua0lcbpAriY3qNAI4UQqiq4nEC4Gp4edeDO1wXrbowO37nWI2rBqs0YXb
vg2G6C0rsgtmgIqwff7nI4OBfVczjEcVg/9NuipzWdRaFF/fMA5q1K3NBx3boubkj8Nslasbect1
GerBDITYgD0c6Pbc6705+DjQGnWFUcIz+n9oquZqAwy/TyrG10gnt1VdEBXGKL4CkCI3kc1nDilK
/XD34xpn8sdppIKXkguXHjfoucmrBUMYwk0xyI+s7Far4GIfQO6IGJfTmjMyLQlsAz3GRoTvxRwz
41AqfjeviIT4TJcLFLrgF9bnP1fZ75R6eJL8yfr1Aq5GfptCgzjLrgZvqU3Q/oMeQ7/wkTklAK0C
WCjVhHJql+LiWPeLbbUKB2KbqZRl7gftk+SXtp3rrTkv/Uhc3TIEkspac3t4vLe7D7DAyJzqHToe
8eBLCUGZTb8wyppj/jNx3XRxEM8vgFjH82njV5xadXhU1fMy3TDpc/H7rAAVX89EKxGa90KtJryC
PYRIJHX9zzriOkpWk3mSC5TnbnX7PfUj+sti7p/wSI9s0OpbXHAnD1X9/gQJm6TPTEaM83nlckLX
D369HaR08O1q4wIJus4zmW0REsTxmYvPm8MhxSHrwroRg+Sl6LBGEIZZGznJF63VlzM3xsYwRRlE
egIJFnuOwSEr7GfaH++4N+Jb2Y680A/EZkkfRieQ4hAkLMYuHY7qaljPb+ZiXtAxgQypke7IzMie
8nz98vdwMzBHvs2tFlZJhooPpJkrhIRfk8wrB3LM1KpmbnE7QJdybgx+x6bzKMK5n3j6ItV1z1pz
GmnLPrTb8F78J+RuXyavDai/NOWoi0xikRFqxwPMHGS/b+KBOwRmXrGtv0h+dfQ3ev4+z5HygjQ2
JeQh6f/4T6S5sWY8vRmcvMywwO2VOURt8J9kYQ7mwfYhdwdaWSY9ArzwpCOip/2HeSM8OfxNciJ3
1lryh5XeZSgQ+l8v4sEY1pAnQy9uPveZvhVx6Hno2MrrEkxIo6VdvtYDJ02WBrP6JPdcnzeG6LHo
/HqSezBO0CwDq+RbtpUR9kwQ6bYA365T66fd63hhTw+7RQNCoDfM4OLuqGatzN2Ud5gdx3Zz5PRi
RzEwV04m22NdWHH3etm8TKFVJsWGoW3wYkS+YGRAxiv18WT7UX5zbphndPn1hJsqqBDNideVrH9W
2BYNrDI9t6ZK7ikL6je/NP5Y87r+vMOOcc0a2t2OOd4c9oWv7szjMbtG/9cQgH6UXhYyyPKaSm/u
V7XmdhmO1fJN7Snxp69EdfXKegvwfyCNCe7AkT8cltw7t7awD5WI2lyB+jbu6/hJGyd5VYsahT03
2TEMGXdOd+HOcl5foJXLt2Z/sBiT499ZK5k6Tq947bPVEr7WWfoKCZuZLwlZVYmr8PkrwNnuCTFl
Y5KARELWwnc9/nJSAkKZcnHOy5JsTHOYeKUA/4xJMMOU08AtTlTtNwURhmRtLjubDlcS4OlxXqK+
BBBRsN3nXtiIp8u3JpsOLnCzlsXu9usGoLdXVmOuk3RlM4SPJj/ZaK3kYk4wnIkTMDvz2+BYK3CG
0ZjDa4pBNxhhzI8TJXkw+ylEkRoFE0IkZIbRggb7MhC1UMuifQQAJI1enRn7/JCEqG3Jhm0XlgSI
pbf0CouK4rOzfF1YYLd8SNtzzvyBaiMGvnHBRut+iOJh+rGjTGzm7nOiU3sIzgMWs+x+ZexHLUsa
wUXyGDhluFh56sl82LKoknETV+5Fqv8EF36aBViZPYaNwNMnclFf6eX5p3mUJW9VIas0c6nlqBR0
T1p2p67p90WSVyWGE4JBK3bPp6fJRuuFQ7m2ta8wAzntGYViBTKBpGf3g3SZYrbHXo+KU8fWweqs
Q9+a9mmCUpWGDI7a3jWJYI4gcj6KWN13gEMOI/rccvvUY/EJZ4w98hNb2fKiDkorEyt/jdkfFWwM
SYA1NA2hmFLqS9NGSuPk/kzDB1tPjLgfshmQdEPm4eZMFXD7ztg5J4UZ8l/jQe2kIIfFqqGxca1f
s4KzTnQmqP/FGt3ExoA0wVbEjH2E5CCQ299sud3V/pvSXZhB6L3HNpjoxXA9yuL5dhFokWQJBGv5
pLYY46iNr623tseK/1YV75rf3rBzXFsjziL/Q0kRViMavXkGPJqL9KaWaXtDRrNflK08kKYzrzU5
yahhOxmOZsBKB8rO9QZhVfC9pywm5nmAXPr5aJrgXs5xan1mQMRMFFyK87m+08KwInT/ARWMVzxE
Cw56F2Out4FqlQrvw9HznK3BoA4sat9jPSZwAQUK/Ri3XqoILhPpUxsWccDuExuYoLag3A81rdmz
ZZLjM7oPuNRx8N4a5+TASIyHfTD1h5uA+Ir1RW7w3l9jafiCudwnQqXnQyixTNpjJh90jaxRSGDE
u6QE8+C6CTmBs89YgxQ7MxikP6rb0p8G98z0IrQpOVPeBnY0bi73rML0KB3tb20C+dltXjAWi75p
n8CbKazKO+pfqaUPM2tGR6j9R4I+VF43oBsfzl55viCu0SMHm2sKSl1u+3Lb1CMIW/JQPzcyyHBj
TROkl2/sIg9WgnqJdLO54r5dlKrZpST4YzZtvr84b0Ixbj+2YwJzLH4x+zmjvg1K9fFcR3Sn4I5H
dTCF4cRwcKgsOIejKA/J7J2Thl2aPcEWpPliS/0WdqBgxhoRlz49GW/Cu7e99m7jGU/NOWwGcrjc
LFf8r91RZgmizCupe2upgIZgM19RbmR5ShuQESzZj3Ho8BlVDrAsyL6rZ9zhZYyXau62x7pJyzYS
2wJeau1O86SccqPJHLEY5fbi3QZl2kgie5mURHBJE8/FVmiG0KO7Y3jIQJM2fo0pePElVZ4cInSY
IRLWV29nogFAhFs9ftPFK8sJbDQn6LlCObw920wMWeIdThgO64i6H/9PmiAacXBcIGXSojrEZTBu
xqsmTPR6BLc7oMxPbX9+I2Ym4NNeVQ0wesgugdxaLq/wDOZOiGmez8rPbTYhqKVi1u0bxy//9RJ6
QAxlcxr2CGc/rhLAtWkcj3mSf0fHx+E5wecwN7AH14JjmmMJyGtGEWxl1cPc/24iS95sKMZnToSj
uIPgXWW8XJ5imxtC1WkmnibbrI4h2VYH5qr7LbT4mgrJCm9Tu2bITpKl+3VhmSK/g/pj5Xbwi1FA
d5tTs06o+82gU5lgu5DVBYqX9gQnjNSfZg+Y8WKOc/i+m6aJe/iclC0BBS1b1qNf/+eomHxgQ2D/
SpzCs5r5Sd5f1hNzafDbPir6tBRT1K9dwFMIYKKizAEvO++l4gVBq2dUxCN9Sqcema4k5cYB0wPi
oZUSeIG7ay+e7gC3kbOoCSaf+mZOFFFsIHfrN5ZXP3HA7Jr3j5dTt8c7C75Vjjsa05t6VdBvrLoN
ZqA0DWy1pqASeIFoYvXUmfG0kW/Ssp07nnHyiHh4Qp7PXS9MAA/NkbHtQP4weVTzOCSfHmXE3hQK
dv6JpI1/YjvZ6FRajNVlzeKRnbcMO9ZieJThGULGFJcjCQVFBZM0xQEoMk/6AxZo2PRW8uXZad84
ZvojEEaCGnfYMv0ZCezbJYQVwRwyYQReXeIPgBOiTt7phO14TcoG9g/QlJrjiyJ9CwoQEMuZOf2i
Ua4J/DMWSkG00cxkAMZA4FpELFQpgE5iw5l/3cowcYOwjY5yy7DMgEBDoAercW3W1mNfJ+g4DJsk
Pyj0fcwsdxllC11ACPHQYFqjb4hSEZqLgckyXPLNycKVsBb7jQ9LBIJ82GfIyw7scvKdOdsN/44w
uyTvcX/snIBaD/0yPPHVmfgPVmBaD9C9wko7N8tw1LH/VaCKXXVnv9MhGUt3tN9HOPnoq6ZBrHhb
3IQeawCMLbEzPfhyIWfkaM4zA2/qgHLxzVzZ5aEXt4Pqft3JKrizaZWLcbrWVqUi0dtgbD4CQbJS
I2xIoqrpgKiEjnOxulUoFF0jMK/n/b3zEC55+3WI3hGKumAu98qPESKsy4qIBddR3nRX+nnyXGh5
+8Wj1puCjt8QhUD52zq4FDXTfl3MDChmaaXOraKfBRKdw+mdOS0UPSZ8iVWrNiPVJXYuD0JVhpgJ
X3JsCOmAZE4VrQwsATwtcxYG9fzo7XAim9sN9aayl68/39fEkFzg2oEWd9IUQ0tlTqk1Q0lafDhr
u1rMbLXeoqGvGLDN1ltR1nhdxCEzRKPWmBVq9z3dBApUtv4oPyUXD4p9kaJ0VARdRQsoRXJO+Wdv
XvYLZwYiql9tIduX1bSH8nusZ3GevG9dp2vVTgeTjv5UElXIqh8d1Ub9s2P1pg1999twjnihFDyk
JCgKrVrAKYKzhFaBJSNZlXDYN92rJQmFbL9EBvRTmhy8g8wQlxSfUPpVZeBWFjRPpIflYEG18GFz
nW9HJmKW/sOQh3SG7ltTUM/zd1PfT4RtPMUx3WR6su5Kv+/aEUcyXo2fa5c1lhBXr7ldc8/M9JC8
QTFLE3xMJX/iQktRDxdXFwGU+0D1VBhkBeuRzQRjg7tveKeTz7nhMGfPumhKgscl8Zp5uI7fQ2B4
eS7ahndVLS0SNd4VQ6NkJZQACAEFRMDiW8CT1N5zHK43+eR+aAxPNJBrfvANO63i0Z1G2snwf5kC
Hk5kGBVmqtv3dcsV+zSZVj5yRA3ezJA4DCaEdYE1UE+tyc9UHEKc2DQ2dmAso2zNDM9nRcTEHLmu
RcXoCTJyXtTnlxQOKcrgjd5eWlknJuAAKUrAPcJK76iRpxim8lCJdCtFpRx5P2OKyvOx9aIcgvwZ
JNYbWgVyFnkpA4VQxbZbeCPI8Q2hfqrkG8/LRi1Sv3ebdYQRSv3BEEqb0sX7hB5uov+aA3dqdDNR
Rmx2jppHzBsMJq1KypfrEzX6Boa9mvoaBVGCYaECoD34zUhcgysARk21nVHgioG6eeE7ihtz6upc
SzitW5CHb9d8b++mUULr11m1VmGpZtnI8ceQAwqnaTC5JSO8s0X/psL1IT7oD2RZvb57G9YW1ZVI
wfU34dER2hAJdhsCdX66SgrScYXCKYsMVe8dr0LbINQccAx6yddv6t/6tCSTkcSXe0Nyj+MVOhX8
rnI6KNPoBGYok8DqbEepYCjQhzUC0oZ9MM+655LS7S+6kOOR7XO0QAzj6VloZZ9Q2Cz8Mezk97N7
LER1wGhD+5Ny/NPRqxbPG5Bvo0yAfM4XAxhPkp1OU6e23bDHlC0bLxDaslQYdvuoRY/xiqHeSyRR
56yrcXKAA7c+glQBFJL0XCf8kj7yXRQrczKUl6OegO4BflUv/FjDBN4/Jue+6Zp0fHskP+lL3N2c
4nrarHE0OIAwa3LORXrFvxh83H8CgnvreFhsiFWEvAf0YLwUxRmpLfHosu04VweFQ/6/KmXYw0bd
YfhX6pXx6rtT+In5605f/tf8uwd3a/9n/fX25itwuF+iXi13q98LnKdJrc16YwjxHN/lrG905lVL
iwhwl8Pp07DJLz+ODHQP6s2YQXVt0sTlCtonc0qty1H3Fm6E0ZJubGSIhletUTDM9DgoEDCkVNpg
/zRPLVw/H0qPFzRnq2Ji/E7Ztz7ikSZBPGJIYnipgw5O0G8JncC8N+h/KRSmMYQY715bab7FTEE/
mRugoxYo9VVv9EopEZWpABbFvUQ0Teqma+2FhoApuW0sT1A0YEaDbq4nwP3PNWkC3+9e0QiPnW+f
R5H28FiPKSshGbt2/YQYvKC/b68T8uU2mJ1hE+PAQ5FSeRpOgk1nacMRFLWCebZjnh3eA5t+Pefp
XUsBVKT3/lp0VUQVHwX4DeUnho4a9t/S9PDBoN+FIpBVZM/gcU+Y/Lw3f2eQb+gEmXGNnnhIvT2/
NCYUbG5TBuKlDtWznoJYsuN6D+DEWmDpsctZNQlhC3sI+GDR9z7cSuPv5HAZAJrlAM+nHp1Ozpxl
DNFRo9hCbZZ0XtdN1fHif5MB9cZH/oDnwkEEFt/niT9BZdpkDvREq3MTRQ4h/Z0brkg920H3qyIF
eVQ29tNlXl5V+fIC+XQrtyPHrzFrwPfkLj7Y+ItEjPn9teNYvUgilA/1l6thIoxaH8DvLE8sgFK1
pt+SQRT11xKzj1UYhwyuUZnZCn8AunBfzKuSvWn6sKiUXSrNS3p2abot0Vu7Pb2FU+/vCMCZj/1e
l+O0WpCPj40GE1THH1CjC8pKZkj/YxXLvUvsjM0C+1Vb5vNRRXRpr9SHuhmHYR+7DjHisdT93/gf
v2XH8PH9OR1NPfcfkD0GjDBFBz2orSLSeYWmG+axDoImxoSSYWSFOY5PUhB2nrJlNneseVNqw36J
aWXr1SNILOGOuS4nQDcBrEv/DB4DTCZT0w375QXMFx3lQVn+IwPjExpLQMlcMq5LXdqAA8dj2TL9
fbENnYgEDGkJYpIHcN+agi3Sl9sjtHo/j4s8aBDYaJ+O8FoG+DMEACxvcyKaHCMPNv38KRnsG04O
i5Mtb1Lwpr8ZeAYOOtJWkWoG5xKOXbsuONcuw7f55sTsmC1sPC2Mc0AfpiLNhzRluOa0GtfZP7EA
eJUlL8lQR47o31XO6UgaRYVup9ib04huE33EZQ2LgGAk8Ylnxro/crIu/5Jb0rREbOweDYrNo8nC
n9ekIvV5jSJr6DodmG1xh/KG77YRUVThUBNSyCWdX+LdepWXtc8lfBdMwH65xi6Ap3Yu5hlIAwhW
y+1MMa9vVtmQtFMGVTYeyUeiLbLX+DX2k02cPuk6mpbKT7lvGHXWvHiGOYUrAtulrXD3dgYBUk3B
HMb6E8g0NIKaOcJEwvEmrL9kTTGTvbZ6l8mGLGa9VtEia8DyIoOrMBJLL3CwG+Y4W18pubO7srnx
yBCc5wrK0Ht55pbZSzqARa95tOuzpo8YOVH0WtWIisQENZEou1aCtHRx+UqGC7DOh9vXneY0OkXp
rLOlviL+v6EEFb+Yq5zCLM7oW9n7Vwf9NkLln02csD3nJlmdJK4w6DBa0HOtZsvNdgldX31/3Xzv
ypU0KqU7DGR5MmxGkrd+r94LfwsZWu2zlOcEtIABML2FNmY+wdsBaJHYCoJgDrMPTXhM3Vo5HxSI
KKR4iJPSeQt4UQc0F+usoQnDIzP/6MVNo8n8C7/Ioo7WlbEAUnB1u6KaVSHgRJD2j6Kk/FqIP5xO
Bg5ATYw5DAzp7QEnNF9scXnvJh2+czVR6cwvfJUbgtonIIbzjZxdwzunZUVdXjipVJ2JqxvhEa7s
ABibHLT84LlVQb6MuRC0P1ugF8rP5R3+db6xsEi/nvicXEEhbU+JHJvFgpOL9NzSoVfdtR0Z10cV
M2yW92MPedsyoIsGxaHk5koDIyPV/zPvQjBr30oImiAtyS+7mMkhX3qpm2UkTHUHgyWX19q1ab4X
ybHx3CZNhcnUGDE8yyq0IUk/afdNNOgiSPse6i6wADkBMiDCleKhDSlcapoiT2a+ndOlNQYznfL3
OzkrPNNQI/HnPz972tpNm4RW6fDI13+cpE18C+2+qvDnud9eWKZjHYiKGHYoorMtBFBgtort7PEr
ipKn8A88FoVOTcieR3gvRjHvqGJ1iatGBAnhpNC+mnjA1dXHnhz65dQiY7bpK8ts5OG3FDyKaxK0
g2t0j4S0MX9jp1oEgTFRHGXjJwQNhW5PD+sN2vdP1mUj5wo7TsJOKmqVJOXkB1qt06waSgMxFwJ3
jYYyfV4FNj3klbocqqsRwPNHCVq0qavoovDoErMMi7QvzqqrWI13JtzJ5x2W8ON8Z/3qfXxUjW2R
xoZ6UFX+GPniK2kFIZXy47CW2VbLJOg7qjLX10t7UDn/c9O8bwruSnpKZozGXCOyGeO53kFLMJWT
qM0DiwTskAZwbRaiHuvC5xzlSc8rTICupoSe7sgY3HVHsrE+iEp5ezc3Q1KEQUr48ZDvytWJtEWQ
GVSQUAOt+c5NrQzlvzoeQ4ml71oZYOly1qU9xZFNehs+hZotusDHM/DZVr5i4ZuyCcx5D03tjgF9
ZOxrUrHhvNgbG2Mp/HTv3qGVEMI+PpGPR8ENCLcIozMEiC1q3fIl7pRdC51qC7cWKUrxs07xfG9S
unEU0RWGBlwyPNm7C4loJIcsSKuS2Y2e/zN/4Bk6EawKS6lvjUXvJCz5eAd/78vKFMCSakU/fVcY
yjbTHk7r8i2n2cWHEKv0VU+akpIS2lUAAhaJoXSWArfVDe+DoD7tF377XfyrpmgjsyL7An6w6Zrh
P3V4jmb/fZ3eFSPwLPFPy4hNSOc1FDTOBTrx6QU4LeBtmRE0BN5I+a05pMfxBPQnuhh8YVUOAQhq
ani2Cv5PkW/DE2/KCC92UpoWRko+KVVVfLg+qbQZ+BxtKkOEK5ecFLIVPpInwHF88eulQX/yqIe8
dLPxmCo122ZZZv5T0yHdMq101yrM3t7jIKGuhWgXp1/UKzKGvIB7tN0vg0sMQD4/ySxzekUy7LlQ
QPHTogWIRyAgUao8gwuPFhwSSsF5IITAGVQurqTdcTi5i/qqPWd7j01GhEVWE7A2cwMQwU3v/Pym
yUkcnA+vz3HR0ORwVPDhFQabXOwR9pxryDJYDBN9QYTg8xGk781Miy/BGK+dADrjLa5WibWKB2FS
krTOa4gUEQ2RtXoe6Eh0i7h2b1Afn6npJHBQdLDhtPIQEVk4nO7Ll5JfTSySeGtrBQ+zXi71t40J
KgRrK/9PyX1JG7IYj5+zWLiyjpjfMTeZyFjOaOWEca9dCBTDleW7wtg2hp4IMvPAWIp+P6IRG9Ue
4SKmPBXb11y745U7iohu0cYBEVZIBBwUnVj1vGPiWp1w9n9ZmaBWnC0KD3jjWjNqZJqN6/4xuuew
jCbFXiTRwBKeh9eihvWEsf+VQ60rhHboIu4DpHbEee/7wHQAyVLIpFFzofkbhgLor2TCp+8RirmC
5YbK6xmxj/iaQ4BV9kGxQcrvxNZlQW+XaqtQA+Txh0YlStnBmW7Um3CF073c8T0RBOWH4ATvTsVc
x5Loe84zZZuy0JEzEa7b4neCpeDpYa5aIMJ0V1se/OUBjHxFAdDey1tXKNZat7sMk3HDnZoFihkz
1ndcbF8L+eKJ0ZbCtHtQiEBSieYVhFc8kvNnwogfO26xX01MjRvEYvIG4sOm2N1S3d3Valgj6gt0
JaRcbRPBrgLbAX5N8cRjBeXDaZpWW4DiDXnSbfNTV860epbQweriH4W9iewbir0aM9E1YZqtsMjb
f/LI68EkNweo5gLBGQQeX1djWHLZ1aVIUBKVMOD3HpjMAc0nkfWlXCVMv9YKbuseBvPH7CD2IaRf
MiRZPrJfZ18ZDjU+Twaivcm/Cja7SifINBJgIQu2WADBxsov6u1RCJ0/8tWCy7Ak3YzUwo2qSc+r
RekWfxaj+FNvJqPJBP4BOkR3zW8L9ovXSBSb3LIUm76CRIRoX65JLdx4NLn7Iz3bHKYc4BafPMfw
OJa/Xx0YtgB6cgp6x36GgAuumbPCJoOmI4A4k03K2YqFACHAPrLJckSkCfQ0YzVciVqecp/pAENR
cTZeZU2pzFrzKiwGAMUHQV+4lygK03fN7y5oBQEJGyMDzF137No36N647yoE7pQnQ3Foq3ZXoeFc
VyKjutxW3dSRfnLN1VGr0BfEU5wLIf4sYsmIYqZ61fmcs2+nhwFc8jVQOsSULEl6KJI3TCK75eun
yfs+V7ucW/yK1iNMcvFtA3hj8ivYjQv+Hj+bO9JuY6zJFy1dqNt6jy+dHXvfZZPM+QLx+UttCtzE
Lcw1iSHSqbz0tQbMClz+XNNQmle6fFQn8qOcul4amh3MPy6v9SLIWUtblPN9h7EivYgZDLKmD90x
uRhhtQwunA6P0Wj6d9sQAGdv6uVyMGLbwWrWL/tD34r+WiJw/aGDKAn9O7jGXQL1SuE/5RPKTpKK
rqYNyWZbrntvUKgrOJqcQ7Yr5QCfSBpLh2MIQu7faFlZ7Nd0mDde5C+9f9Z1MIoBdBcPg29tFrYL
whpLvqDetBNPiOEXUAZQf4QbtisUaGhg3zgISihmII2MTBBE37uZzFiUfJj9GKK6iEWHKB4VE1BJ
mWGRh14If3krc/J8mvT7j/DrbvPYTWCJkBpcYSv91IqjXZtf2yMhBBsybRm+e8REi8rn8RpQKvYH
+PxuWcRLBW41iBik0wop18v2DrzQ+oa4rzsbkMM005J0g+fl0idiXNW5aL/W480OpJps1pAWTsd3
Xq/4s88XOmAzBCqtZ5Y3XUyukstGclDN40WJb34Fr7XvNP7Rio8v9wJ2dIJBrAYyuj7sJYWDszxb
vsE541S9jgX+PU037GLTuxGbAWK3iC4+AZ+AGEuhP050aI+HOqX6FfkMr8NYai5HuEjufr7CNr13
tqSdWZRm8E2gYPSUuvSPKMhQrsBVD8kkunjaAyh4OYLdIuKMfLwBKysi15RA4enrxgg3H5jQ5Yof
EOBM0gr+CWi+frI9/xDFgoq1tbce7rPxEPTacwJQjcFKcpaMcdYUddqZ774OmdTwUt7G02FMwE3r
A8Uc6o+uH62OedZW4uMdmBW3LZRf3DO2iI6EmEMtYImZnGFBQBvGpn1FRP/9xYs6TiPOyTFGvzqm
8VPEZsfyWV6qFAuiS6fOdgWtN6/byGHZ1B/N+8De4dv63IEDUx8uItX+EHIJrM9/3cZ3OaoOBU9E
zfSe5X0eCVQcrWqxIbd4JKl7JewkZcoxEiQJkIOfjcSqWImktXqgQjvEf6SlolpVmnVnf4drAusX
1+jJpiq8wSgBn+kWhc2DYNM3/qC61DUNKJrIX1TQJPjS0IIPUOZjLdiwvmz5IaGlx0QQ8HzHyBfa
d64UclcSpd9cmwSxr/bX7SVSfEXV343Q6zX3WnsGmOyBsV+U8lTdglLp/2edAA26O+21k5fJdzOZ
5hxk8N7Djdt1mOinXIMKqmODX0tPhmT0V8MI1xQ5QrVFaayZkmw8MVBlHJLaDpq5IXVsY7udjJkJ
rQcXpycKqlUNXYQnpgDofXZ+PnPTH5YW0G3sgU5HOPtqz5/pqlvMQt4mC4BKU7saZjqdq2a3Qu9j
WZxWTfVkFMMVd/I+m/pya9E9Y2PlHY4tNwf0lPfoBrnWwaYLBEnuPhKiKnA7YpYBCLZLC77q8jUA
aXHpGf+8pNC7+UZ6vvmKQ/fAi7SDn6PqFsQ4A8S3F6epbY5i3U3NcnRXlWfAZf4k4yUJikzc2KME
NnCUc4iJmVylZUiROtjJ4DQmPL8EpXDENDQKV9MTUkyXH2BEEvXJTKLH5oXvsT+yjiSqmTEcaJR/
oJT1fIiJVMWFMOh/VFI7oDRJr1aqLZF8867yOxXLUVW8kLmCnsrwxK+nKvwidqU0pQ2TwzRna432
mtu4o5gFuKeshkpi9llfKGd9zjbjWV76zAnlHQmagIZT4+/Kp8Npn784MDP8lUmI3PAGGXo9vEWT
FJOe5Qm34/qT2GVYHBlBlOYpRS/RpxUX+L+AEPwlm6O4Sv+Mm7BcxHVksQn8ERKu1zTXM1hws2q+
K+/A0Fx7FXVUNBGbdzQYcaMg0falBr1qLwd6VRrchDfOvVW0jS8bkmsITynQOyq0pqb/m0BuIly8
P2rX/oVbIv+tbNFF4K/5e0oLRExxMbfVEDTt+z7VSEU0BJ0VL1yR3e7PLQYpTGnWGULT8LY20lxd
Cr1LF8YmBxbAsdtqT5aG9o7qZ7ImgN6ouP+DetMbrLXivont0N+ScBGz0bJwHAIJ9tb51QMlmXtm
5tfu7zYC5GQqqR2DsPS7K2UNmr5/Cn2rl5tPvacG3EvpVhwgCUinN5oKPYwn8bQUsOg+KdUfeJ87
L3VHQPvvo6K/65XjaI+AlF3Q2EaluVTpbI6rGDVRS4u0CaYxJ4ixcUMMsSNETitwgDvhhKBu/MPN
0gYM42pkqYjfc7GbY29rgqXwhlKKMRC6+OkGetc5OHcZ1eslDHhNmvbI7ulHjbDmFxwlIR0LQhlY
AtP2XhsF8ovvkGiVh51T4g2J2flaqbZ047xKs5nhUvoQVlxlQdu5Mk5ZNLwtvpEiuQKfpWNRuUKN
Y6yQHOFi/xSY+LkNcVTThyoa2Zoxs2MgVdCsjnx6JmsJe2f33eT2M12O6jnYJsdGEwHWtHPU55Hs
qfPAUg0bZGDp9gW7FOObKylko7uOfRe5KCGU2rXkHRMIC/vvI8oH6512uTow4wVyi0qHuY950ncD
y7Rrn2Co3TVjdhZm1g19emWXuTSIAxqwDt+Gym48myhvUrRcE2rvKlHgQIiV6jlOoArbEUVeCdXO
wcHnRbkQCveTxIr/oLZXDQxLzHGCM4vINvS3ZZ3VWAg33gx2jfHGNq6AeILMbsEJ4CcIf72XyUVP
OI+mbhMmptvh2b7gFgvLvMQqMdTZtwMl9k2JX9eEVd3g74VdMFnft6XyAbDVA0dqf1d2kL8vDJsr
2XpORPwvwiGaJBRCNyHtK/eviwFkk6bUrjqx0KDr6Mv4qzOJDJRhcylChH++hB2gWoOCQdvbrg70
/77rqmVeelAakHFjaOLdXm3h6L93iuaRRhS5T3yilp1rYqmslW0lXyyVuAAhcZsyp1sOc3LlXwWU
b4a/tPb0uEhJF84N6R/7vID7IAwgDLcbf7r7qo9Ge9Kq+CzsyXCMW032mr9SlW/5e+hF3fk4UWwf
ZHXGX9icEjpaC6t/FE4ynrpSET4qYE23CIWkCgEHaa5IOJH0B39KtnI78N801GAWh/mCDUW70UtQ
x0jjoHQF7lk2mekpZ1TP00L6QDYxsR2GTPLaKkMqlop8Hfve44MSHY2BawnoeRf5xP89VwTStHUc
KLJ7JAzc7izliCnsq3y7Ch6cjCt6JepJdve2NZ7zsvM1NW/AYcVRwqya6vX8huGabmeQx1XCk7F8
pr5zREFtZ8hOhiu3gk3HY7KkjZxKOK5dHyErrbLzR8jJhEd0YVhWBQ8w2NkJZOkIkHjqrkH9umPl
aiAAvtc5+u2ZSAxvvEdR2QFEwwW6tBniJccbpaLpTWVOJtIhODJsctrXZQdS2upH60Dy2X1vkcTE
WkcBmo2L4KnL0xqeXXEvOXJ4EOKwfcOkCc/3FFYMannazE4Hj5b7U+sRUWkPQG6I7P0LQnZmEr35
yyU5luTXPXg7wcPUDNtsfj7OPcM/G2OKfLqjAtIEcQJ74ojgoVNuaTP0pMY6xkuROwV7mVtfnpNm
664D6MqfXdOU12H5rTnftaumn8M03raYEwUXxf3mpA207mwWI2gA4rBbSAiEhHuDms90adtGm0EJ
V17dO7reAVz204AlBsS9V3eZWSkBwaZET1ApCqLNzwhSmRH9Q39D6BFXnr6H5zOCTqfTanqEDm8s
3nT4OnJ30fr8VxaNM626LI94bJZakTeZ95X2QIMR0OQ58Fv2o5ggugkVLIQ4VTaEf82kRb7ih4vp
WKtFqyNDDwzQDJfjRNmrLXDlfDjy5QlTC11bho0BN5/dLgFMIfTVrK2RYTb7IO9tQ3dGRNr0CNDu
htDF+Dh6lJnvI2nRbPzs/DDQY7AJ16i7UDrzRGPvMC9tVgWvrH9FmSzkwt0VWdciRj2OHfMThZUb
ZD56WumKKib9If89ilvqIknzLjL+YtXnfVFSlwhaZsOR5VnKFza4F+5H3hViENUdOzQaCQOYF0Mg
3yM/2bV3Ftm1PuYzqVa0CM/b7Gu6JaHVy/DRO5b1irBcBMfjy6RzRg/vxNi9t7eRBh7txW+JcG3/
j1ZPfE0Et5zzspVDNdqKNHqWNXCADx+FtJXvWFhy2eavo/LFfQPXVhxAyrfUifmvdQZsHim36NZL
5OMeyjFUD1N1EYNMs1Qqr33FQEZeKcJiijxO3iaG/ICHmtYebSSeuI9h7Zr1TO3Pi+qlWxldyFeL
CzJEGV8fOX0msNK115L2EpC+44gbAZuZGsWmC4I8Zodtm0rEMLLMF9EK4nlV5NMK+0OJukD//vB7
Y9srY/j/rcBbZstY79Lawy8Z4n6y/SbhH9Tf+XSGt4Hx0oywR4wTPYuND7xq+ZtsmuNe4HRsjkdD
OyLwvUlQ319TPqIbtUEtO9+TH/ElPA2TE6ABnQLoaCvF81jiFgTT5JS1jE+VNNo5Fm9/fLqVLiRL
qhc1mMY8a4hjmFZiHB5NTbR12hVaVVb9Uk7+UZjuevvM4bbp/U4wokwtVojae+Rf0HI4ayvBZb+7
A7idUS5x3JnpSGnUy26GHh8TF0+Lq5M0UvNE8x2xdXe3+Yy6bEa6ALpq9p1w35cxZesQtszYEXwj
MEYsnUN/ILQg5+/nACBCKNzIoyUjekyQJgZzj+WmZQll7ieD8/jwLIOeZM0rPP8ykk3i/IOMSnaq
jGQc5Ijhv2o2tHSL5Pnnew1cZ9cq4fz+Bw6y3Oi60sUYIy6NhIm1sHMvfTzytP03XxJWWz/Un0DO
eNg0UNYJ2zJWtBnRf6ol5NbU7MquqK2RzzawSnr70Xrp4UmuALGmMSsN2EVHm/ZoKcVvaGHbR7GD
mMvtMyUpBLcQh/wHhqznSXVpkYYs7vpA+agWXyHer+Zl6oLrGZSXLu2Jf17VtPF0qR+I2rcC90c3
ROLxhY1u8qhRHrpmN765NCk1xu7WGjciwcJ9C0no8p/Ob9EXNuu+/t2b5Of9hw0DfWxYWnZ/4zlw
cQy5Lo7lzGYiIayMBfQ/arsPn/fVNc+HICW/S5Zvt4xmffXlExhzgOzeC67S/80Lan64AGNFTkis
jJW69N3JNGbJ3WDAp53a0s4Ctgtg/1dP+UocW2kjqFXzo7h9JxWNAN5Nfr6+DZG6GtLANuUcbMDo
5LNsoGNx+bkdILY5ikcWdEN80nkO7YkrEf7OTeX7LTurbH2fYSzB7fRgISELfxATVaUETjA9lH99
x4LkAnhKqmoTligCQQBG7yU7b2jjUxnHp2qkMz9BTMjUS4laKdvz0O6UfWUspo3i/A6qKUc/tZ43
Ptq0K7xDVXBZh7rpJkHz8IGx5fH2+a0yXEvzC46gF91btsZdbAfQx/upjCTvnkczBAHhMayWgJQr
1LvBACO5PJGFFweneQrIDWj6ZtZvIcDbmDaj5ACyw2EXzrd7LgWuFY2Mqe7lu+8B717YMJnTyClg
J48o15jmWEqujV/GWM8YaUhrs4CsdXz07JuTGZnz3BzDYSNXEm9xJidi5zuiQPWnyafYWhGQW5yj
onsGsYIHsNIp+2IHNn9lZyMeD3sR/7w6HwOP06iGXOBhD1YLve0uN0SDShIyb3KDD2KBu8qce7Ea
WdwbqXtRanZfdmkxmi2oCrB7tLLRjYCEuk8yD9ik97fjIGI1tO2rztrfd9Bld2vgW5oFfVsWX1S1
gnF4YehlhtnBqjDUhEbUmoRbNmobFWEjESI8kkszCDkVIflEqEXPnWpruvNNFjEPsd7BxVsP6Ey+
1x88+KBljAz/Z63Gmwbx8mWYB12ZGAktuTrj1zGLL0qiJSEjmmcwYw/S1onHFvIpYqttkOHWJ0dh
PDqru4CHmfa16SMQF1cbThcbD2/VsT4TECpfUmK588Exi6PeZ7JyeYDs8QPI6++McF6rbETbCej4
SGrW6EbsDLMa8hmzqDJPliW4xR+MRqbL872hvmu9gHM/ExI5hSNnsrAix+v+Tyjqr/ax+HSHfGM0
HK8SASRxTNJW5fsZ6/7WeqsAmb4ZUKa63jprWqbX8RXbfLJEEkEatRvZAEyyj388WqlYrz1eP21a
2588+oFb1xTbpMi0kzw7XEVSDmrN0xnKuQ+B4YiDSZK6iKUjCXrzf1rLupE/ats05mLVyc2OGqPv
XPSyuxMM1NIw0W2IJj12dDBn9CoC7xg9+7HwwguVOUncuth2jEpSTpF00fry/VZTWvsW7OK7ePHo
LbohkK3jDEqwc5Z7VdelrSHr173XTRgorexB3SfWsOlHkWnpnCmPT/6DTLynMvvwRZeAPArQdcYo
D3vDv/8OM2XWancfjveCN3NBPopCMMaqktd9zRmk2SLrT2Q+OQ2V0rkCdecQV634tVydrwkj04Zj
BhcXfjmiAfGiveg0oqRQ8Mr2FeR1mlKt2ITrDOI3HkBWrSwPc/T4NYVb6uf90qN4SS5t2kB5qbXJ
g/MCREYmD3jT6WfWlF2xo4RjrPFzzKUYG9kBPgeq6UP8/BNUVO6VjYOR3IyfoVU3ci/F+I8q9QSQ
XmvELxeKSZOQiTPxbsM0oyMGCYMnX3elJaBsmsahxvGs+qcsSKtpJ4bCrmtS2+jHuLQZhMJN36Ty
i6kPX8q3+e6mwooexM3m6DS0JW1bQcq2RXeP+YeZ+/Ilwa5+37Oo0HZNjQU0PdD9cJjfTyreLFkU
fZVoSwxxE0EsWxL4BZ3XotCYm2wu/N2CxRp6POflg4IR2CQsUIwRRCdJB7yR7dW2Bu1GgI14RoDW
FEzRxCaG7P0Ab2PsHxkpWiTHPeC4DEzwDrDs8xv6+OIFe9mMc3Xj68HVhjvifUrZ3Y5IYBljFUgk
KGweqjN3PqShvBEslFH2IEX15ebbk/Xa3MUnY0varuVSGeA+fL1TxGwa5ShosgB5i1EPFeS1jSHC
0nYDFzsWeueiq0XRxD31mpfmVIoQN2BPolWDAtp2Y6qHbnSCQB5Vz33nJPxbndIfopJL6d6JWuJ2
9DQ3tr22Y8o3w4+mUtZZF5JQSisSYFB7gQJGxnuagT4lMt3UtSDxFmlAmP20hvGCRYzRW+PYt4OD
7ZFuLLhMbcmZUOD8q2ouJPh3yJRyNTntCNmHEMikNi/0Ru2nwGzAOvzPV8TYke/rE3x4W+jwqcPa
Q/N8pNNEN04t5tSeHCWEJFGpQEAvlFwhkaatbDdaLsT6IShmlWuNrXn7RWd58CKoGLAP1GGDFcrT
dL65537GYh7psRbv5YPcPO+wxeiAJhWh3njTAV9ChhHiGop41m0T/e9O5nFN76EtEyW/pP2OYoej
xGDUGbMZpwCkqbue06QD4P8qOiBz+5QTe6fbyUA5OrWLUie1FMZzrNwXwt7SJDfzMRAnM/Lt11Yv
XWXzchhLolaMnu8HO+yIMAwrXIkdXh4gGCq3opef9l9LlL+7blgHGHopYav4jjgXN4ZTlmVwOmFl
oKG3TbUGSGFU26jAt8fuozjxKa5Ss1BOgDnKeDMfIxT0jNbxgTFCQjSXlLIa5TtOwgBWbXY2VKV7
inDiYTBkdqalDeUNiO8bqtgt2KGHdpuuRdU+csqi3bIhY7U6o7i5sJxzPdDGPTNj5yDuCpYJ5rsL
D8SUDS2M0GxV1nCbY6gIUjzx9+RsFlRzl8plLQLKgzkBMawmA4LEUqML/kl1avG8oIxTz88kgKlK
JKu6fP89D/CjDLqQR7DEyG9xmOZVYqqqnJPmdk8gfLXGI/Lq81EwEjbE3IsNgG2iKGiY3+k+CREG
zdYmnZbHY681VfYbuNrqQGZVcXRFfjUXnnvhU/An/Zfhi4+z7O1lxLBzlKAvk7GAT3ryLzWHQ46S
rvIhh5/7VRt4Wf4Vj0WEX27UGwPitUIJtJTUm6GbxpfC/hd66j3pv5Alk+HDPYbOC+n4Y6AtSNr6
2gEdMlZ2D03olQSmH2SS5yNyn53D182hliJGVJm+mtsPiv5YDLIg8cY1sfBH8aQzNEIbWs8UW2Mg
YT2dWXh1tpxdOOpkTCEtokTO1FA632GO1FjLvnHIbxinWBNBBtxDGDIA7qtyiI7J1JB/M+RRIxLo
13MDD3CIaGRgbnKqK0Oi+SOAp8UjLF4fMDpG4AH8KUJF9OhQu6KpyoJQ1Hvooa22xp5B2q/V8su2
013Bst/DCQGmeLP+o4zF1dl2uy/54yGsFkXPaHwDrpw4S8Y0MUbg6cQaaLBC17KI5PpabeAlsgz2
ITAu39EPYPV0XnfZTOz2P7uF64IhsU/Jtk1Q5yY6KYnwRJA0oedll4UtocxvJWm2QS10MGJTWwVk
+uftygl59EljQfcPSX2gv83W6TssrBzVpWFWZaXrfrczwCaHB8py+L4s64wEvW71Xy+1dvXzdgww
WBmh6BwkoDkPDFpOCr1KbpA1W7TjA/NBRcBFAOuLrPeH6C9WOZdmIJEUZS8jrWH0va5G4AMDzqFL
RFdUdz3toFIvrqllR45LZ3F6FZprGm7CwS+0/YocS1u8tCFF23Jb3iX4Y3GSe5apHrWkpsyiNwah
8tv4/ek3JX2GXAQOdCJEKgPZ271XP187TSKlGraXnmPPCr90NvvqUi9ALbcK88Ko3e489554Vp5H
6lLVbu6CL2Rk0OgDRN3gIhtWQxZr6vvuVHg/Dyy0Is4HgSXWPVYGGf+NMKPwsNIMN+mP5sFZ4Keq
1ePZM54VBaB+O1RAYh0FpaFLu8AeH3SL1qdqdJzkSWUboK79ePINQYVfiKUGFWcynDz/r8OnZ607
nSaY009DZ73Oto89AGuGGG86tRfLPJvON9O6K7kuS0XGQcK5VYiCQ0QJ1R1oSDc6u15F+uAYlbzi
eswWr3qblgpL92wu1ZnVCBxSWBkQHTWSW45ULCoYZ2HPgJmCX8+xZi80eQyDGQz+NLl+b0bmN+ik
didglOg4OmvlehDBVmS9ZbAAPgrWxF25SO1Fw/1ez1I6On7yPdsD1rvrN8NMMk0hoTuQ0g+JNutK
Wx+S4HibACD3s5GHQRWzk70KY0XoM2L6YRBan6ETNmDSm9zfhSaJuaYvQLPbB3+9HQ2mDXrQ4+xt
jJM5kJkAhn/muSHbm5kmxC0cx9bhUS0E0YHssw59LzM6Cr1A4E7qzYYbDcYNnZnzeVxdpzgp9Vv0
nT2iWknvwqKAP9qnxa/nXI+JW+TnqSMEezHD//lOID4ADyDut8yCoRxKaWz+c+ctxpBwHZQjnx0I
H6husuZzR8ZHWQSU4XCc0qscEK3RKLHmChAprI5+F6qBwHYxt+/O3eFseVtEtropVqKaQRgQztLg
I95zR1VVJgbqOuD0f533BA+aoqPFk75WE1xsbbmTnQ4jM1B7/FewSfrZJ8LKQij5rre8p4E5B4Ch
TiSwyiT0kaidpW9ZETlGw4meyBGdRW9pGV6ms4G45B5lK9LzpfwHAJq4cBhE4X5FUviNh/ce1PIP
VGu5dXMxwamXrwOgdPG74OxSviXwkonHzmxo+M31yJD7jpGaJItqA/I1rJR5FnemvyBCbnoWNLZK
h8FjIBL4yIJs0voP2xN0X+RIgg3BcTfHZw4FldHrY4ngDR8ssRMflawqe4j5rB9McDa0gdh0+Dpr
ACcEpu6Qis2RzRjg1lAjHSRpO/22g/hkJSJrTDvIGMVkz8uVyzKhn2t01ZE10FdIpYrgnebKyG/a
qPO49+jvpEFNijlXvanbFwzR0/sEiQ5dS9lgxgAMFTHd682NXgZv657DgiJ8R6hYTtHzrTjy8i8a
nvKgRa4raXO7bm451HANHSdOkN7c7SO7rV8nJl2LWcY7LqCkBQb/010LASpnPbdSW/Hn70fzJ7Cz
JiUsNdLgULcrEWY/bMuM0yh3jE4DmuEa32gs1yCn3o4Ap0RYVnW6KnMhGZFXohjmId61Gh94HVxc
tOWeGc9Z/k/xocVcinQoLYdavVUfGmAAG6S0d+am7+a4hG92LXPd60BMoc5lcybhz/YmpuSUSXo8
a6xZ+Gjo1NKyjagEjEzyB/BbyPffQUjYui56iKE2a6vv/mzTqtqJb3AA8bFwdYe2nvLW9y56ilix
6g4XWRynx7NJozOv0QD7tNaMAtz71xbDk9ffYD72AFy72H+RZP+klTR2pm/wIH7OqEUv1sc+u/ty
dFq8+xqs+Awv4z6/b2u4xqJkdVFRsvhF1y564TXcUuqahqKTwzPy2dzKOB4n/tCId/SYfp0ijOus
NGNnJdm4becCf76oIav2NT8BEsmNGgFJ3ObwOxBU2jh5Tf1k8dmkVqe7rVG3gH+Z7LH5oUyrd3rG
/33B3RZ8ifg23p0p2dshC0ue2RwpJHXqU+V2Ykd48jGSuKA21AJ7AXdHU7jtzur1YuP91tr/XURN
pHEyoLViqUpry0ZZfzcLkVzd3MOKALJq9RC9IAcmJlW5VFoIahIH+0Dh/I8LkY8mRUho0MFkS7iU
RbTytxcyk1QpM49z6DEFHS3vATVEuMRfkK0BwhhNdVJ/CzYTmwRFvTdB5bI03oTMDSNA0aJavxde
McrTuYmOaSgxUYAQKjZ3CR89oCzcghI47Yy7cKIZZRKdu3HtCmyZMKH/8rc37TjNA44yAks/E1IC
Y+xmA8SpSVqilwaNwf/lHzxSYNOvmS+gVS6pL78odTcBYOKIz7XM+LBHnT1xOHT34U7flUUEyHAD
QddqUhdckbDBy3F4b7I7kwU4LHY1yeAdn5bj7Bq7xrxSp7Ocv9jHslPL0jrwR26SgnKADFKuMxRt
xirXaJasIJvW39Pm1awj2gaQmBA05zq/sXgU8wVzWMWlNFuUfRx+oiTIBvOxkwMLb74CaaIQmG76
HDB9EFzE6PlzB5k6ZtSGOmd8jTWLu7HE4GYLO9Izi2iLeP4trb5htOhcgHjeoBA5YaDlEKmxeF79
bScZ1p/czyp6Wy6Pnepoyv9IlHJV/jpuQmBbemGvn+vLGpeC2tdXdrWMqmuq1l9ylA3OHoj+yb1I
sdPRARDF6FF0ALrDjQ81SivmrGhbjd9IR7HD01kOIwJ1OyiU4WnnbZZvlV8NKITea4xNfIvrMR3F
aUtg7su2kximGKOYWjkC/4A7fy7hPkwNEkoVoGY9Fo/7Zcm2TjgG2qZLSJedx9vEmKwLjMZZwXeI
C/0CVCAMr1daK/+O+tTOs+ybyXnN7coQ1l0Q893htwZ3FQj6JjD0rkg25VmMv2JAwhsieJIKQFJq
BlWLuR//Q/5YzgtP2TOKatlHqh1vWZHyd1itYkCJ8eha4gHfk/BnZHi0vfexE+xMQ+vDjryhgcVP
IP73QdU47KX2AKfQAFkqiu2WiaCtY9eVtzxnIEz01lPyT/f+KABIzYzsmBtz5mmrJ6CcC/t3elyc
pYXmeSYOAnLHrPWtJTpcbaBvB8NOFNk4SdG47qQrVH5fvcS1K/CLezSGHvccfB6Qd/Wp3pbjj8Gj
GnoRPtw+nokgW2xCYVc7qUON0Sep+NlKuYA7wQEb8CKAAOT9/usi/+ougMNywMVXPjsCRr43Sdc8
JVhXp8ODOx/A5MjtiLocbeajNdFQ3Z82hnxCWduljTImzYmiGZAos42T1RGO5roZ41ow1hswijL2
cPKB3a36U+/rz77f5r1frBs0WXmhqjigeHwEhPwufR1kK3IExjbLE+Plw6iGKb1uvxG7iGRu4Pma
LsJ7DSBfoTdtHhy70a5fMB2JrwBXa/uG8aR+HtiMOLLoJrHep3fOmP96xBrPbjjUFqote8Oe4kBt
eM+rO8/T0DFfg70tf6AwJrOiCxUkYtG7QOJogLBNzd4zWdI0V0ZqbrQMQF7/8/Er88YwigQbvKJM
ko+95pHhicdR9I2qJ10vOzLMcqiwjEyQ5raFEt5RLBApKWiQbwFp/2qOp7d3a+YTfUsdeBhpbzF2
Z7mSYQncHCpKLlgKn6ZRcud2Y6xHMmwfj5rclghvWrB9gaGVwfrw7mmpezyd254W+9MtuZTTAZrh
AsQsbNebmHn3n9dX5y68TeOalLqzcQEzJvam6lEk90xKppdxlSENxoCCP9KCOfPPt7WIB1/7YDJe
6/9gLpMKEpEccJGdDVqF2AMM/lfm1ZsbA2xAk79P17QprTkGycFrh6i/l+IrO5z/+AwzW82c/rdD
Z0i7l9qXgNf5x2nwk5SLLZub6503O3KeAmorgh5wqG5M9IHMVYTbwPCosEjw/Gm8u9F8SQsTIFfe
8CaQnQrXLCf20tusULunn4kOL0L21CrlmzuJllsoEGjS+6n7ROIgoUWDecius/UK1QpzfYmFTiIP
1NbfqtQa2SJqvBNA99FZ1BuEEaRICSaRn+SRzKW3FuyOrulAfPDgmjZ2Vrjt+AFL1LvEc2gr4FAj
vhY+wftFhRRVY6eTOrPtWxn4v6Hs97Z0gIkvtx//0xfSok03BoQp03P3alCz5LpD3gCcsR09jd9a
0YLnORBW672InTZpO1llnOw5sXbfviClaL4ObVfLjY/taKzmUrElASL9uJQqhpt8oPKLBgk73AHW
ErSDd+pABgOm4+VUjtTFv7AIJKO9hehpT+P6tmoc12UAMoxYVKhUL2UikIvhHhL3R2r7JZYam8Hc
RHlS3zqhkHWyca6BG58r1daZ6XsJhdJceII7198PRSKtZM1uB93SrIH4kyZ7v6WRhEWpoNKos1R1
GCD+Uf7KajsSMev2jIIP58NLRmKRp0Z0SPMl9PkVq4Rr4lyffgtP985FXAnzeYdlLJqAK7jiRi0J
XZqNqTSkHPl2IaI0ESfhunAWWkQ7yFcqbs/0DwgJsr6XiWBnjn5EKJFfa8M6FsEK5L7GHpHBF+3X
WltQ4rfc+8W0gl+BFxV8tinNAg9vsSahLRdm/z17Ugk54tOax92gmaFgarDBtvKooRNVgCmeGO9r
UbFGrbP2+em5rNe/yQnNAE+ml9fCKwuMEaF0jazNyN5+CNEb50xcnvXMxOB1xZNHl85ZTbhkKWu/
yABloa0WJnAeF8XDkuqSrIVL9j5mA8IUIhuHjVA+jyqzcO17ySt86pfUmQT/GAZWcJlYUmNj0TFA
i0hlmlljZaR5LV07ZRjhqnMwOhgwBP2zJsYEm2cfcsduNmTsG2h+504fo4PO1PNeoFLI2FSzo/yC
1nzzwGPEXUYVyW1WES3knlEhQP1xDHE1Zm+lhzQn9NyvVY0dWHHsnqThmxgk5ruFnCec8Rwtm8Pg
8sVEU3Be/x0MyIY1GwQMsnmLMTngYo4THvDlwUZa2J0i8WafeSXhf34URbl6lSHldSo7E13qWLl4
+7HYLS3s69AHvqEXCW7XUCWuPu5Zb135920Q7H+bkThm7QsBHsYvu3edwyopTBpqHVbSkHKJA7fA
PlTp4wWS4ty+pAhW+bw6m3AO4PmjYp0MCJIfEq68Zg0H+2P9rDBSQ6sacZ24LKbswChyFDlyXV2T
X+NKjBZBJtquNGoYF96XMq+1yNJfxNbxaiRocqAmSrCak9Yy4IRpQfeQTWyDpRD/occbUvG6j6aD
utPk3H6xDeugt4w5WejLP3ijAlvD4ej9jMpFMroNueLaT7kKad5sDwGt1tNfZ8Ec2GIuNf/Pu0oO
0X6ux25QhgGDwDQzyyGJ/D7mNcwHI6ilEyMhgQD/xlWOul3GxS6WLXK4ZLtQTZB4ssWwB5DOW7bw
+QL6fg895KX8ufBGAaPUiCpr4q8Z1xqSAEXdE7GW8QZAqqj+F/tiO4Yju9Tomv6f22p35MbWdnBa
5aIrrBkAQFrIyB0ENf39THH1c4i+HFO7kzb0dDBlPE7x0vueh/8UOVAFQ7vi4UdM5vLd6wP8aRnI
5CNLFE6waz44rBIPcQxjcW7EFuXPB0PWmhsuyeZh4IUDilFxHAz24RIuXJYi0Gmbf9SVyA2RZjvV
jXWgy5rKuJ+vy6gDOJlZC4gnz/UWmSx13GTpXNb3tOZze5bG7fICk3E6k6r8qQaAkfpDGfHXdmsM
R9bLz6dhQ+KztPPm1/QCl5GXnTJ8Rers2/JBTc+WQrfI/0L0BM5wM7w/ia28L25HLw9nZkyz+zsQ
ikvsSOg8HwFTx5CqL5W7W7wZa0Eaaj89XGoOsuahsd3gdT+YefqYMINcr3gtMz8RbzFoZXbVQZq3
uRb+isUNV0MwZUDVInYROJ0dw6gz2Q1rzpTWQ5Owy7KlBJ1IKzBSsCd/T0L3G0pZ83PfcvKFhpi7
IQwTBjWTZiejRdpDj07Gz0vdp0uq5A8XaLB1uBBPn0zqJn+GU2R/uGHgtWS/RzB2UexIqudzwiVK
uFmsvBlVuetiNiDXMphSmWvhiBDciPaC6ovmGPFMTiDwFZvd+YbhyaGOfybwWyvzeBrDmh5zm7gG
h5fvcuVb4NB5AzF80bTgywfx9t+73Uunz7dduRzQjTkGY4AE3n/9rLYqk5jrA6zkctVh3U7v028y
fGaJGB6vmHnEV/KmbiW9CrH+/yC0slY5yIgo9Q+nPuN7dquerO62AO8Ut+Kx0d7Ai5zMZB8/6jFB
wS1zkxbdfmEIqZo53vYjG+LFTLCpGMkqc4wD5oXKePObWN2635ZwYUplk6X2dKSDug7v1gqSqoae
7ThnuXrWyrFWv8mBwW0SeO9oqJTi52UTFmUXeFRCBjW+BFgM3gMAUKnShYrfbJhX/SqG8coQ1Tlq
OGMCqkcqZ06ZwCuw1j8XqjPY29C2FnekD4FUNz2yYVVfNoWInH4TS0OFKO0mRYn40H7SuDQzEEvX
CUOOOfY6DGhDsKGFZtg5L6AIWFWS93CJUtsMXOqFSzvxuM1JyoZNH2yAM4FwF9bvFg+cHoSNsAs0
ADzYTXXBa8KCwpDPZGKr8OqdMDEnidM3rNXzcLN9u8uDvLVU/cYxPCG6gFRCbB4yJjaY189n4XCo
/xcHFZ6C9oms4XG8XycS7smciadIQgOezBlJs10MG3+SAsPUZ6mhERf5fq60FzHghNDd3WANXEar
1tg0OVyMuXdO01UnKiF3CElTIs9+0BvmmmG23AcS0KPGE3zzxlnqNdNRSEHyBcnOKMwMK/+ub2lx
+6LCMqwX0bPTT1hHZJBmZ+K/FI5etyXQ0VkFnhDPYLL7EgER7uYmCEndfXfxuBJ3wqmGsyIgL09c
8eJt0nluL4PgoksWHf4QQm2oKkAxJ1J6FBOmTxDzANfrcC90XOkqgGrmFPHxe/OKfZ2b63M96Npw
vvzR7GCZhdV08XFAcHTCGWj1LL+DqYurhajS96zX77lOQkzsHI43yTxpXyqNDWdZ64UkyTYVtEyH
ej0X7SK20G+xVCfBg8XGS8uEb2SMErWunpFXVp/Idq1kZ91Rv7iU1hXrx3nVRztc5FT2eCzSMrca
sPxDm3Hqq2gvua5BTegEF/SkEp/8PnZpgl7V0U9FWzFbV0zs1li2SOg2sBWFtw+P1EYCw6fyB4ec
HRbadsTi7PmWzb69IXcDrcDVP3gZDgyDmrxpzoHno9o6dnGTz8wGfIhn+/i/EYRKY24Vlstr6TV0
ovbi5wrgc+zKfvK7feehl7aNbjCQuyCsRtxlzkC9eEFBsgPgIm9Q/UoDYlKnIGul9qmvhtepDyYV
axnSgxbAKafvQGInljonEIfrH0SSApZ7E1n7y8lFjN9tJbMoXvjgakzFAk35qcXEtqzBwisTn9O4
myGoAW8XErE/Dimg6/mADU9yDM0ve1q98XIUlvZNYJNgO3jKweVjYqIdcWcJUQydUfurtu+/jg4Z
Pis/Z/CHr0GKxG7x4jrOG+p8xcMBRPIEhYoJiWKkc+MFbxxQeO+k2B1vmiimuE/o+UDmpdxWCLW2
OVCbTOMZq6WBBd8/dHGmQg8Hkdb1CMTxf5gZzaLSH1dL5kvNc2hQLEnzSJuPtjL9ij9Wdirco9jE
CO5YOUAQemzMad4jzHnfMk+eCQAL0OqwtGOn/Ni8wsGr8taL/JBSCAAZc5ebsP7RfE5x6sTt+5zI
Iuldf5fpY9rS/YgeXNkN7ZRr510z4XV9v3fn3LfufQk7KYlMFdGu/JUm0Jr3KprkhHLeAcq/BXIC
mWoJ+mEo9OdhfSzw/OdkN3sMVbzrk7GitNFc1ivATJGUxjE6+bDCSFiO5HyDid/IeWca86WuljzZ
Hj3fkHnBqDCa4Ca1JgrjMllX3yYzbsbno9/NOPCuAzVTROAIo0crZ+5Zyns8P8tj1w6jqvW+UOu9
NquduoLmb335Vupe1kFle4BSfv38Z066z2vg0EpAHb+NvTKLg3pJlQlU7SZONUCzyplS2oXmIvk0
Nk39soRtOtEZW1rccDpHpA5EsAA/iVXzq5sAERA1BfZVDmjcs4xKvAfeHbWwdIJ1JxxDGjkegkEm
dUCdnQaSSK3ij1EeZbi9f3y09UCQZkUAsNYwXgBIkVGzXI21hlxdQwizwOGy4Wy1mR8k2IBFIVXD
C1/N1p221cFePboMSmZnVZJqx6hLuZAi2EiiYOUWcEnaGM99AP8OydX0EvgGXnEpFQ3oWZLXKJJN
WNrV7YoCHe4h0t0PitmhXVlWKi8c7CQgsif3PP3KeL4fGxjgD6XTpLBZZ+qd0g9nTiq8XwbF+eEZ
+K3cwPC9S271Wp8NPKFIlrRCwav0DkyOB56HuBd0NlK6lZYi0627D5ut2J/hJPJs2tvlTSSbquBc
yaSgVWX1fL29E3ClgcWhD/lbo1szzaTyjrTr1nWr7YlfkB2HY8DxPamSk+xF5s9E14FQeUD5JSAO
LjraOkNj9poQhhv/RIZws7mDcxHGr9pq+CctvcBuYVSmbcHLZ3c3toVigaJwkdZgBvGWwHTH/Q31
cFZArJszFjZlSFk0Js5iwB8UH1jZ7iU6govf8RSuXeqmiOAcUyU1afpSFhaYgbWXeKbnz9/Wld58
lkIILfO/Hl36r7HTuv/0Ns2mtelSftptJKaXy6jlMO9H8IDnMO+h6o64MLgQmG2hwChzxPVeZ1+A
nDB+O1RsDlWWgp3SttY+1hawDZxCnAPWN2L7InCOEK7H6zDN8FvBhOFJsQp2Vg/v1sIJcbzrk2qe
uBtkVH3Mjggw5+rqN5JHb98lGUaBwvMtp2sMk8U5WDhX/rZGqwctXJ6prmN0/iYEoSzxDG+E0wpo
3iynvgpRjNTLVLT7A3GmV/y9LTLiwHKAW6XXMx+ADwEKQFUStCcmvW+vc4QYdJsCQvqfaTjWQWSo
HzdjJPix2QYfu+3V7JVFbsF2gTG221ymtF+WYvUy8MkI9ogMHruupB+IyA9WFGZSoM38Y9WRRb5D
9VBpF5IkISR+EWDhDXZOv06Jl4g12b2nkHmhDIR5dFWv9wDPCaSaPj7ULhhMut/U6Hqrj5hXEvFo
fadf5ZnfBx8kSpGLNcp6YGb0nlpZmgrtMhfDUigYVPJIa5hTSjVB6SpBUlHfSvk3P+5ztMcOqSsD
6/WinjoLXG2o3JhjsGox1qq97eSrp2TVvX0TV6neHCV3fiBw4xrwqGy67E1ua9fKhkOTzsoiVTcf
bpxZnKOd2+vKquaURtL1+2ih3S5bVMzVKKlqh/7T9efwbIR9DLAnBcpcQrsj0B8kEHYb6r3OKYo8
qtW8sNDOG62pt/6wPeZkGyGrju7StC0GWwZx4hwJuBv+iaDmsRI2XNofoJQK9WuWa/cszJMc3Xai
cn7kVa7KI1rW+E4dGznNdkt0vltNxqLIi/9CZW4RkDNly5K4IxjvQxpFLUYbqEPlW1Sdhne6BdNt
RC+jEqZUA8gaRfZn2frr9sMz5yo+PTgdbp94g5rXsJ0kl5XT9zswiKlFnFV1fWg/mjq6Giy4jaQD
0H81ejs8eG9EhamZgiNDPWH9xQNfMnPntBnvZ6apWCs1pY8hR/2v7Gj2wPkVyS1Esfi3kaxt03mv
2YQf678DbZuTTJJKLVVZzAvLZBSbxDvC8lyZTMhrQNK1pLlWJUsl3/I77+UU4eK+4cUxFj9r72FL
NsnXhhbEaOkuvd515mqgG4IbwRdZ54EZ2QIKVXOXTkgpmeOr1WSJhkk7VCTlXG1VNl44SnNixf26
Slrv3CbIizBXvzfprQvxtZPhmzU5wHDOTgxvlUqxsXs80JBBtGXWt71w3mHvjthEPHnuUIhkNtRI
yH9s2CSviMegHegRdtAs2QrLh2IECes+KArFVeHsq93zAM2z72x8I3hqBYBD0BthE9q9FxoZ4y9j
2XV2fXbO2oO9Qi2LL88+RFBYiqYu1E9x3R4iKs8luxZETq1Tu0YLYz4pqkl/WVV/r4ZWFtWocqwL
pMXLQJ6YAYq5ow9radYtaSy+glGS/6ZVdbqAAgqiPmB+sssa6nf5u6IzvY653g2YSY4WQoGRH2MP
R5gGsjtNXm08YxKobjIUHgO4nBINyjJEyNkTuVklvIhw9jfdKLwaIhtg4GQvrn2TCKHJmTTi8ia+
qK8kmCPsEfdbyebSS6s3j9cod8R+OvAKAsdADUhPTnic/fBZ6HahWsblL7JaIdRrX7Yxv8GN21UD
o083/VCnIRDJwnK4VUZN0sEamLp3WllsMTl3HUhmLOWpjVpXmJW4ZNGSSPJowzirTN1tYKR1T0kP
Qaa9Sn3O7X40dThMdqiDHIp7/QRFjOMK4/mXfF+o1lPHm9Ss/579wjxWosZBMohXhqznKYKVIGX3
t9bmL/ac4216HEZoqZI8ljnz+cPQ5xJY9XMRIYQSLmY5N+sCV4WpeRW08MKC+o2HUGPjnZgZS360
XFn/Vvf4betuXA4FWrAlmZ/1hD/MP9pdo1YMy9ts6n783eYYpDL8mcU3IRiKDj8m9xpidaPhGlQ7
TC25BXGdBJ5h8wJ+d3YcgDnlRHVSM9BslPP0HaLAETIwe9LnE0+YDEZm8zEofslJQD0jcVJsaPTa
1sRSPDsjUBuM70snAq3Ja4JmBaTIUAJOM1avLmdB16zOpZRAay0FPdmzNwrBvQBkzcDD/Z8nZVvV
Cly5PQZFDwrRhi4CYitKhxdBcDKgjDzo/6cqRqKnhepHBrzakkyYIVHuqMr6wqVDg/pL8DSO16rO
33aOH71lm91xvQLJ45nsZiVmAC6kITu+uqM3+nwp+8PTlg8JKTKfClmbn+5YjeB/Ng6Ayg3I4T6h
O5hGcH7GKFimnPORMw/v7OE9JVQdqP31tUADm1m/0Ucl5/+iP9KBJ76vOD+hwiw37JEYDHir58JS
5iQS7PKdk1jW/xVKO373Cgx4oXrNAisIfnszRWR5tpld2JsF7Ydvk9mplVpbTm+p/SWjB2Bf07hE
yHMtyXGFQsb0CTvUIEjeKmXZs3pjuzECnjzuEEViTJt/tstdXsKJDM/0MWSlHzTjfZwvvCSmnvVk
YtjyvQiPWLNNatELKOJm88ONRhNR6egpmofjE4SqUzHswztNs4OTCsoNYYPmVXQB/LRj5eB+o/T0
j0+s8mVcbuLwUk/A3oD3s8FfpVj2OGAoXWOaLcnTV+Mv+chr5Lk/p2vMNnPvOoyUpCkeOvB7i49o
UyZCVd+R+VWTVqx96xnhEhpQY+ofD2wwrcbT7/bM+9ZLCQLszjFSpso8QfIlIUJ73p7LSUnEW3TZ
FMFihs4+sSVj+TL73SqBPBqqwJ9UbPbqwhqxvw7loNrAUligHsrQi6eFoctppEZP2XpMEpGA5ZhK
Rr6pIz0Kva7jzsesuGt59tZzg7T+t4bal1fRUThFpBGgPwgfluwoOYrIrRMBWQsKqQ3nex+0Js97
nRVXXhCaLXUr1JLkvENw79pGtTAURVcii5hpFqOgh2aoJfdY564swsz1n0CTItYmlZ+eRza+Io8M
fseCRI3rq7slJNANDzSkxoebiKrzLrHzx/yvfgaKyWpRZ+sLhIj/O2jVr2KA56ow925+nzZSbsnF
9TLb+cwHpEEGcb8gp9e6dncB6HOm7uQLrxikTkeL1/G+aa91l1ZXHP8IE74jFooPldQTX86Sryia
tt/WBjRiF/SSKeYw/TH5FPtRhlByJTEPHZUoT+Eez72GiS+NWqu6exiYlukZU700TMSjscCbs9pn
fJFl3Zes33ob5nUSGIX5riCrzoBQCiVtmcd4JPk+xvIsFb/d49/fxwy2bJyPEtx2dOGqdusXkW0n
PK9XY0z2ocVfgOdTLnvaFbZw6fd0Y7ZRPChJB2WArOoahTXK0xBD3WINF8cesoxNPBXduZtd5wO5
mjzvnodfHigAWOjSHA6Wi3fsA0P03l67dQZZ4gkil07BFYe/VAQtZ8oiTjLUJFzbmZxyg+ONw4y4
CTbhS+EdYKUlDhqjs9V6uaWJEE3MUN1aA5UFWtWjn3y5r+yyznPx4Yzu2NFunBgEbf/UjJd/Lh4n
QYAhp2XH+PvC6Nf9wD1R5jhybM49Mdv5pndiF9x0PGwPApG+l/IDP6nQlsE1mVsMnYXKxhdNKlB0
LCrMiVkQ60stAodB6NPdpJiuTybQKkJ85c2+sdi+8wiClmkWQ68k13UwEJxz2SPk+UnM3FA3I2Sq
G9la/GTjGDkfjr+LCg8ncOXFSTDyYPMqnX9WM0wvuXoHl54IXrivHQsWoi1rUbt+VirZRxAeOjPW
tA1inBkWGV6qE+nTmYVJttWJ/arxRXy940zjQkF84RYqjLK+4rf10f5O//vS20HAxsZIIt17E9zO
d+svohDb+mIzAvSNJ5aoOqGGQWKAoeWnvlvBeXYR17CBKvhCDHXCQUd+f9I26V130KW35wKes6lJ
EdrFSdSD7692YsrXXWa3YIfcjaXAVqpVLRiMSdFxrNBVvLXhpWOSWKMdbF54ca5V9BsPT7dj9cq4
95JtTKCUkKlz05hyIPiw2GjWB4951rlV5m/pcEQCEYr3MmkqW3bXLiIglK+5S6BMYbPOtoN+KUJa
QFTbyEtTDpeEBFiCKSFryqd2Ca1jGBSFsG32JSKP65i2lxQd3YW/7lZQrtS+MJexBVObUBAzIZ6k
XbtqY4EltTyltaHxos7r5lGfxicDe1w0xpONzV3WIoMeeDi1ZkJfxMk6EkRKuki3k+n1TCRtPzkK
MwnCPBP2rigB42E3tzwHDgd3tFd02Z9i9+taW7v0K/uwbwfF2Qq+6RVkJJYrNm+fwKg2g0l83p/h
HyAYVYRl4HbaYVrY4d7UDTc5krp1kFtTdAQxLBrxuqWgnkY8BXFhLBIjRx6GWcs0U8NRfx4WMhqn
iMSiMiznz1a5j/vYS6yGKpXVLdEaHycN3YIdptLmfMRWeV8TcCC0RPla09qDptmUOl1VmZTeGRpa
3D70Nt8AMc5Xdx/5eBo7ND4/oQ81T7NqnqhffNHq7I6cj0hCuviRUA0Cng3gkA79FpLAvCq0pNGP
McVSGEOsIWvTwP2ozXDnbtaIsEAOSR+BLBERg2mldjLEWtDcXCB/G6Jpd/UrR+Zm8x3bA/JL2dAG
HjSmxoEcYwjHa1sDsF+FzRB8b8Up6QAqJ9+CA5CT4vVBRcQ3Ejx+FR1DMIakKHfOmNTwpmXoTVIZ
mj12dpKmK5oh103pc8GcND7NejDb4bz5JyPOW92CSFycPeqMGHU6icGaCJKGduHTi9sCH71eFOmB
vsCWiXCg9z979YAENOXjaxG8LaG/wX2IoiOW1k/GbevTUoc1gBdQh/A+m8+Si214ohIIjLorIF+H
CVDn393tw8NYG1cA9yQwCJjAxNZ2kHv2rBI7hJHOe1L1eMbptVNzVc/0oKjEhNfLz7ZFV9Yi3LJT
ywkrrDwSbBqXpage0fxYS0DqUzS9Kitqzm1p9QTJs67yNmfpo7I6SOFKB+kbq4IyPU2DTAwcWZ3z
0SoRZPf2klwYhrFewrw1JFaLGry6j46mAAnEAqw0mCwh3t2wGa+9yUMZx/UCxIHkhnSdgXake00v
0Z3CiQvnvL7IXr7nfqgcbLqAujaFizgBkLUFcCLQAy8JwrgRg5sYO6dAlNMr9l2EhYdP3VDgYhGH
B4BpysTW29dcOeuQz6KDdDi/r+RF3EqwKY1MtaylJaY1sq/4Qbdgm+OiqkEVLRP3PZpqw/90SuQI
cp77U5bBl+5Y6i6UTIsw7sK78ePMKqGGWY9NIHc+4At21LxVVjcsFPhi69jBkkaySB9Vybsa7D39
jkvfq771VnfRD/NCABu6BnZMPD07UCYfjobrxjiA5GlctXdIfeiwIQ7N5fRCm/biN3ZntqycJjwB
6D6bWBS0hoUqMH64TrVDaKGRKQ3n3oxPJZGevHlwUEMrozJt9DEyDO4BXH1mYa0Wo1jge/1mrtfc
WgKjsz0ZG4EOUrd/BI0boBvPNCuPgaddkk6qN+eaR3p1l3CYcnph7Fa3MJkZs5wd5G+wGnzLwL57
gMSxXAtBVdgBRyV4jwpLNRdogUjNi/FkkM7dIe3nDbm3p0oVMqO8W2W5Dkp/zcm4WgT7TEf4r6cE
lHK1WM0rGdJKaoQWcobbIH6OGvwOl7cptV+3UEoOaiwyU09ABLJPtCAOReJFVc9DECFdqZicbPiT
gh4D/eHt5ADgTeKf462GZNcuNWTdtESGCGxoY+4MNrbnQwEyBDtjuxG5jzwEKSgyxfFR+T6NebwC
Q8yHZZabGd9rE0Yg2jvsG2i30g2w/0hgeNdAOPFBqmuY9/bfTnOg9WvZ7DaFJJiyGliPDL36YSmS
S94EC5D3+8Xzt1R5fYJxI9KWrOUNtVDgDqxIYwBl01AYVOuxN5DmBntaow4sYGod12VIkywsWbr/
8MdOY2N34l9bFHrhncAS4QK0t3rXiB5uEHfZhtQNvS1Ww2nV4uclcPmE5uWIIc5fIx2u5hTK3biR
uHAWJUBpA9mYQZ2+rm0STrc9ELesTG6CrYsN6K7zs/FHmiEHuBbRJgiHxq1Y9Z3OYeWOzao/NprJ
8xBa1uAi/eMk6rdyLskyG/z/YJGi3i/WAtI7JmBgqdHn3BE7fndnxs+zRGnwunol21x9dNc43bLy
ejUzLmup7TmwRW2OASy+Mpzakh9zPaBFj6qwmJoiSmFk800po0/cKI4V5Ze3D7Pqnz/Dm0598YzZ
IbwmnWxN8mOY9U9G1kb/2QdwUzk5VEttBF6iKS74DbAVyBSxnSt6bAul5t1cQOvSPtBHU+vMQO3F
/IciTvC0MXr8AixoRkcKdI3IMZXDE5h82hKHmlPzV8KJKYhCXDCzfsei4cQSxRyGoTHLLD8FVkrk
gNiUhBM1awtIq42hRTEOlymDuohIJARorW05f1ZyYDpM61I0jWOqT+enrhZyEqADCo8rUdS2QBSP
qV36A9s3xYxTRtwgOlhpG+jd/GjOnRKxzyIlHgLWNIZ9F1jqFyy8v3j4A+zgM2V4//W36qBLW+gF
3ZzRpVsF+2GbDet9fi+N7gthMlT3DfjR9dK/OBl3O8jTtC4xYAv8BXoQixQc+SmWFLHO0Pd6JXcU
4CbG24D+47RjeU9CxscrsVsLBWEkZ1L/FHA/AHQOhhb/wqnbUhF6uzpptafBO2+qCgY5FNAfjVQY
Av9zBhF3qNNfC616PLB+O9PYDNsbApn2cfsoppMZu4aQH0g2y1X0boaNrc/Nb1Ie/q6QutbaHgpE
JzwWkTBKioCTD3EbGs8j9+agbEIQlyEF9tyZkh4FXjsURhQhcHzs/M1YWlEDxcFyXi1U0V6pcUkD
2bMPSmptfTtrysdnr9KuGBR/oR67kaYEdmIg7FJNoW8dUrvv3r3eo1eMJWW688Tk3YFsfac1g2d0
eOGjNkQygQSmji+/0pkv2IkNSMgzLKHnp2eWx9M4L9UT3tpU45+TN+LRs9sg5HFqVa4Hngtnwu1D
R7edOGBFkp/Id6lNM9REjlmA2XRufrqGqS50CGYgzSzZJaGG2kgyQWG0qbaeg3eEKOR176Q/P8EG
cN/EI4oyQgh0s45v5hrrbDXGoz+3AMzPpNgVYsGczME44capYmaif1n82OeBBdSb849jERODw+oH
vIhwiIb4OizJm/4svmFvlXN5bqTgjOhFGHO8ntvBy0G9GCc/Uk77FryVqqf3CqBhnOVeOaZVb5el
74AgbH2S/GJwtEfjt3nuIY6MsGVGerzYftgRauEUYPXkaZPAvk8QyOArzDH5OE1/qlBYtgMGvPHq
CzK5u8ieISz7CzOJjmGh32a3sclIzPwqY00EZ2sQM7bemF4x9ceruKjYgbx4bnmSjaTtBHtkeQaw
8WXExhoJw7b4W2EivgeqmV8Rrfa6zyqb/cxgG709PmCwxjIeQ77i58HO2k5yTOjYnFtPKlI/ag0P
nYDypqyRkXBWI8bEHitXRazeguZ5UHWpYbpxhwbZex4IRbJJTJkCqqzZ6Q6DXRYETEW9C8rlC/8/
ow0ogMFqVr0uznr9OairWzDYfj8d7bVZXPcim4axxwI9WPe93qwrrwsqT22SnvJ8bBV8hm5GX1YR
N+z/TKYHmd4wMAV0GGVrIPzjGCUcqqDWtU5FJGGdhXDYQMSkGFg0iMF4HWR+z60EDZKPdl/KJTQS
MMKFnJdWNp8OYezr2j1gDQgeLQCtEY1ntxv45z8FtgfWISdgcFZFzBWMV0xwS6F1Y6MzaFVGyCwx
RjwB0aartKs0IbqB4WsjLAsgQIj9HiNin+cHHB703yEVMBPS4Ln4KNAXVC1XTlh5rBLiYe9bULuV
VigGr6rfKEhG0JY9tTDdxJUCrcQ25C7z6GBDhjet/RgHElaE0cisUQpTcSRFBSWTWqWEN9E3cd4U
S2zAW3NMi6m1tG2ZS0U+amQKH8FBkbQdOutqXI5W1if2xz7T6PKFMTuQN8kmE4YA2x/KCxlFipyQ
hMyyH7lHP1bhpdr4Rf6Vkl2ggpn/MYrHeSXHai7Mlrc0K1eF1jzVrBY6lMNHC39X57NrqO5RyZEI
WFHdDx0H9GAyhaCHVHJt0Ogt9pmI9/KXTokDLAFVhk82hcDTfJDJREiOjLqpl9tYOwGzR47a1kNr
KUEl7yNuhjQ7WbKV4eyhhi8NRhQILNJoY2tjuv2npR0EKGm7J8i2qb5V1ukiCw+npSzVg726C3Bp
rAocUXfVWKAeLJ6gmnngNSOAdSLOWQLSaKzOnlMdk1y+UdRktAgnMSA4vWgXLm5vzt0DbtZ3WifZ
qWz5ttwX83lE496ttUSgoSrEb5HwQrh4FSrPZvpKXCAZtrXV8Mq7LcIndcuvAJhuIL0tYBOpjU3u
VpSA3XrgdCyzl5uE/SDvLPLVr1ywN47V+ye07yyjNL/EBCpsGvY9ZdAfwsBhveRXdQ1fJTra+c8K
W89cqlSSzQF31eAWQC+5PRmMzUlaQIRSlPUm1LahPOsESrjzi1oe7Ka1BYOy6j4Dgx/YavAQJ0vt
ZEEPd87B/1lYYBWOPbTa3LT00vM2afVX51G32sMvaZKY3Eh2a+0d9tH+jZFdlA4R3TudzAOwPa5M
uC8KLsEL/GgntY48YhpDLxBjS1UnYdwo5H83AT+5iU4Ef1w5Ta+k2JTYElaIPklEczVcZ1D7vC/v
lbz/PMPMuvQefOjK532Jjnf6f2K7s1qF+dQ9FpnpJOEt2xgW8kLEoJ97o+m6A2yvULUgwDPJRYA0
ZWSmkT+dD90GOOpnN5pYbKSUuISh3gsNyzbDlxP+x90FBXLS8jsPAeKXM9FuyTP+lS+tEiWaFyw7
/LNyJ/eA9KQJ5IapB3QC5uuxM52cfbJTbQ+4nEhX8xKpcOqWVcHh0e4q2LTzm163ueKE2xnNudmC
dRmVbcQ7NMEKFVr8kDwpAIfyVfez2WbrWubPpxlF9nowXYtj5rJ2paZB813NvkZPLFJC1t0dJazV
ycxjq60Sec8LDbjPfjKHhr3Ytt4dwAjWjabwCk36qEi/ZPGimN8TFVAy6LywtDYduq6QY36O1Xm/
wmWo7i68oRqF+2IJ/ZUSGUK0kUHFg3uq4ISmTRFBKNOeFvR937c/5sadMmLMTnpuTRR0jpeclx71
kS6KDWlQq2Nt/FkzHpw0qMkZQfXYshgZXcvJ5Ywh465Jd9EbVqWy7OfcgpdtNvtk8NOGOzR+2h7m
LpmkN/47gpn/4lhJq7jbv3WZAH80NVKOnxVd6zp0hZtfYnqeLeFX67LC4hLRECEQ/IDhIBAWsZZ6
fTFRpV0buL50s/1v8jw6raiWskyQ6izthCjAiUybO9/WGkXSdLYFBfRofYRSgJHKL7qAgtaKRydB
c7Osqkp8u0TPSF673H0mq0RvPdebeByJjLjpSj5EPUi2C/ByK5VHyOGoQD+Hx8BJY7qJjvnjQ4N4
VlumwNXvBdSfh7/RSSm+rWJ11snTWspfC3omaKS/4plYYsV7odJNcR/30sAPb0wVLncoh2Tby0AQ
yfTti1tSqgr61Xk0l+wBsEwW0JdZTZp4D/yrQbHj+XGiiaajVVH/M4m0yCYrCMXc5n9tRU2m5EHb
9lh2OfIDFPetESERqOgjjPDt36ce7DiZfWrPZLzbYCBhWILXNooJew0yqkSTtsZPJGVMzYZew6+/
YnOBsEB/4C5suUrK4QC9oosMnIYY/WriRJfnET2PU00XfN7PRRvCm8BzA+7dC/RplTyjTcTlkUdV
hlGRn9dRJnAg1D52/CwGTQX9tSG2n/fVuTZ5vtusgiWzJW1Ob9ws/CNONvd6zb48x9p5Y3dZQ1Ji
7hKpUAnEG/74CpJMTLkAK6QVWmMDERdlyxXQUbaTlR5fy0zQIqcjn825UvriZ9duxXgUtaY130MM
2gqUVqRz45J1kD/e1lOxxFd5ZZaupaHhaAkKLPCuC2FaUDEtMkQAftzRl/zjSSHDVP1eWb+dJgQu
3QdEpt11m3294u3iKhJ7a5XCVC+XtBfYAPbKwBWzdV4F37AG1jd8hF/WpbecyS+a3dfxnRrotV9d
Lf7C98pPwTcluLn+MZqJYkpOfzjB85bc9LH5QZjCzx4UFe1cKOn1O88sdv8RLjuA60bC1eNaoEqm
K3KmAdsNTUHTkUqHa3Qdv/uh95pFgVj6Y0yxGw6NRlQPK86b+AjMkVF3F/U8ij96pxApWGCN48cm
RoV9oaTr61TD5hHaKaR8e/XQjI6PRksS+RvnuQ9yN3x9T0UWMz5EcrK/C3pIeZ/1bDJjc3dQZCEA
C5Phbj1Yu9HZ8H8vSnFddM6wUzvSB/ptnpzw5zIDe35Zo9cV3sgUomrg8VrKGw7KC70PWY5Zukwj
ZinVnhGfXV/0Vffg6XjS0YISY1tvWvskMvNRi/dCeZx31acHUbSIvUai86e1WujfPR/fiEFS9aa2
VPSaDNGShcylA4x0bH3/dutp7Nv7nG9DGHNVuTusj+2FOde8AMy5Q9oJYNDuMucdSGTo7Q64XiiH
Sy2vScySibK+SEvyLWvJF1ini1aBWyzqDl4aVJOa+gjfDrzDCwtyEt0oY6DjrJCtDND54Dwqnh3P
N3/b+K/Wu9mqZFiB+k7u6jzcB+aRcQAEHvxRP40ydvTffaes1oyfpw4UDC5MLhEn5gkZUGgzWZyp
aRI2QJWd1pXlE5yxV7T86CasJbsZ0YGhBUKZSEv2KOQ+SPwnRa5FMFhv76Se9tlUFqxjQ646auT+
uLyIGNALiu8G6QHKLVigRoAJiRtq9HVR7Hbwt7NJz9tZKapj5yaNkEo/Z9Pb7HHa9knYKxuhm2lG
skB+vz3wlpzuyCSSVLXEyHmWD4LVttPekC0Uin/Aj0vK/l2uXLW2l51TzrXhtSpuMyY7FeIH1aqG
6tJwNXmRgN5vmjXSP3cTmJTXzuLeMEyO/4CP1z0LODhKfPHquaOK14CuMshkYCyKnXXTtV7d3M1w
rl27kCTn17Hq4owVl8rvcLtG9br2+VByMa65WUDfICuTJOOVShuzOLrfsoJwly0iXndVfmZFLzUC
EenzQdBH4YJyYZb5E8zCUzFH22mzqn11btWX4rFWJzO64KRuMPkz1qWuOiTipJ6NLRJRhDrIr3VR
RCLju4Bn1TYw8VvEVDj341GKwy6QRSrHDdnW3r5a0oHrUSmmHKRh4/KRZV1pLT7u56czPEQuQAIy
ZSlvaUR8TIt3jIKvdR9/QUloTzg92IKOV2YYqHhRno90q4uAp1gt5NF4EMORozxCgV25Xk/p/CNP
zFH8XF7NehPKatOjxmrbiAp1Qzn2POySFcYx2KrNpj42FSzSQ0JzvHbfAQfrGE95uMYHTUiSHp4R
FSYx1mFEvulCDzRRmv7KuEU1l+xdyghrS/JeWyTKaF4gJrC4XlZRXiBAoXKEGBKjACy1aIu826RV
y0edhk6FkbQPsWKbadzwTGVxVYgVP2hAhoOis4TsNsJ63I23cgI5iHcDhrI0DCrwBt7bDQFQskpd
AyPfsm/Tq0/K4jkY9n+W7Nc5wcWCv2gu99ltwuUWCjJnj2FJE+weOsWrJ5tcylBhRvOWgbxdNU1/
4ZpYGTbH6VlGDMcxGNDzDI0YT4pjf+QFC4EmEj6ICOsBLNgj0+CKIPfQX73J2HE8TeyjyKnzo3Ef
342krVt3/p7XlgCgchyL1elHNBhNcfjHo7Nj/eSlqEQ19LOgm31XJl5qHpwQbAWjZiDQtXVaKLwE
3o8Dh++VrHpwW6aM7dbnKktE6UbKGp/yqf78Oe3NzcouusyrYOd+QDfNTxZeN4Hrr2ApaDD2CyDV
S4Tb2fvF/FuW36GI+jKUxPbv2nZoT/lrE+53QKonnZX04TQn8MpRGPGQOgXtPh3cw5wD7lJbu+CZ
PyaUcoObp0Ps5KkGWVxonNHHuJg6aoH4Yv0LndT06uq9I7lfbek035EK9cXsVlFladEF64yyUyGT
O3hXvdSDuapWXuUnSjxG5R5uQo78Ag5oaWJDuiu6dz5YMx+CZWPL2zf0jt6NptMjjeqKk3x/pYXN
seZ1gTd6ToQoVrd7eFXwYw+6dh9B56p6JGlAO5cLWms5PrM6QM80BvePHAZE64IEweCFTizEJKt4
FgG89YKNWKWzqppKii/czfRqmw9caBJKyHnIb2DW140hzDII2r0mTjjPLvaQeot9fPZnN8zwbKKD
Q2yjPcGc82K6P9cMTrjSEk0Muv9MNQhF8nymwRgTYbcWms2ed0zIjoznf7Faggjz3m6FUVRVOrLV
OCSMORYNpJZ36iwT7I9KBhn3smacoAPg1uzWH4NJLs+6tjhQFqZSxwA47n4jBXugJMO3aHu1Yusp
PJSrNDqstF3XqAU3E39Aw7h3vOUGe6vPga/zVndff0qlGaaMwK8+itbegZS4VBRIOt6+b0fUglmc
S5yraSquv1fndCh8Ii5ruG0gAIsxSVOfyHg1VLsBhrZKPzPksMhYVj1/dMn0CLtk0PUM2x23IxQh
Y9uipapu4X0OZglzt7ACY9BZKUVtxmUtukB4iynnBjKiBH66iIYbvPmV7m42hG4XjtP09BBugTxo
oMLt1/m1bv9RmqUchM1koxJWNW9jQeNcre6Z6IZdDm4qvDGK33ZXtWhqoks8dhHuTk7Z5nbI4qPy
S+xTICAO/+aONI79EZ0Nm3u5C43QjuwF/HZzP3AjFtly3m4p2kKQW5IZNnmGW6wGR851bhtw+Ipj
AhCvKJ6L767ooEp9wy83AKIWe6ZLWMN+ypCczC1w5MG0kO6tiFwqUwWm2/9lSdw27vHt8AqftVtZ
F+f7jS9ViQA7L98r2eoxP7c4U0nBBmPMRF2mAi9QkprfI5EsB7fyMcjTBPx+rz2dtoqj9RsrVz/W
CK4NoRE3427usPAP64TGNbz5p/dit4IlhJ0By8go2Fa5WhY9mRV2N5W7cfS71t+DGm4M0+dGF8m6
PZJ+E+dUsb2Uh43TprUb7RlD7MxpHvCuWu8XReHmnbneeXsfslEHYP4KUaUcNUOlkyLUPF6U4uVZ
wVRKnSGPCQ3tKdpeUvngTcsxHMpL7DCGY+dk/6kkxawd6uj37tnKQXacsDJn44JsKkbzEaIfJb4Y
s6BGSNG84JNii6vJegD6G3lvIsgUz8V7FR0nBM20Aex1akcsBkUHDKudtn0wyo64rLF7fTt4WKVB
jzJjXlFYUZKE+VXmsa9BknGxJBd9b5LiG1N2zUBVtz7s/bXkzOaRidJ4xhF8z+9PhSy/5pHt//YJ
NlBlyPUyCTn9f0xKYR0pzO/I5sByYJ6KBhwsMw0QwHUq191z0IKA7WXbBmrXo4cNfWZRIk/P3B9h
ceXdnED1KjPJRBrH79560LGZVWN6kEUviIe8Ekldjbe64SNIJ440WncNesALlqAlgx96xnBXKR3v
tlkYGROs/8dHILbcWF6o5kYmKMB2KqsQmb1YY2UMRkIY6HT9g4JuEXOWf5GIvcS5IvOVFgbE5WEI
GDxl6QKQ1VTXwUniejBOKYw6AWtn2Wzjmbfx3V6GHyArbJg99gwOPviBiS4Utd3pz+ZllQKiMd8P
yW5sGa8HeXsoYBBMdn9E0gABhzUUOePesmRBzz7cvEJ+GeU2W397KRxNBvk2C3Q18VQKYutQ3Bm0
YdD6y4Tk0eVVOUCKS7jsfT4A0RRQa3qGPlg1Vez4Nzp9/tZJMm/3d2tMyAkyoo9F3cRi9sTRt3FS
MyJdANd3a9Ksk3NnOipeHyNH+Hfr1y6/5jAXWu1j58Gu6RG6WMsE0HILKQ8nw0X1vTaFcUvd+qd0
dzAzUDZUnVYEaJDiiItIWyxGobiHt90q+7PV8LIOEVJHqmA943Pid4n0FAQlVKZdAvav4/St/dgD
l+QBw8gCjGOviV9FrjDkHXVlI3DxWQ5RPilTeg4QOv9jNCZi2L6Z3Wzee0VFsTM90IgYmYtyHp0B
QBp531aCCqX2TxuJjcQU9joP/iAUlU8bvre9JpkyZDNKzGUtwexKbsmNWLirgh0V4C22DiN4BfFx
fe034YJuT6TWvsdK3pEmSYPzXNSXwrFgeL5AL2ak/q+WY4vgnyANPHk26hgyMeL2V94DGxsJ1uD+
7rff3EfPnlgu8KurfzYwBPz4fIRUuTKkw+MxOkL6IylS7H+tM7y7e860o3cXi5qEbZX3hGGNqUS7
e+DQvbS61ejtybGbkyY9Lr2JL4jwONI+7KDbcUt0JXpHs7RFaKqyDVJQ0RJ6SwwR0JF+4Z9q8ti3
kyFcjJOsvLFb0vSp/jG40lVqBlZZpVp8dR2fYbD/OSq08uoG5EtsQWF2swWuwMGsMfSWXCTq1WvK
1wwqKNtNDJEhFEl6/tasT6jNhNRG9WrcLf5tlfdnqClJ2iQSVaZelF/xPXclY04GIkBhZmWcTrQy
4QWV4a8Gjgq1aDMI24M2Nh/B0M4yy6wmqacy4ezjufclMY9jXLLaEyduAXjxRAlZlBEtNOSbzHxV
diHqtwJ2ZSFnH02mpiRHN5RQfDpiFM6x/T22eAMjLs9bMYjLCNY6R1Kl5F5ZFHFFg8cfYkm4RdwL
HwtmYXCy4bQJzAHJstjidGhOV3Bu+B6OtaReLO5jNviUIYW15r4SfPd9lI8icOrxuQRm/fSsYkaL
Xmgv6h1++Cqh5AUrBrf7AbTET8gr5LmLUsseHf7KhEPHAo60zKKg09Prd3MtKVUOW12FsNgBlDJl
tN3IGNZJ9PJ7NWUaCNbD7MYby1Yuu3io8EvdCBnwhWdhQt5Eur11FlKlsYjU+DPBqQNquyVQaLU+
Ugqj8++We0vn4Uzt2yhM2I+zovGxNb1B+r3JwNEyTnThlm/bs07zngdbI+bdnjItrAmRDr0ttWmF
vserDq2QK8CG2Z8IZdRz8qXlrgjC9Vv0R8Z9Y2Cv9p7MxPO0CRcfEyDxF2ZTwtTJ+D3ZHM5LBJvZ
bSxEgOc6dujckSoopV0HM9ixEzakbVSbK0j4tg7Cjw0A5S6agO3UjhlMmMwJSlRm/8MllaSBDNok
K9YEp5k61lUFKgw7xAcI59b9CKO+Vr90kuqPkF2CGAs4pvXcK5XGpGHWGldytUy1VDovLNJCzg7a
c1GtmzY3QOCOUoyVDlrf+7o6HSsCkPpdzR389Y8TBNnKbq3b4NYxe0l5GZcE9hly5VkM3zSFHf/y
KB4SF0s+vIsUr4YYq8a7dNo8r7Ev4KvvEgLUe8UG19pvlOrc4iQA5M6zS7we6RIjMbsRjl/h2Jsj
ZNqzq0UWV+PdyKxN1cBtBcXRvYlpb+p/9YrY8Wjzsdh5uMB0blhh8VK00Osbm86YuWrxOxVR8xkm
Ewc49fpv0UkNA6D9b37SDYEvsxd+vrtTk81YFlgka4sLjzx0zxuIXL7lj8HUQ4aBypz+2W6NXfqK
QvA041oxtdekj3M8nL6Z549DyQ48F0qjeA6yxFXnu7P06wYXRFqz3AayoPLt+6H67qbyUoXhqe4n
Wr/y1nOu1HJLas4mPI8/O7ONcpaEgjdhSmJwRE8bXAfS2Pqvs6ye3UWZUkym5+8cY2aHdgskgFRt
2aWFSGf8N3kKKu68R2FFEu4q9w9XnPG5QCA5PTkkNv7lbZQiSQxQD2ySfpj82hoG4z35kWJ1wvGm
Y9mkKavUHK4VYO5Is4zrckn7X0tyK8CXJz4bYvA+V6bAYG+k5LtZX1XYy4Qed4uztlMn0fYmfbsM
1DDxmwclLNlBcYGtmcCYatTLpK9eDwl0hqLZAt1Hmg646aAQ0vAPe6S35KJa/FFGm3yGK2exj68s
prxVabGxLWQ/rreCH/5XgnLkKAdk33EFj/7n2t/TvffIWr7pAbFDgQckvfhY13VA9Rpa8V7rZAix
zhyI9VATsRL2DPeRJ9BNDQ3GLRhNQ81ruE1OCJH1AmkqW3vPFUpcav0BHdjJ+t+0D5UojRD4Me5D
ntZlvAVoRTrTqdpNcMqbOa+/V11WQfY/hhH5sGJPZGQlLkLD8UcMRYp6aT/22LiNJ+jqZ8qPbito
vD7Qj1yjZTh20TgBSAJJAVLWu9uFMWBikLEr20beesZjMCHsYCb0ZJWXfljhOFQ5EOyHN5vLEwwu
p2zcL2OXM7Jr9bgRVcei00DV7dnUgjqr5gJqdGaYnaLZ13OAuFgrytXOYhTmu82+ReaWBPaC2SgL
TPxfhKSTw6MHZ/R/dgAQa2FwXya3WOUU1jgHY8CXHHEf26Sb/6hHs2EEblyuD1l+WeCWLUeRG6tf
sroHUezxzNkWSyCUjeC72tI1t0sBZnEk5RMsB326O0jeo148mLNR+q0ckWgyrVN+OATiugw9zyAX
evAiD8KVA1ApB1IZttM8tgOLhgY/kmI7oGdHzYGCTjoG9Hyopw8D9HN4hieKuobNnnqCNxXzZ9pb
8dudlIMgc+dfl0X2QicYDV8NOJ7jAehOl9IjEMzVurLpqxCLyc7tuxQzxPtZqt5dSJ3KEcBl5mtT
xfB372HSiSlyp+UkpfE1tfjnlENBLeJ2t6vvg2lccFST7ONl/evkINI/RvfLBFn9vsc/CtVUJnHq
70F2yjvAH8+cBG5h5+hO2DxdqAd/RtRdT9+87bII7dA3S5DnVkuLdFVGlgkkKczLhaF04BshZDjw
0Z4NehQZFBG67z1GgZHqLaJTkuLM61TY7Q55Bj3TxvNse9VMVYtdOeW6EK45qI+ek/OXnKILZwwZ
avYBwGBJvMu+rSqJTzg86HO6CoTKS+PbpQNtC8FTiilb8uPe4HY0zcg99hOMIIJhtV+TsH517c8z
6+tP4JM/mV4cPRCoQdrFFFoIFzhLjjE8q8nND7Yi46OiXJq/T6k49JFqv3BJK7UukAWS2Fzn8HCa
/3V9LT6xq2ldZUuu4G4GtclSFWEjIGZPzp1+iGgLtX75oQJ1Pp6DC1NcniHg8GnzrRzHLR/xXVmI
zxfKRCe0zIjrISlya21mGA3fAKpm8h3iVHuPPT4qKRYQCyXH1m9OVHKfjgdPVmGu6AnkdLN/dvJ7
GEi1bASM6+GB5YqXagPLSeIt58gc9jr1QHNHprI8tePstYrrxcpRlDgH47y2e3YeVNL7ADrts9PH
wuCH18KlyRjya2dxo7eS2KAbdM5tpifOLOhLWDa9ND2++flbXQr+Xk0KjZ/z56iyPnQcNvfdiGlQ
Ipmf3eno23ZzwlFw1a69gXxeHPio7hrpvv1QxZieW7EBN93Kco53d36KNWvYcjmsLpeJVvEZ47QI
L5LEfmzCDeh0PTck6YVomCnXZPSyE9VHVf90E5KCa1Blelrc3wDHMGoDazhhEGBGgXhGRNjtgoCU
lwHEdf3pqEzlMSabVOW1E64C4hO0H8vFp/1F7gahXQNl8L+A6Twc2MLFwNUwKjq5rmkZZOCQkkEi
f6fOcEzljaPo5UMuXUJdswnGE7am2sSatU7LfkNnNH0IkjBz/+2c+dpw1RXvUuIvCKGsCykLes+G
pa/4thyMKxQxB649C1ozL/xAa3NBngDbVBDVu+5SChikucRV6Qiy0oRdJ8HatDN9KZGmclDdzBBb
Fd6Z4Foh9WnCO2IYcNFE87uX8JOqveyV2Y0wJ+LruyF6hNtNp/QNZPKh5nnXSHRcdpLet+yceTk3
/n+lxp619wSVSHsy7zUez2wyUEq4FXRr3b3HUpVnQVGM9rHMR2INIy0rQWFC3ebVKSs2jkdw6u0t
tlFEtmA8JXZskxrmrh0dpTapTvqyaLBNdJ+RC7+407mUwh9H6uyS7EVwgL0RbmVTyxRZY5Yt6ZFy
9vdU82n+5WtVO5Z/KpvDTiASzjWBF677GCk9aiaw0LmA3pkDOdvQKIh4ujtt+83Uf6ZXIgBrWYVk
M4U7qM16vcKqquWTSNUuY8mLP7OP7mSOmvQWBSeJ0CyqN+9UTLXjp6UGAk98rHCLZXGUQFr+xaLu
HtosWVqlEs7+LY4AqNY5gt5Z0v3xLlBcO5IkPMoFrYlxVCIhqwktKfok2XqdbSvnxvgI90VZDH4L
jiNxurlmQrLjIKlHu32fH89S+aXwGqNgTfXoNuNaWh3LKy+ARPfXtF6ZK1P0/NmGYacZl9asa7DV
eOU5S/CU3ANw/w0DNo2rRE2q8YYqttRmlihQMW+wTBtCMmk98DpDZJ1JGlZVPbBUxVyKDt/BCJ7G
87gYpVhc5IwKM8IXn6xJRUO/mkAKEu8Z7p/PGfIgsCcjX0JCR6x5pX/JSh/b8osBo+Auljpo0vju
j/IxK+iRFjD9mdz4NDalE5/XKPzgxZHh4rWBUOTd/eRXOmrp67JGsNiL+Xg55VbG2KS6KyUd+7rU
WlUKWVWF49/wjzJuo09/lF8XS4Op3LWDCwRn5kdZKfo0H4Rh2ivq6LEI229/ZpRiUydGQO97FW2n
pKauugyp/vG8819n9JlZTAQ+jwoHSKfcdGv0tYMICfySA3tbGHR48BuEH+5nGR1EEx+S17hL87TO
xots5ECGT9rLaqxtu1XSqIjZJlP/jFzsSA+kK3p+OO0MHHG2stI4XLHD1QK7mtWECRcbA+hZEtQS
YIc8hrylE8NLr2Zgn47AcjQUFXnE8LpL0lyGo+O6gJVD874ZDJfNbbYruPW+JlVFDGED0HT+cGxE
a89knEPRJr+yTQKqiqJ85DeLSB0OgARzn2GBv3bKoKbf38bBa8oS1jjdbtrIFp/QtmYbg31pjkcB
KtIVWfhd5Zf7EdwCfD1KzOyeMtCvkszAk4ToipAqdI7SLpOPJYV7vMDzsFePRjSlgzAPjY3LZ28J
/zxNEI3O9Yvq+Q+GUM07Pw2V5ywzeWsaVKWrC9mpHiPEXbSF4dgP+k4FSnIN1g44OOJKoNdurWdG
+ZjJO/lKmJGoFn3edgSqhV6zYYUbs51cJf1fWa0bxzqT5p/F2vwhMpff5kkjUxI7ptpYLuy5s+o/
QqspAFzNcnSgjqmeEv/IZpIGFRgN54dxLVvOzh7qqbYd8eUY4Y/Mg1sUw8wd9cR8oZioEmixQxzZ
R23oix7qJPaHv05RUO0I9AoZiHXPJ5DXiZJnnnjT++I7rZbhFamLNEbeJRagzuk9kCwfEheh+sKL
CQBprUJHMtGs33NAcBMgBVFKIkbYqLwrArK1nBkNR42k2PKAZX03CcHYfhDJKngUtqISoJBHjS2m
NlBeSOMfNeh3zTfJbppQ/Xn2enJMMo6+EtILyL2tBCN/tNi1J2ADq/x5npTVI1EpqMKCcrLFz77F
DQfLRiCYbhpMQp0mDKaTRRPYV6ieTlbB5BYMuGMyhHDBGzljlHt36pYNrkSv2REX0TSO25OaJKJB
3ISr9NHm5q2GAm9akDx+lCWLR1EgLOXl/ZgjbTO64ndvoQlAUutmBQSheI9bNKBJOsFM86HH8fsW
kmOzmwq/gmR8XdlV10SWvc5H3dUfDIXha7satCXDniGbn+8ywlhtG4OhPVx1fK+K1h5TtZkH1vIY
uWMQn/FVynF3xmHNeIm8Ewh+/ASReDdc4YP46oPHEgEFDaWruKccD+rtEuSesjuZqqQF9CYUCwRE
lQ/BPg0FOD+j5woMWrcuM7OFYFw2FGZiAn9QmJIMvweFcRTpqhZtmH1MfkyA2ez055PGr04g+bjy
UaXQA4rWlHn1xmEh2+a8+/exq/CaSwVBI8NgZaA6yho23GP5JIKFCrXsekzrqlMyG4H4AJfs6bcK
XleESjimG3iSVloTGHYuhnM+dn/51OFZK2ik9QlkO2lJQR5FWZv0rtaJwaZWc37JKZSVvNNQFR07
kDhQBoqqehtlGOuGpolNWUzWbU7yNFj/4tQVvytKG+UPFHY0yT1j37zOi3cLnzLcArkw2vGNQGwT
C/3c7PJrPQgEPkYVvNj/+f+yAjkI8+rGnLbocEjMCHexTOpe4I20htmgUmzQGZO07mRnTD61v3W4
0bhYYtstwFEVLWymoFiVMcJ8x9/Veuew9+eGP3bQwiFcjSOhiSu/v1tkDv23llITzBi1U3R/56Bt
b2/haInj5J3d2WmMLofWM9kTQulRaXngjBLRvlmS0P9DVhjokt6zU4XgUaooKdCNlvlrhPY1RkDE
rNTiDcpITmKV0XFg0a6eUACTxgDynaicxno6aiCzbvhiWfLdnlCT+HGvGKSeWVaW000zk1Kle7e1
B0f1ScTfraoOtShMaXTJIJmR3o/IURhd8qsel6zGcgSv6+T513ZnIrv4GCqsBWwNzlldwznuPLFy
7giLtDM9k3bOBjEliRr0/HSjjUQEmJeAoj3Pi3E8dX2EybOy6aFMXB88jdlC/b0m7ek6XEJJMW8f
KrlOIoKic79j6IQxDuYOrSnpMr6TPYZLkq6VAs0cDQvbTKrK5jmv0SZA0sGF8eRh3AFJHDJCVGa1
XigddpuS+5Y0uhxWJnAXteeoIuF0W1Tps3KmtLgG69hEqvwzNQWNHlxsXDX6Z2R+EW8TeTaMpnHw
O6HjMSiJ7gBRt+OkoJrNyNKDR6zNJfen4G8nSRjUxNlYixqUwu/lOpJfobPk8KhWVXaBmdHSZDbX
1gusVDS5vRpVrq0U2ayyNE6Bao+Eg7UpiIJpfAMMvwEIhgTtCSkwUueGmSrpYRvfSniY8FuLCn8w
GQWpPunCHVyxlKfIMlwVhLMbemYxmfUQIretf/jk90eJLayPHt7pEiUxpLd4I3Jrau5WYoFCshg2
HH28C3j3B0GIkS7oubhyAeq2FxYsmc6SjvmGtjBeXuqrrA7Gw6A+57u7v96hbsjfYclbyLuTB0xi
F+mWJ3IWpVcDDEcXwKboTPsl7t02AQodIwXoR2HETp2egTAFSqdhyFeILJ+VQNUC47iyspcLffTL
s5Ow26A3I81lEoTRUoBWFFvg3Z1f+cXJbGKKmFzBVm3D6ENCxrK7cMsBjBGUFF++mKcXR30mMWMw
FLOXT0fJ21golbcZ5fS0XfxLxxWaXbQ69BwHNAy4VgFAGVweX4oMaoL/UnE7GGeWH0G4iquJ8C9i
VuKaOBM4f2K7PaqDuXQBLRLiFn8vFmj4RYjGqRLLypa1tuEAL7HFR2Y2OjoEuYR0TIL2Bo7VphCZ
g2bQHVyD6FGLmbqp+wSnSt2Cqy2zZaZRWKuCPNfZgIRy0+EecHbCQACfu2DMcr+GXy3mItuXz1eS
Ti5Rz48H77Mxcx7NjSINHt4ft15RFpKcZGpmINjdZY0U5N6XD+KZZ+UQ/GvgfeSoydWp7DZK1zOo
SjIxDLY4ARFhd4WBI3Jz3eH1JWaSIjME318AkJQtCYIWORWZgUvI+7YTs5Qy7nVeD8HeK8A+dYes
DWqaHyFWnD6SQgFh9j34txvMKOmt05s5HtQuhlw2tC6GXJfZa2IXbENQvsfyeFeXIn7ngdiKhGOF
Yx0+HvN/1nc76RS3LkdaxzJMRYYVewixbQMJpcw2MX9AVwS1SjpMcEV2W1latYUkFjE34bAY/9Vo
Z4Mg/Kl9CHmrCNQG0oV+Ik/TxdMgGirUxkBrUr49qnY3RWr07UkIbsNxKzt5ND8TbwIWqbaVWG1h
KGTiZBR0km8MCdq4SisTXIaSyKd68YPsyhKfMO3W8QlFYaPVKuDbMk0+O6Oz5gnmgz7L96YC8YeP
uqqOnFvFUafDKoFpTXK8ZqNe7ZsRVOBZpYaVbjDFLwUlwyB9MIsaidhPjwq/Eg6NLMKtnk4nJ3ah
0Ry4oaXr+UXX2SW7++49owOpgFQI/OCvh5qAfsyWWyLR6FAYJIv1cYWPY4IRl7ykjwyG3YxASIdf
ICREhMha3ZbacK31tHXvnW5QI9EJQQCXAC5DLoi9IYq2PMGDx5owrEVLXgUA+5tUcj1dFVIA94B8
uwWUi+TBLHUXLJ7yGDAnKBOUW+WtEguHbyRR2GajGM2GRTkFIXqJ0AP/pclXhS9hDfl0hjRStZQ8
I31HO5fjHl/oDgbl2Jk1d5YWvWMoWEbFx2mtPXqI4JmXDVHCLcCXTQANRVaMq+FJuSzgUYgHnZa/
TTRxVhDx3OJhub1xJpPBmGRr33NE/LfSfKQcM6ZXxF8ffnnBr/FLKdrGQyW7lS+PMXy/XKNMYdAc
sEsvcsTfPrHuwXDTDNi0oHY5rvzUfSIUiBWyiHbzBU/9ABt51+OkQb5X8uIVhqhaCsTCgOk9ZoLq
q8hH2S/5jnKCDyk+wU7z2xhQJkspx8HXWT2/+SDJIVHE1LD/CbgBsV7/06RTglkdw0V2faMfCTnv
xlnak+d618VYnwW+Mh87r7NQLA7ErcyPfFLugCL4tpKYmomybNt3Ps7iQrBRrXKVOMs6UZpD3EiW
h6RSUzH39dYioQkmBpYHdaLx51OGvr7XLJOduN02q9NKym9jkYpZ+Xw7kJxv5xpduQbZUE9Tutun
JW4AN5EutLIeKtC3y/78AcY38dxKHxBjXRGc+QwB+r8bObv5OhyTxPM3wVIFdVEXn7KdqX9a9oe4
l/Xka6J3DDJ3ip3/ZIW2MxGtwawPdktN5FuUekIJnmfseYOQupzVMxgeo82X0PpzxB/EodLTi3ll
qhFi/hjJJYayNErLhUzcZOP6BxuTpNr9ewNFiHip5wh0OXRKLRt8jrPjReGE0t9PbmpcppXUgog4
PaA5WXXS2xLupYFNIVySBHAaoM1F8lIB7Q6gSuqBdRHuu8fLQmsx8j6BcbD0WFwYraR6oCeMuVjb
yhOpIkSycpcUhvyBjBWwi7Un8u6N7d5u494iyMA6oj4qlTEwNsAfsaUgLlQsPPoE9XpCufUEFcpa
Tr6uTM7Yz+ebpBi1H+YtyzzQkHi18aH/d13MdDsHCN71drXo6PdjfX8MaqpC0h/SBYMCHDxMDPC0
84cAsCT0nQYyMepo+nBBF1fYb8ttKPDSG/4kemoPNoL9d0uE2wZ/bc3Oa9eJCaLT+ndKY7nK3el9
AHzqFsOObD8LD/mf47X//Xy1zDWMfj4omR4xWbcWCHqtuPw0M2+/HSk8hMBRwkapdu5gDkTfd3MR
nAYgUEugtvSFhv5Eb5dFhg+E5YkmvFg1HEKalPpe/P93wl5o059fKeG7elBiqQitpJR3eatQWzkE
bRtPP/veJ+2F13FpHgD5ZDalYi342GuiaCnS/5etp7aP0Cx8fsMGp8NM2DcnbiUyEZsDpSimELy/
SYxTZLZmYmQK8aLCMscYudxXMoKwex0iHIyc+DecFrDuwH0FVvdoXvtu8LQdlZcZbdCJ5pIkdwN+
+GwzFj8sx/UGirViajVQqqp0mrxHvlXo6srxnNdzeehiWGwwRZKZCJVC5BvQ1Qsv4zz9LbjT3Syg
T1S+gl1aH+QR1AAGWeq4JfZKFrwFaCMjp4zN4cal6Kng5zmQ/e1BMzsxtMAo5obKnMniZ/XGJMxF
631NZieVo5uCT6qtKzbkQkbd0srm4ftrA4k97xv4MjZlhvaekAq2Gj40CBonPYWXzOqMIpohbdKx
irh1fZnBDTKN0IQGJbdLKQL4kmS1pEBm5ZKopOIrP/ax33JOO8GIYgEi5RxtbmJTdaZb6s3reenS
tmrHlQiElAFuhf2J5k6L1b/ebMwjksldiTtxHoSQaknXy7xQTGvcDmfIGzx6vD7VOHWs8LgdEyCS
OmZ/OcoPF1rLEIGZgrR+d7/YFDC2KtjbjbmqJEKy2+pXY3g54gFKIpGaYsQrnzmiRNFebMiA/iO0
cTMrnoa91H3aoYClhKddpNov8DlbkKK5BwHXIlmP6ZRr0Fc+PHjNuXziUNqvIwg23X7FiCDPe73a
QGXneopBwAf95+NvwU40YAndT+h90mSuGKfUdJVeZLe9ru3Xs+cRWEBSTdVTDhXpQkMnlaAoKuxk
cG0RtPUWG6j4OZskcEVfuxo+zMSSJQwFXE4mC068qC+jTBbNSuzf2YYQFYKhvXQwYmHwsG6Zd1eO
yfeQWjtyQP2SeTK/bQjNo+v5TpynIq1SK51MDmfCn33lNQhKRq1IG/WVKxG/GUAqG065yqdCsvmV
oRZJP1HeRFDloQ7cg/SEcMCb++XfJd3WMdj3uBcFRcn6f0dh8v0BqDi7lLP215UvwlxxB4aZHgDm
k9vlx7NP7onzFJZ3/CRB75AvshQoIc6moIUtnja1ezgCASwdKN2Pq1+bfinzQ6zVA9oDl1HBUjwm
wG2r+tVYjIjFr2CViWzz+ZGAJ93D/LPC/j/f3JmuMShq3VdavhDWEjCtT4bpcAcO1PfAfrL+tTkF
1GfoRAhDRLYU8DgUWdlGwTq4h6UbhMt4nSfdpuL1K/xWWt3e81Y5KGjDv+q6PhC0ASs6Wn4nVSh7
DKdIr9i6KeFD8fNbvrJtujw16OU2SRUCYbmtGOz3cyMHOJ+31dTwtySJc106yhIkAbDA/d4tSOTg
O/SPRl06loKTZU8xxpORVTpx9re8e/bygA+1CSGisy/2/GKVh53Z3jP/QB4l5LredxFEFXwUYiIJ
15yi7GBrLzUvsz1r9MhIYk3LY8PG0BmR6OIcQvXLvhmZ5dMeXQR7KHmTEdhpC9HJcjt/Un1NHQcH
1FQsvCfIy0KTzfvh0KPcQ/0nONR21khdPibhqRlb0vuKCWdwHcPwRcvPmlXXNlTfIzv+c91BGt3X
n16UupLBlxlWaUxKrtE7UkOA8JHI9b0pymqPUpYPe9hx7IzmDp1y3oWJ/l5VfhjW65de10ok0Evj
bvIzQH4BxT7kE4OHwFFUYDvD4xFGaGvQeLgjmwnfE/4n9VRehuhuVSFH7TAfKO6IHVpAPBcCoKHt
RcGuqskD3NA0WkNeF1pAVxxosyGoSp0V5YAzcij7spla9pKueB/xSxrE8uT1UXCKNGbyXoqKUBZK
vjj8AdbL2K91geuGKJyjySoWKq02o4RVrQsbIt6SUyx51qRZCP1Lq6IKXI3cNk49uY1CIjhBXfKy
dw013ktAiqDvhG0A6NCTVqlC99NLHSEG68XDk+4J2kNdLLrBY3uTBvEfdR3hokIx6NtvMvzicWtP
7Kbukp1bxTHlwlIXMGk1Qsj3yIi3froRlydz4aHCMrLXV5pNOM5Xa2V1Ge/3T0JnW60oJl2JOQQR
BW0R4lm+VbWMHa3oDT34ulBNeCoRKGw4FsM1BaFKQDxFpmKa+WmgL0XRs5muoQAvpaejtTwbN/3X
3x+N+F2LkTfDBQ4pdKVfw/PwRrJfvtJUxxW0fZr+3f58WMk1TiItb6Bx6qeb90Gcec7iwq97c+AN
woECIL3dvQeONkAJ2RA6+kV3rIWOrki64quI+2EYW8+gHNWUj8LKmAJ+1xGbGTmqbuxwWzQ9bjS1
yE40DHQrqQGG8dt7cit6RPv5THrLW/qO6mTAE/LmTqrFjyj4UX3JUgPMnY02SVGit33j6QuJGr57
7LIGj8mQbJ8Sxc3WQFANSTKMaJfWGgOR9LyiRNBMPOAORs15kuNBIdpi2doxGsJCp2VvATvfhAeV
IHLJxdWPbvje9+yGu35rXaP8+W6qlVO1BMJuvx8vbN3N5E09EsRrUenXEDNxemH8PAM3k1QCo8Kw
CDZebUJH4y5695jxJUk7FlgW6mRDgMFWjEoYxas15Mt/ZtfpM/VgyTDvKBkhQxdHj8UNwwCrS7tx
xcskS4alDiR2P5+SNdPC5rGoqylTT5rqLiXv2SOm/0PTbBI7HyaguMpnRuQS5QUgUocb4BySNj3z
iv2j1y0jpNGsVtqzjUQO2NLJROyD8GhCyp2txoTEI7uVK6yB/bH2QYxLn8Q9j4DELqL1SaT+GTtF
l1Lzqp1JdrcUxwovi8y57f3BJplm+c3LjCq8HAZcj+zLu8lz6/G27etleFHXXdnYFI+XFu7RBmgd
mOsk14PsSjdoR5ay8d1UkOCCfTsQ1qR3c3k9jsueD7atvnkjEmrDg7FaAlDhyC7Wn+kQ6PPYx0xG
9RvWGgjL8LdYlA6Dd9pgo1KzCebl3rOSwHApfuVo1TOePetC1P8ITGNyhHvhQdUFeCyPOXgLH6Sb
EaDjL4fW7yt1ZlbMcJzHtfwZ4hxuKnkCoS3aMy1RPQAOuhX67eEt3M+v9n5iPVOHWcjwr+acXvCz
js3fpRzZYNEeUQvFImKD684/9hqYJc9vws8Jjz2wm/SsmyipRIBcoQuwGk0iXPof6mMs6ucdK7HK
/LLAxKalCrmT9NvXNmaP+Fi3aKfxBXmghU78GP24H85gzvbjPStav/kob80dQ0iIZS+iRmIl0pkp
9BJfU3ZMhvCHM78NLsHyppNGWF6ZFE+4MyhIyXLJKT2J1f8jguRtcyXw+g0a/EsS8JxEefWrSnjN
w7VKkcK7ReGbH5bW9zpTPzb3NTz2MGU7XH05WooMnjE/WE7bC9DdDlkr81ay1aju3sVRrvFM2vK+
JdgmxhB8v//RXZ+LwtWm572rjL0jpDikiFbcP+ZzUeXT2xD8HHoMd08NFpvW2e76kVWuRVgA/pA6
sXo6Gq68yEIYYpSUIdpwdVhD7j2moMFEf66bGaQYA82VmR96HR7khErIAuo2Lwq53ew109VNoy2/
jJaeTfxnAXFX4Yq4Edz2PPgJ0taOLFhyRj9QZlAm2rcVXOP1nahCKeHocj7d0QLVS/f79maUfrTB
zcBxqTUtA3uAeEAXiMLo3TnX1RkWlE1JDvVWur/OlpQsgNZ+V+eBQnVX/OrkWf4wROnKp5AL/VmG
cvGpzd5UrSGGwdfUH32TFMGV/eHS/l5J6YYktEBGqNFxSP//ITFM8tOFHuFW1MQYCVJitDDNwKDA
+CoCjPEZwBNrDzShzMT+ZPtWeMjIEz8y7MiaccvqA2R/bl56CUaQ1DRErwu8O7eYiaPuniUZ4Ubu
8uy9DH0h6ycT6dkMg0KWAPA4FIjefiQqJs3Cl0/nyG9UQLbJI1RMpunKEBow4T3EkJKn644K05Sv
abe4Yxdz5ultivHrtpY4yZxlU2xpqdLaPC19I36vP37jVZGPs88bAuhQaY9IoO4vXvFKozEoioao
KvKLjcCVWgo1tmvsh6KAwZDue/NJs9ICRbDKmph43TVfkl2orQaV4IGTnDOylh0+jIzyXafuO+hH
zdfRz2GPbR3b3aZjbv0YCVYhTxQawjMTPupUP9CuBeY3liq3/8nHiZVQuDnPzeoExArN9SnmwmMh
4IVg8qMJAaNYPM7XJ+4vG4FFmxpZ7XIVnTFF0a3KX3+ujusfbR+teBlawvb2xj5zzW8T1uijqJek
FHwRYQyaikazbECQ3VQ9abwXvXNcWlUeoqs9LKRl2y1pKk2EfxIEqoVp8O9SzmZp6M501gxkOnh4
Jtzd/NSrxjxnwgBvYo2aQPvEgUC17vX5duaaCU1nj+Bvtnz2jsh/HGMwTez1ut3UEHgXWisiZuTr
80qBh3RMc7fTF7mNCnViaysGm7kFCra3iF8IKj5580ypcvZjCda6IR9L6SrD4rxVO228aCLaTNsa
d7Q57GwUVpFIowW09hFiVa4Ol1v40VO0K9Q4ayzuwQSyDc1E1MHvvi9RTSDAxGI2/yBH/UeBhdNa
ZSRwe1I/NjM2j7EGhJWIUrMXsvnvikUQXR+yYsaTSeR8MaSNjW3sbolm6RZ+Dn+ZFY0Hsg23rrqN
WlYcyWilmpbSzjesqPPd3+6JMUOI8E4bGoKWhemdav+dfSyu8q1lyBdwAxuPPKpmHS703nn1kD68
KxJkXiCTU4c3nAvTAuYCtDd02BlsxfIrF+Hi1bet5vxJ3uWd7c66Vd8AICDN9QPeQYjdsrcYlhLK
k7Q76NolSu0l5MGgTPTbYURBonL8o3okXeZ6h2RDLUVpGIOkkNOr6M/bWcNlHgCn5irKQBhSOWdr
wunltFUnYu+wBONHR6YJJWsUfZjMJkiIKpsslZzLxJn+aEI6nLes1BPJ7t2X8OHNIv4XkM5gK+RI
LrSyPTWW8GckfLpx1cGN1cwETup/xGWq4mL1ap1Kuhq8Ia7/FRmCnaQ/JgZ0Dm5C+Cc/sOsfVQuy
lGP+8ZOCsCCVjm67zXryZQfJllw0PUMMr89m420gKLA0ie7OUWQwzW6SoXwV1LN2+CZ7iRmlP2v6
5IS/kKyk1MkxptMGGW65yjmXNX5zKdNY81m5MCduXjPrHndtP/iLcLWRuUxgMc7UwPlOjEVE0h+5
l8ukpP991Qfrr5PEjs9sTZmdEvtbtzIoh7g4WkJZLlUH49KC4abl8sin9u2HxKKXc9a8WNgK3nJS
ynhVIS+1HuR7gIA6LPpEP2/WgRyALIFlg1LgL6kBRTUf3uZ3tpInuDL8k+7dDxpdLW/+mXtcDmGp
9pAe/SrX2o49xEL/NEJ9GJ0+x/wfsidHkC+EuX0+v/pwfH6hDTMafbI2K3RNBGtzaU7RqlIeYA+8
JnAgYjj08f+xpykD+hRib31LQllIVOF2Sg7zqcXv0a2kgtqd/3Z7dqwBlrObknL0ySv4I791ZrQJ
pjQmLvABw8vxQfmdh7Vm3aT9VTIdk8FTor9C1AngwgfhNcb1Xc80a7urXo6qv3NDBsBOmEtfJZW6
qYSrHGY/HrcP84VgET2CEcxnh++CaYuusuKJtyvLqNOX1v2zo/Lt8VsUGTDOvushAEEXl+y7eqo8
SiwVkof4Hra6rAHcHeN7urMSt94n7YPko/0lksoVsJIEd/pI3XDgch5ZpBA41O+Tyor6CRzUoPX8
MvYcKOb6omibpXkTunfJHEPbX50v388PNEtXIztwRwJn0rxFY6m42DWKXHm/KKmhHMW7CknGh8Lo
uwlcdQRifj3RQM4flyC9NnSt6kPbrEvKggX09VZv5N8DSzn5TA45ZaAQ4y+Ua8hix1sH2YNNTcmB
ce1ipoScLYiPYUeksPNL5bYLjoyCOdHtYuRKBbqa+A8GORd+lBBarcjc+6arv2XniS76X+IAcz5F
akcYd+QsO3jW11G5yR4WoGcyLeVIFMbbjt+SK1YnlzlnZZ9cUKNk94jO+xiMw3kdq5g4SHztoMJV
aSh3oopaeO4wBoRYreOXqUG2YOK8QcI1TOzCXQi+YvHlgcZOBs0ATwnsQu4fQr+Y2xMjCdoK7dWL
AgHEKOLZ7KW2iHJtMTnU+Iyt5ABG3yFk8p+gnvvxYMVtmOANzxBpVFZA7bzT91i9tMY0zdtbL15Q
CnCpzbf1GVCisDm04E9GMOM9WK0hN5Vi8OikGxsKzODKar9OEYUP+OVI8PRk1F04s+fqrMLYRhBe
91uxD9549SKcHqgVknHVsiDtn1IbLaw00tuiGIJRV3GwXATNo+snvSSfXMdh3LRIc6fK8f87J/ig
HNw96y+htxnDzHR5EKgJbvs1JCycb7RgqNc/SrAf655inCk9DBIYIAiL5GlJ37o/w2htGQLvXA9P
0hb55K05sM4+gSjX7V9gv0ANCZhN4s/lP596oUXwWzVdfW+1EWK6Bk6iLhQjlPK7/yMSeLses0D4
iWymbibYBsTfk7DA4xb2GMkbEw9pAT9QPLhig3SltBF4+4sUuFdYY29bx3aQYWcoVvSjvfjr3uD6
9clUlX+H9eTre3kpuTvugPZ+cg+0kUv330hj7z66RDBaDWekTcoezZ7r+uqzeoWZaAX5RhMRlXBa
B5jvGGw4P5lPpc4iYOtju6mcQhxEkjJj1jWIBwPJEW/hhwdw9ZkSoQGtICiZ0l3qOHKgy+7qQtOR
f0icQiQJ/ZqANbV/CgCHELofm/Rb4gX42288AwiIqq8wxlVzQlCylQhONxpcjrJ5K0PcaVf6bGER
El6jeRZJ5EsGkkR7YOHUzBDVHcgVZKDrVapVB/ddGkjk8R/UBTMKmv5hCMgkms3dR9cLwuP5rdIQ
qKdn78YpMyJUVZXEetdZDrvmTCv5EBDzawfB+SSEQT/cdk9VlrZ9b50jQgzkfHVXitjERAUbQQGh
HWm+G9bzwWTuea4M3T21dFwQXN66x0EXxOME1REfosYaBMYqcMj973z0nJgaeygyIAP9CABut73/
VIKGWVRrtl3lj5hJnMt2Zg6RXQS5WR07sA6SK5Jc/7Bgo7cv+D4KcBe6pJeG/3L0nRAmXmIOA2Ma
zj+dvfnusgifAtY0+Ki8tgZ2taqD7xhXfZq8iJtKRNTcOGIUwc6XL2iDOlFMxBqTF+JP5MXRZJ1D
KnVDDWroLlOvdBAqlNBPdr93dlVALetHU0fK+bXgPhJn3G+BKhsIag0+16JSFJ24sB+OtcYqGIAE
zCPCpvaUBBYmhBdfR7O88voVinvje37MipFK5pN+gi9FpRYvGscvkvy+UOY+SVqQi5o+LXTtneQ5
UUDkj5zN1GZZzy7ZZZdg55oTM4BqMTV7F+wTfk0r5fVYczwZghw9HOZGwX9+A4IByUj+lDWcnZFF
6GRjjbf4PZyR4B6J6fe/vdfaG7xriqAVEtmlbe1QTwuT7K836/Gukaevt5ZRTr2gtQzx/3WJnSX8
toIenPg5arLsdIjDkAXXukv+ZSmcGwDZNcxDTdwXGFrq5uJ265d0zBXLZJx45BHs8zEIfvYhdrMb
tLrKVqVJif9AkzBfHnCEEJRYcS7kHQn7ezVB5rCOxptvFXqaY9mn4dSFN2NjfKFZo4n8ehc8c3ib
Ag6pVms7yvXGLg9CMipDnMbf2fTHuGNdDB7wzkwVD3lvEkn6c/htqhdQFfo7Us3DwXABgayofN4t
E8Qxijuacit6uUCxtlehxn7gl3OWY3gpRpSn4i7tkgFiH+TKeHQ3nJIqvAsSII1+XfajhsBHTEns
K81/lF8j+GmjTbCP6WMhJOHGJynCoubOcqam2tIU6YjBfcbLWtFdfV0ltMrGMad5V2AFU8YbcVHw
OjoaEnRJ+35rn3DPBOZUw9HtPJDSaCFvgSiywHW66i2pyyp3PGrBvTmac9h8PlmAiWAoeqVQYfQI
q79/fGRQNG0AT//T0h6/yjkcrFhMMuEEPNK9TSfou2fnq/97LcjoMwsOIquRM/VSjaro137FnR90
yb81u/9xSQej/S7i4IliuO2SGNiN8vMmN0fnklg0tGJzpTYwJMs3uuIKK47TzXcWaYAen4QIRWpt
WG0Hkvrcxm2c93CiTs3dqAhn2EF77TxCTe/1rvWwJ1QDmVEJAKZRlo7GlDhsn+uT5ZYYPCRMHdpP
QV2x002sjwjPXXh+ADnKOg7kWSUw6Gmb0CTTjPr6mlwKCoORGXODrPzp8xJ7fu2jrk5cTiTo8gBZ
vA4geh2xD472b5br8HoBcI882LUgUBxrQNnDHTWbcWTJx+d9buaBsG9ucRBOaHoXqJGpZYrCbuco
3SgV2zNw5e8rLe1/Xt59T0ZIM7YeycszZl6ffWfvIUmNiioqZDcZZqS1J4XY2PZzlx0k3wL9fxFg
Q/Ulh8qD2dDaOijc5Qr2pnb3wH4NduIMqW+xMdkb+mY6NDmqm0Mo+QelIPtbMylg6noJ9vdJNgP+
ISJCfsFrxdFQDUxnrsdgSiFBQVWB4EVxVBIzCQBf6kTsgU2vZM+ooslWI1+4hKi1XdMBQ6rhXY5g
c6oZMoAzF1a27XfUxlL5MdbMJu8nmQfgM5CyldlgJgsYSs2Wd1pyifmjwsW6QLX3OtkTmYHzu5Mb
ShdsswF4jezwUsnuPRWcEWgsJbe0eU36xQYpFEq8xQjnwdriYklDkyhnD2tuSkcBJ1hjvLwxwRSC
s+SpA52/C/BiFAStclvjBy2kf5gP8WFvDHZHy3oKJhciltKB9fUAy1PE6TjrNA9pHWiaaSfWLOim
/SyJRXnk9bhQ7KW3jR8ma6mDtE51AwkK3tWYX4dw7APcOJZl/7HTdbjgGelOdZlGhy7tIVk/rNEh
pzBjKw4DUWE+U2vxHJ7R6AlSrZnZd6QBzXVr22969NAroRNmLdlA3laxyoBCSHlAyMk8fapgb0bt
jaxN+To4vNvTrsrrYHsi7sbr/llTXaiHu6mCwohEZEPqUAW427B3oM7guNf1Pd0eNrBoO2Bx+2kS
QdKey35y28DQO/m+lD9yLcYPYP2ib72P+s8PDZ4seMlw5J+GI2OigHV1Gu8A5ufY1mdqB//EfyAJ
2cmSW/LOHAVTloXUELjuU0CUzUJ7KB3bezQ/DFCgfFn1QtBq8Fnc3Jsotjp2XEPra319KxcABGYw
sQwEmbgpPt3opDWDdAvNXnvO2Z0blK28y7ZnPBL2JcvmrXsX3OTLRd+xGn4lkqupz+7wMz3vgEiN
UGQe8F4XZzmV2Wxk4KXncIzy31RqqmQYi/69uwoYnmzYAZXwOsWHO6zPQNl8aJ66exnpjzxcexib
DjmJOd5CDPe8bROyRZPzj6TublxavV//BTUkri34U4W5K5/drnkvrMBssso0nIziW/QX4Gmk9Q6w
QdYA648WceBsXX4mhcYM80lw7hoIGwWpg2LNwLKqsKzK/eBXIdplgL3Fx1TwrVTE+2or5ua0+2Y2
cSt0ikn/vqYiTVvirzhvDtDRARt4ryTspCzLSC0WOdtXhtnUeuaj1+xxSmCwgaDFVAV+EsDc1vZh
pZoLd5aGVM5gxpIwSO1BomlNkyROA3EHEDnU+OlNOEk0vnIjQTuxxlBRJ0j1M8Ew4FI0Ou0aeQ6q
EJXBsI4byyFUFCIcn+o6OqxyNSImtP0ub3jsMUd737QYmEvQPv4db74/nwpbILgl1qFlVR3Un+Ou
c4kFGIF8QfaulJFIVLLNfPf1MKkq/kbmK0QyJgnS0Fh1WuHiILJ7uT8KloWnCeEu47oqPcf6ut6z
OM/LxnDMkmmCs/PwZ46ivdf7is0ObPc82e3AwQQgVw1PD/ptIQngmUg83eADBf5q2jCPgYd4o8o8
a6XqHqXccSisNWVPDUaZ+qRbAQQfPzMYe4tjfAB5btnrVD71cWoKLBPmi/4PUPYMTKmorOLP5Zd2
SzeOydS/y6B4gOWt6o74G2jIalZ86lO4szTJvfc9O9cIYxkHZuk9VlPTovQqLjQXoiqOpQKONhA8
5oGlzYtii8CJDfKzNQXcwFIvTyz4mFxb1IB+/x506A5HQoO0JOam1X379PuMN/b+sKRrVVBEjdmX
Xr19wwZMnQJSEECI3EifhUbHwGwvWO2ZrF2sfzReB+jnn1ppFZ57qGl/N3NJpDjNLNnfdQws779J
v3cgqAzghduFGu9EcwCOFLs9UhBFslLJnG+ybOLCU6FqNid+MvuUwWQseXSEb/o/ZQTebctYCmtt
MhAVf1QNE9j4XPqbdI2cS8Wjxmcgkq3v3xsYkARL5/0xIS7h+OKdd/sdIr8yhsYPstI0sOmFwiz3
Xl6hDtinIRJtlW4twxX9a+PCU4nhaVF1XWzULuW+Pm4gjnBVFz1qbXKCZkBDCEUd5zDMLt/Q8EfW
8NVlSxrTb23aY4vZzMQVY1TnlIpB0xl6S49NaGiCzq20I/mS3QHPKn22cc26TEhr//x4yywG2uSz
vH+QQANYOLNg8C1CpMIc0tB4KGQl6FTmEsXym38BbXTMz/rNN9ZVt1FEcc0jhb1PWZJQJutuK/cd
hjR+Aoiblr4UDhnY9dhP8NaaiaWiyhTC02n9h0oQNwvegF0r5yu43FsrGugf5qj5zxyeuzGKQ8h3
X8ROI+w/uXpwaFCCN8HgUrE2kMrrJjmOjbKrjPG8Cs81oQh+1OJ6TkPsi8vzYXuUqI2SC90+ok1i
1HqF4Mu+BCr/gi60m7Xlq2/veoxEOtwaKVqBFsJi4v/q0zsW4j32XcKlAS42nUVTo5BTHAyXo76f
w10PB/WdMsEjjsAOnxs+8WMOt/vnTNGUFsKSeDacUR/2yEUij1cCYVQqfgy91WCGclT2j4hx6opx
McmLYOUZWcGzkkJ7Rj+13DO56YyAfhPOoUrDawaCGKOoqo31+L5540X1UklahU7Q5pVD6fTUbxnP
G422hmv83WI0S32EOINLih4ECifzZZdrdmeJKHuFROO/6nMQedw5lbuCBz/XCWv6Wov9Zr/pd6GK
0jz3cNgi1LWyGYfMLB8V+mNdNMrACj7Xd1gEJeALMOK6cEmmTwseS3BDIBkKpgTSUPopPd0OOiOj
opRrrKcNvSbo1WYU1EuVIv2zPuuDe49W2LrrvPUw+TrmIAjzatvd07jASChFRTnpHv738NuXOYdo
XrYFWa1Iz4NxxCqbxWWRCwDJ+4nfbJ5QmqXRDhkFh6YfKcLp/7tbAryN8CcLpHpu5zxgm0YeEQq+
427V4B4qDbERfMcxNYL+rSNxP1yC4fSj1m/uZqLul3WItzdRBVIpOHbDpo/ZWcNx6ACeLub9swr/
3u0iF3d2/mHX6s8DAZLQviB5beMBtJM3D3nCMUGLrMtVuDT41egDWny2xp8FL3Ml7UuMg7Ks8KNE
UYTvx0Udzzcdhyb8NHXJHXbbOMlKpSHuErN76Pe1cIsx8QDa/0lheTphZH2LV9OCjoRgMCrhIbMq
VHsDCrxEXdsTeIoLl6fKcgLDlbowADKlPjfWfjL9LkUNwF9GcyPRh6pr+UYqhVfnT5JHYnhVwsPa
Cim8Naq0UZKJgmyfNAThqTZ3oO9z+EBhMQetMAaA+Np7s9Ov0US7EJtdGeBU7hY/53X5zamUBzVG
Fa2DckWmlJ2HSVkxiSdK6YCR2pa5rVVwKyG1+hl696DXqnbua2VB11/djGs0CljkQNkI95AD+DkH
St/xvwTmDV6QB+2tsMcaSxrMQrW6nA+MFe1vCgvoo2TGeQE7m9Ie0L78SK5t9OBd98xiPCwMplur
esNtFy6gc4BmaochAyZ0L0DNXIzRg5Enn+WQC/mKNgDmdgUQG6iVQX9h9EJk6YbB3+PMdt3kvwhA
geCbEVSfMVKbvy4uhEGb2jxSfCZaS05vzYNmP6qSAFhCIQij12HNwfHFl+CC4PgjJbNpPbBvPgZJ
dJgulcFGzMMl1fJz5qMGGSIDXVouQKGbN9YYuVVL5sUY1fy8ybl91MbyqeyEVoiMmCaPoI7NjFaX
f6GeORA5OBkhJapopeBNWbgIst67YUrq5p9I15rXKZtMI+V/B0WOAoFP+hPA5bmCWfyCiT0Hw9XA
St6WMXRUt6srgX64LD0818ZUG0KALow75ezwJXGv9q4/Iqm68srHOZ6klLMZV6HlQfCBR/Ut85O0
hoJbqd7Wx7DqLB3yX7cNz1G9kn/zyuKo5JS5CTzCOv4f6E7LMvnoW41utybRuuw9NHeBCK6C8BJV
bSbyhSe094Mjx43NBNyosXHPJ0UgNnYnwWJ5Il/X89gt9tlZNkyQvoz6rie2u4ylRsUtI/QMAQpr
O+2yZWEMbTpt0x44b/NRuWUfj8qfHUKq55Lad1T7wBuEruOSDkzSe7t+eJeokuYr/QHYG2uJj1Zj
vus3Eo/arSBVOpTg8VkP+v9ZNo/1GKOUpwxhDG6nNZg80ptNYOVxr8Xb1peO5Cw+KCsJ4SlCfEaa
G63Arf6Mt4ZqqSSI+28QCxtr8uGmucMJ1gjLcNjFyV2Ft1WCM8Bn/lsKyx9pdxLSLz1UEuF9SdLC
13DQPiqXxUnhScek5iJIuYTvuLLG3+JPvCtudNNEFyOVNZBVLXXjNI98NfT5q5LXXA6xhRGFaYrn
eSz3MsymdRoLTb8oLoXgtyFG4wbkU3bzmywl2gAmDsdWHSr8G1Jl93myxp0tXqwYpAOIwWmnr+3o
prl2DAl7tSVhTfN1/EbN3erE/flR9RrTVVUnF7bNukfuGmuMp9IV93iqu/RzMJ1fXWvZW9OkdFHd
c3Kg5CWtS4wD3OIl0N8n3OG89zoOJCXM4QpSxdJRyaTS1k7PAxgmmKiUFJSb1vu43p6l/MwX2SRV
3NB/u14qvuIdMzMyUtrWJTR2YEUrZXa3e3ThEzpW+zOAmKX3kze1Poh7uYRvRYh5y1SWBet6P1o+
iJ1YIq4WDBjlc/yHpDnvv4r1tN2HSAF7/MAg5/Cf2S2/KUy2nTJYQ4lEv+L+Dhmk231RdEJKG9Yg
V3flJ/gidEQhpzSYxulkn7mwfBik9vGCAfqZg+KE+PI7FxgzQjL6PzIsBXytOLHehLGD6qwIsFS1
pp4O9tSkiCjWrqqP+XmixEjWss6hf3HGSMgjnxSbBr5RXNxzJGcxrTnu6C6cerpDKWuKFPXpUBK3
hnV3q6JEA96Sad1miqbeMB9OCKkof7eB/xM4IqoYo+kX9Qhkfy7Mr6T64FhJM/bEs1/iQETlrzor
ePJpZBzSeIeLqgU8y1/7gHz7FkMSSkCppAEkwavhU40m5AiBVTP3OI+rA/sqQhbq3miSE3vznOVh
CjK85DDoxAj4wEDB6/Az1FMRlL0L9q9t7Q7MU4I6Am+wPZbXDd3waQ+D86Kn/9bFOp2rstqjd4Sy
QiBnt5or7m0tn2bBlPVAGL3UJQ9IboTIbHAA3G8DvfWSYeGYc8GOuFIcivORl3B0m5+N5VbXVvs1
aaeZkmqCXEjAiFOJv2ytgSfyrNxylLlD0wa9H03/bYc7BLNE80fJlv8ax3Xpek4AWpmUqb22q24U
MwiKp+RCPY3tVmhnKlTzBxk61hg3FfDc1kieqp98NRHjj9d2QGd2BnLuGAfPQFZzajUigNC7n7I9
Y4Rl4xmxiBdol1b7nehyiaczqMpZ5gskHtlWnIjDPDsiIcoei8FWe3pYhBdR1MPqSDRyNae1vnwR
EYoC6jCF0led2v49st8+2JY+e8HAH/KGbc9hQh01sU1FjhTpVgsF5jnpA9JhbSWkl4TGoIyS2T9g
94WEj2p+c7kpS2/Qv7TscU8++OagZwaqr7UQtbAXKWLwTeyBlA7N4oIM5XLJuKVGMD9K6srAmwpb
DEB/W2idOZ9T+u2MNbV2abHpMBqv94b91BTNqSFRPiTkU+gMOzbBTOHoy5V2KfaB2c1VGsqNwrft
cGkB0IzPN6ZVj++6BZ4+4KyPOeARFOkjmRehyEXfRruZOhsd54Rw9iKnQGLASBuLlxejtsh/ObXJ
6PgRIVzusYyiMJYx9cX1MWIJ/a+h/HZZmrtIoExFK6mqyTQ+pS7a02QtXzUTJoSZxAz7Rg3vAKC0
MQu7cgmE+6rRI7LBVXo0i59fiNcLqOrUavM60AJhFIKDTrfCezfjzrWL0WQnloCUtJjfyqj/VcnA
eweq+UVNZwsScLeWScg2FItOVdcC9PmSl4D/9XiVNBpP4tmKRWuLFMYMF8f/YwJhzyBZU+EKOwAw
2BmlgZBKHdc+gkx0scCdjX/RC3CFvymRyoeimF+06lVpR5TnnkVAILjVU+IS/r3LAC/6kz6NF640
rkutJuQDpTgINWs/MztdyUh2vSJtS85nMoAE8iEs/T7ekZx5WrcDrnQa2iWXeouZ9AtGeltXl4X3
In36eHIZzQ0Hs2q+3b1KOuDKVOvGyYkkGLg4UwVC4X3GlaImzR9Am8lNs7dko8K6kIDueRRIZpGt
qhG0Lu1/NzrB2f9unH2stsfkkA5+ZwwRZVv7n+iZuh0N5WYd/L+v1UN7L0ktKflT949TWCkhIuEB
IZ1ER2A34dW55cvMC24PYWaPQeVhQt4QqHxqJK82QnxBnYGfe5JGojwpQ7yy4+iDC6ATGvcOopJf
aA9leUJKAIGaCDnWe5HnNrjoQ88JaA9gNUF1kGaR3rhZiDxi0MjhvyUd/7ir/RlRHetEGsmb0dbR
ovN6VO3xPzSHAt3/CWNSF/ihk8wy+a0F8GHwEqabHPS1FiIAErfowYLK48ACqxoYxGbWVvFloatz
ARRfqwyuKaAIW5XOu69H5xtQCtOlrsQct01suH4VLg5b5XdSng5aBdMghPqT5jVq51c5JbJfGkTW
EZIWitWVvfZ9UJCf33du+KKFgBzDd6n9oqR/oz+tc0dmw+bW7KFm9i3GaqlB6ZPifmCOO20OhPYS
pGlIKt6Ktln7ZW8s3sqxPz2QQGzvEkxGCOy8lAzN/LeWRxoDCB2enTFR6Rocgpp5LSg4pBKTHA48
6UZMc0jhj5xXwhELQWNUeYUToBsZC6piWRUgb1Vd//Nn1pwlu8ncQiGCc8ouEUlgHIk5Jk7EbeFh
hpLxv919B/MAiJKB5twmhyJ4HiiiRwMM/mnX9QqBu9OEcTKZq1uUyiBn1qsBwncwHODYz5i0xhAg
WWsE/VOJ9XN6QRIFHzo3qeJlzSsq/SYq1M48SNIjLxPXWXHdS+fB0YENdYjS1POuotOBk65hNAcx
SiI3CVPapfgAmJxO81H89oy/k54284Ix1SJx1gyHckmx5+9YRvA2w2m7Aaj55bK4yvn0ePrCu1l4
rgMVnaV9uKEY18wlGyd/7CNUgUmNlFFPa+G4B2gJaxEM3KaCsC3S3twQVdMPvv1ktKmPCWeKXhIK
wfCk/JT1Vy73+1HrASIYupsgFoVJh9UKZpPc3YhR8xg/PaWHpm2P5GnDdADhiIFOi1CTsK7FZart
lY2WTrDh9TFDX2fPxQRJzed9qxmL16ZSPHBValTArMTF4SNgU4AEzhR0m/2ZyEEsMl2CHa/PR7UO
KumTCZ5b4vdhMrD/v5ibOY2f/aXZKrKF/AEBa5KwYp+ahsU39IG8efaR2Pti6xJ7UhwFe3D5jD8i
S/rq+I0LYb0HyRfWXYPFirT41iLSTU7xgFd417CQVrEZjJuvDqtdrh5ZSBnEd4K1HmeMzsOg5fd8
gXh2bXNPgmLSFAHXjlXRPkURI2d1GJZH8axILsBBiVYEFGICqmy2L5TdVulMGcbchKaak1/f2Ui8
npsObrTAgXyxUALNlk5WQ1B6ITDWASEhH+yg61waYPD+zK7W+6RCqkDwhDexfLTEOXL9ouusa9jF
/4yuxrmq/rTxG+V7JMvM8S3gDhRXaNctxbZtFj2SKq+aSueHp+lXUlAT7X6NnPjbJmMhu7EsLrzs
GkGVRVram9oeWgy+F0GxnDO6BfJLaEboCPc0j+MPNuZQdVNfHrFdjTTxmthmSE1X+ZkXguaD1Tbl
AbUgQp6se5pzKr/rKhVvhcYsvRMD6kdAnfWheDjS77YNxUwaS+denAVEFl728za7MX/rY7SidLaw
kyIX59TEcv/qNXI0KFJJcHJMjxYtTNH2lPNvD2sfR2AyKYaT+U40NBWfAXEjrjpd+R/E2OIOpB9t
U/AKzoYg0Vn+gttqpR2vxoFx8+NaC27EVcYRJOjqWrzNRFY/yQMkdIj77V7hW1YlOKhY3gmWkU3l
OaPVJSnrQuJ4urRwJXyNTBSQNQH+ox0eqpUBntHKNlAXCUbthe/kDh0I8xOVytj6roZxD2KHjm09
tLcc5nkjlyXndYL/bRwWYMQIabRjtCVw4hYXflVmo7NtB7gxA9RQgAJNjBGDlm4iYqNt3kMIEF1Q
9kqTtRCpcLFMHsaQ5CSEdkxOCkytvbjvT+7hW2MKmUHyBLjySjbgiLM9cgsNl+6J3RFH++bguvbA
BaVhABMyAsnGUhUSvx4q3g090UyJFUJpRmgtZDC2zCKI88AP2gw1jtdhqXbzgdyvPTLhkAI4zt3D
0bcdRK4d3sQywwyUnOPwE6/tlIAImQG0ywIYtqd0Oex0OMSfGPD0cSEU141k0xRh4T6k98LWo9kl
CC/vg9chfOg5L6j5O1iMgrS6viBRPEgOtrUia3yFCiBhP5YzLZq9+zuY5tgdGGp309a9XXwFwwCO
0XWaseClL/9Cy8qhlWtJbdsdNd3J2kmtMwrBXa9FjDgwutuV6xREQxw8MDEanbpzcsaFcSmfBZNK
/u66O4R5DDSivppXgek1cVeErx+xlYkZvd0gLp563mq1B4GHiAEae9Z9I8GqFoO8oJyucmkOWx9i
miIXthN3f+ZnJ2YE5BUvbDppba07ALZ03MzXpTl/PjKF7Yi7pMVPbWTRHtIcrVpO0Lqul5RFxFqZ
3+otL/Xy/OMtjBAh16qDCh5FCYsAiXIUsh9KJsImlM3p3xB6tehgbLAqea2S71f5rtpBL8Mkx9fh
5nIAn+/6yYr0nd78lyNZH8py6W6it96MiejH/79NiloRIiYr4cDNE6L559PpCSC7fCQ3X/l4RoeU
MyQslPJsWpgTeGoqTvT8KqRfaumD4W4AsETD9UHX3sNUvrNx3uIiKJ4b57+OiDSuYoHgcN3OaLom
ilV6VP1B6uW1i64d5bKsvVfcMY0zVcg6OyTO57OalYDUeU2MF6lMes8uUjvnyhMoBZCeHt80FLiM
CMuxKb0DXj9PcEcZL4LNXYtmMgyVHedip0yXM+NkWv+T+du3cregfOGrX8De2Ihu0P+xINjJk6l3
uXQZ9W3JmfMSBPe+aS4jdnIHaABem0dCVbjFH6jjzDhFppRvlL8hjGKjB05F3q7baIPc3QH2DtkV
xYcmNsVDQSgwJSSWFp5dysVABYmUEAR3qa0hWwV9JVoXWPPMqrjXTCnkBfY+cEPIUfnYkADWl1Lv
JFxH5bsdwTKtsz1hbNYih08FlusFLrf34Nrk6gNmJaw0V0OUUKbWJ5bjtOt/1n/KAQSgGezX1/b1
NP+1ZW0sA2bTfp3lhvs6xNRw4ldVhE0bIRrSXTAC/2EvmPyBH5rCNnxsipny1pJKaKmb4aAfVf0m
LPPnunfqYuLIqaoAxx+R7Fx/tfD7MmlF8J1XdI/m24mOM1f8lPwAbE3hSdlMBgShzzPa0oNF7afH
mupu8vr5MLxD7unjWUGziREXCy9HJXUP97dP88RKKLCct/KDfdSd3n19ABsWocSrkYelijiwRrMd
3+fqJud2yF94ruKyDWnWVkmwpqydwdVe79Rsu7sjU4zR9BHXb9pLiUVN0VhnycDH9Z3NaXWieqF4
qlEOZijbYzfhrsby17MZQSzq53PInMnywELPGEYOhHBTNlhCzxS28ASZM3f9+Q8XR7KUhS10AKai
qhiq9HAxhf4svtKWH1eF2zJhcJ89uXlssgDt63t/RVoxIDH5Z/WYXGweX8BZkpVPLfkVJgDp+zpZ
LjYSS0f3HcTW+nLEH4Q6bS3ncF3l718D+92vlSobr/44hNv5NCgWIl42xG5KBxPsVIT343vNx0PX
9/IllfHUKvFkG/cORx8+xPzgRONhTc7xfIsFIbbnAjmKoFEvnoVUV2cH6j1bIRgo4GRTgseDfKeU
z8kaYfJ18futi0lXwDIeQV3icJrH75DGDMd5JquJ3xN5K7lTqJ4PWlI8uA96cTAfFtZ7xu+mV4em
JH9GsaLFz6VHYfpf71sjUbTTU3GqBzP2NWXvQ5iZoHwbgtlX1usR/WJ8JwQdcKwTtqss92GFmWYW
LihpNxYy+SfdfSQGc1BR2yvWa5YylDRhI8AFy/QV/YaasfkijTvLjb+E/PewEGzk2pYOaz5156o2
nW0AsRKOT4hHIStdf5Z1VTeFmnKMwwcP1GDzrc3b99EgrzojY0A9/38NNc72u0I8+tGohj5DJTNw
QBbSC+Y2QDB181VNVaN3uN1puQVwUUiAU66fW6I+mgZEbO2B6M0n9K51ExgOGHcLzG7xqX+GlDVn
6dezhQkce9ItZq82vUjr+0wtHbIRuGQFIwxg+xtaSnoXlcp9JDT6KmYRxOfliCGNVzgiLKC8+GeU
X6sedLxPc7TkYPBZpdmJ9VMT0z66h02tn5/bXr4sjiTqi/wbqeRJNFqleZkvoErIhTazkDFR1Uqu
qPF8NvtDWWLsak5xqga/xBLEgzFmeu4qVIUOlb4eHIrZjOfJJ0LXjwkRPUm3R7gb0H0EQp/tV4ml
XZEe9NsuYZcjbAW89ouvBZIQ5e5WDEgcUg+zHz42DUD5sfjG7R30fTKZUrAUSsej1Tc4udRKCHeh
B0Wr/NbEa11Ap6qRhRse/Sx4NSZuaztZA3MkXYzs+ghpzaygTmXjlOhz0+5Jg/OdYBmhcgBNcBAl
0pW8dUjATiwDYwi5rG80h4FATZGrCtnb0saUJPr5Nw9U8749JVwowoUtRenWrUFKEBc72Gcwp+Zb
kWc+kx9x90H/B7uLjqzlrWoNb/mWb3Rg7QGrZccSFYEguJ6VouZwMnDwElZ6ChH3mDAXA0VM0asd
kICJ2S0SeHLm4wD+IkytNIG47juKJ74GWWdtSd+po3uhe5EHUyApqKclcot8ONEkhOCiahvqQSS+
ZbYre0zQ/nFp0F/P20Eu8Fe11DWW7exw4XqxznVYQncVeiVbv1hajDtPbOmLfT+tqM/6Q9hZsiYz
elRreL9yxsf+1u/T9k5B2tsWx4F2vuM8qs9nVqjsW2evmsZp1bDY1bXq8JCdDGi02NG/yd3J8XWI
fzvA/lI4K2eRnCshYS1amqqfebUsMLng8gFLh0wOv0HQfAk/1mQwjylzYOgE8DsE4F5B+TBLcB2z
36hZawwpmlEcrGdX38L4MP+WWB+4ko4H1A+4nivaSCT36iKiHNvj5ly2fujSPad3iiCGKeDk+OMZ
HgbufhIndRkBas6EB3MQmrXofJzxdxnBw+sKur7vPtXepDLuhDp1wpCJYawQMTjd1WqFhO+k28pV
By/TVRoAQqd/YeoeFiPooREP9DofsWfePnF0uEx55Lm0LuHzmD9ROnczhcyB0J7cKV9iKtfKakhN
WRFjxG7GHPpnGVya73BT2cZh5Hta/u/wCX2EidlBHme9YwvFeY31c+kGtCq6PusC0kDYlyDaCnIQ
OKhlbvbCZ06AXMnk8XyCeij3xG8twOm4fNMeTCn8+DWtZRO4kEcKJdQGi3+WAAeQJlRdhra4gReT
GByTYEJalQJsbzgBzRzssOtpSx6blJnQw8/x9RpeQNsTF1vV9m52CvNAcYYv564c8IM+ej3Xe/PV
vvxObdfF98o+W6zch6fSATiYhAochxBV5jfUHVI4XcH8J14S4gxz0RYVPk+2BVv7wmR7Q4v2YiDR
DH6zj1Z3hDvspdq+VRu4h5oamjpziA3ZmRBNWEbEJ4N0Aio/ek+dMoVW7pHo+vdQqEJOk02dQKSi
ejUn/DR1kv5JuVDdtY3izmstBa0eM01UZLXzTf5j24uu0Pp6o8r1+c/ovIRNHk554ba7b7VFZoiX
jUJI/ZMq7aALWEX1v2DonD/vVv8vIlzRZc2Q1A94DJ4DnHKVGrEY5IQ6zAVa3IlR4j7HCQ3Uep6X
r5nPV0EoPEdihcvn+wgu78x4jJ8yJgwnXHnUvvxf0E01SF2VWINL3vrB5WB+mOezoc+KdDjFsLPc
a9YzVkgg871YHkHWFnz69ys0blUv0MEp8anjS2pdRI4LXtIGZFj8Ty3pVIrp7khG4JF/sLTBHHr/
BR2o4WolPdehIoJ4fomnsZyF9oa5ix7uO5wT5omiKbBXTpvxkuZjOXf/BXn0J5B3umKWU4pYk1Gy
AZiqIsWOAqpX4rum2s8ltGdlLLyvtebXh00Th6rGKSWtnazBATwQMEQDlv/u7ghno94s9nqzRo0N
1Fxm67eFel4znjWqaHHcA7kNwLKetBNgqFyaf7qKN8BDbcZVUrg11WiKfP6itJ2QlVO63T4Zup9G
Uz5YAlxNq4I02kNLaWpGgaQUzDEo5ITvJU+HG5Uiy7aKNM+y/mw6gVEJLNAb6o+Yn6jyw4S3nUsN
6RktPCR7BOlLdwYP7FSPaJ2RKXhiMSNELjTj8Owpc3UE+HsG77CzacoiNYM8VUK6VJDk+Iekb+Sl
k8KFKMp2IAzCRxFnIL5vZvWVJQ6HX26OpU19v6nOUDYDWNMVn9A5ZiOCBHW4kZMIUnvS7b23IAai
ZzQADWByP1/lqphGzE3xETvSK09Mfogpd4pqQAPIQn6RkY4j+hNT9TIMXznNNT9nllEwUtc4qJu/
sLuT7T2jDD7fpCpKWgPTxUh7Rq7TA22gmO/XMT5v87zHNTG4v4OfNFPdP3D31jMjf1s+vo7iXFr2
USHmuronK3RXByYcrondod5HLVul0HbQasWDaOrENx34uTIrIep9N/FZDozetfMclx2ksBxpuAFV
UB9sirXKEgrsvg4WpAlHj8Q872eiJUO8D8Pc8Cnswsw2AIAwfZK/n+v8UnE423SfucMFjZnYbrKY
MYUmLT9jntD1CbeOlzUW8StdSodkpj2vaSSvNQNNOtgWCd1Xr0KYgjhhm6gKM8dYSgu5fsHE3Dup
Gw2v6kXoTKOqDO2PvM8AzV9ZXlaHGBYZaqLLaaaCbyyI1nYJZtvm9bDyV7kPqWt0TZAHx8Rb1oK5
HDyWDb8bRQipHFeW8KVifjvtmXsSz6EnuVN16ExngB7hZUxOTsHhUD0/uhgeLtJ8JEnJfpk1Y/aU
6wd6wrjEHVuY/RCwyxidON0kImIsmr6qBVbgJI+apSutdwe6cpb/ET43HtrtnCFV9kNv2cBaayPe
smcZlr9NOd4O0lypicPvqRPIE73b/C98Q22FclSkuhesih3fj1/g3ZS53YNvbQIwwtKqmmXhu4jS
XwJy80ur4hFE1fT8RwGKpgO5iOyTf2kCEQjzjrc+52ZzOLw7zFnnfdjv9qpkWUYik84gBv08rGgj
/5LGueHxqi34HehFO3WL226fWO+yoszx4lO+J73UpzUoEiXfIB/ADl3WS9Wn0+749LdojkSmqqT4
1gQlQxvXb4bamFP7q4b521WRfyT/nXSuAhgSNImoecsJnHp7ImwRSgHpmN3H4sXlECZZSuLx6Wu8
9WL7BN9sM6Z+XUIzzCkrGjeQJzgYNjjzSmF37JBr+DrCMmj1MPQYkcERr2KMjcij9MSFM/esJJGp
dYZs+azsihg5Hu+7Vf9BdiQ+GUdZaaht0CLqq3M8dXStRtUpDMuGy26DlRCj50KF3tz7dAAsL0iT
yBwgtWiGVRoVMiW0Bs0DSGuUnX0dqFCxg6TLudpLzAuAiQnAX17FSSC+UQk9z0VNKXZxjnZRuvJ9
B7iIJ03jxisfkg6R2bULhWJex5/NbjG9wL8VTUqLx2v5W8PnzYHQYnJwNW/7aoLJop2di0YTJcSq
lD3/0ZeWVBq49/GwZc9D2tekJop1Z1dNGD6sUzcytc7q32RQtHnNy7dD9K853HheykbEmxsftoOD
O+aX4qYhIqaVHcQSGdVA4q9Ke2sgMZAsyW2yElwlDObb8cnDGdvdJatzYKrp0Rns20vlSM0EmZYS
Zyq9WN50kl9lTNK/E9vz1G9KrjfvebVLtg1m9FXWfEg++J0cfaMs/+XbhoO2LIPMrVnI3XUqYg3M
61O1FuUygkCDICjtWyHOD30wMMWWytOibZGVh+RxIEECb2UzUr7HUrLPpE8K0KzE7HF/1GUjMq35
y1iUioULMJPpvnZZX37jgpLcMpGb3uYcNuS3fzwz4NZbFnBu8feKB7G8lpt/6j/KT1PPZ+2tYMhs
89jV+Hfib2aYX4rYS5AehyOvfEVMSpW+f05UZG8Hw8UMKJjqSalyRDs74Y0wLFRi51+WwyhD4tbn
JEXdTGvp0q7WcSdbqy1TGDHtWje7Vo/4Q8lYJOJ3dWMUipm4I/hPQCraTqg1S36egvf/oM32I6W+
u/0tCUwy8H8a0UBWrLjwUdvo1a0NrRGD9pPABCCK+KfUodybuaHa2EJV2b50SoMPKQqBSGcAX4lS
Zg5EXsQb9ow2bn+QNL2VJsy5GRpJ5+0pilM4f7wuE36uKLUNUuUxzcHl6A4Z2I+o0V+WXgHP8t+/
vvoOVBGr3RXv5XdA6cE0vd/DJ+c5jbeCboDSu18uk2HWoDvA7KM878X2X620SkCjv7tBTTSr5xMR
OJUQRxEt/5mp0ywDdJZSgB9ZQJwxEL1rHDZLinHhRD+Kn/AwmSKaOz1yzRSmuSvSLiNZZQGipv1a
IHS0Pm7rJ+dzZz/aC6Rq+Y7i9zloeOn60ONEAM/1mC5rx7QjuNt4yjMBflsG4iAbgS0+MYgQoPG7
LcCsNP+ZPGyUXZQTNwgXWQv91YAAk1h76Oyxj7PBJl6m6bpJ+J2/9EnsyhuKSN8dmxOU22n6ohGF
7WkLFx+M6zmvm3iFkIyqLPfGt1z/oY+abYfFQIvpwEUYEejcVwM1ALdxYmcI6+sz7vPjn6rgbLcm
B8a689ql68VMjR2enp8aaEunf1ZFAYfu8jKrW1AO0BDGE8YbxnDNy419EYnSI64udcmxPb1SyAqh
UBHuDf7QYn7zUGMfkrFg5J9rqKNTJomeafI1Y8UKwdTQTMq1AqnDZih6flDZKvEDD7UkMbT0D659
NDU7CgJ1y0rp9IgV7RrdbPahUOkBU4t70cJINa7qLAJOuLDlKW3nGzXuBeKI8MekalT+bDQbC2xm
XnxHkzgNGtNiIwBFjfc5NyVjoSA5o1f2O5qeRGvIRYPb/7Lu8uzqCz6oUBTV43AWEzA7NRAYSaH8
lS1ajz/gpQPbj+O5CW0/pAP8fkLPf1n9rwe79VxXv86leFOsfCSvEKe/5fbyM5kaqLEgmMZPTEkJ
Q3VBuizKk1XZYhOFgN/qlO6YErfQfy3lJwUIchBl7ry5PemZbQ4gGwxFFc2spagBcLCPbm+Yxemh
h+4P1KB0ja+L8YAkY0GiutO9m8DNzz6fkrjhUYE/GOhhXmhS/ImwKZvz4gClfkc0SDQGCsPDDP3l
LZM0rPjZeyqeffas8tScZbICtIkzRP6edipoPD5TipXNQoaSeoyF36HdqoyGZA3XlsQFf1sq5Mi9
jFPyinYLNkX15o7sgOUM47adDJtIsWWkK3O7NKQ0z7qZBf0v1n318b7QO8Lo99n6To1MsyipPNiw
rgP6goX089yF4ELDsDd3Nb/FLctzLpF9sd9vJxBGtm6C+rDc3CKVWxwC0o7R+RAq8MQnUNTPxr+6
UfdsFqUZ+qJcTBOwxSjvP8NTM2eH+Zt+w+W0qoosQoc0gmx0GlKMgriDu7ArBB83INtYPjr/e7Lx
AWT6MSAg7/bDnyfcxMzaYIY/U4wLRuTiXnw9vKj32hwyo9sovBNA7mqM5fqsf23y0mZ3TghZj2kS
BxrqSeL5PYCTG4wdD/u7CYsOhqgisnNyixo5cePYWmoEo61WF/W0fv4lqHsJVPAHKCaz+k3uqH4a
6YkiCJHDDR07BYn/tOx3uyZipH7uEyAjVphadttdlhCkHe6+Y0fwq7u1yva+IPuvkFYSrNWa5qxK
Q9qQ4FgkxAw0Td/2q3xfTnfsBXnw9iFjZtsjmfLTMsX4p7TFPtbVp3QxOMkQ692eFxC1S64kQmwr
puRb6KNTGrEQIvXkG9aUZzFXtVaXmoE+Lm0BN6mf0KlKWCFu0IBflEF6vj+ST+b8ZKF6usvvC8xB
chkzQjynrH9sbZQK7dualVAUNfPUNApzYmgJJNL/mVWcv/GpexzE3KV3PQyAf2pGK4xy5JFOKPQz
QdiuKB1BHc3pbSosl3v9PvFze35i3GztjTF0SlchUA2FOb9phW6Euf6bIqRBCI69cptKzxxuNLmu
6dzEIzBgQMfVHZrLQy3s8t0GgHYvY6lSZCI2CVPZY23kUK0ECpl7q5ZhWoYF4Q7c7bvFZSdDaJlA
pNNNqsAfxAwlbA6AXe/v6NCHcXN5RY84hL6gkNGMBGgf52VkHGmViBQ0ChL1vQqPZBDyx7XHZded
2FYYVh6MJzTwDXSZBryv/GIiHdSY+Z6m1Dtw4/mIyO6B7DDpoGQwNL9isYOa88ikNLH2A7ThlHc3
PVij/ZYf6+FuX6Xvqt3mF9mWna7428kOuaoeYYG7gosxKOm0W+pNyZGwPZuUoXxveqKoQnDReiws
9XL/PsPklH+MEDAPUQxQLqt+zInzJ0F36yu0k4j3qPEWu/e7iKofBYvcC39TwcSTVZ2I6AZBCTBy
vtoZ+Q4exeMbA967C7OSpYVaSvliRe9ChIXJ4i/LIN7Xra3F2P2C95qV6dmB93OcrugEpRcOF8BX
gBE4AiUjySP+GIafAqAvms8FuQHObfyZLjOB8ot5eu973aFUjnm3qQ6spRU/lVSvO1sJh9lFiN+V
I4bW5oz2Nxb54JJxnINF3DKxvChoDK2TBjyj4YAl2OTqmro+yihg2T0WuTJZAM4gLBDR2Xj/w3ER
FhXBbV34Br+dM0tnGwnvWmD6QSjbzhHeMiUJ+o7bKT0cvautPQ2td6AyyHXH50nxoZoBmxMNw28f
Dp5Cf9GCmm40L7AFTq+ZA9RGFwLG1NKn4PgVaJB96ll6nLx3g2Ri4meL1DIwsm66Bsb1h2vDYdk6
5z7DzCQcWSHvPhZzBXw/SvnEfVfGEY1oVJ7G0IGoI8YMO7IFr2WrZxnySeuVK1hvwyZPr02onslJ
Na+2lGhM2Bclz+lXLchkIAyrhs1cjYy9exSms7SB93j8ZrcpxlPeuIoqJHmqvMMtlfb5DGdx0YHk
ifjF4HJeEq83H+nZ+bNuw/zYhffwgrjxY+SU3haxUK/zuVK93si5FmNveEuSexNWa3r8bUcF3glp
hGzh+G6A5zSfGarDrpm71eerHTd6du1xd8XpR8mA3lfaLoNnwLsyAPyZp6Au+eCRSaoJwrYXzLjQ
EW9qSwn6Rar4NPk2+MYrqvZSy5XMAmI0MFeTB0FjrORKE8jK+Wsp29Lxqo1/idrL5+IzgjwhYPwn
e0uhuss/pPvJS78fnBCozmEL5qMxXwY1st0Pegs5L5cdyROa076aNRVeUPE2lvMnHk1MGRo9iGTC
QSZDQMOgn0AkH/i5bh7/cgzSWP32PTXNcmce00toxUagcXoi/94KM1oaZQWVv6wMncek++O5am6n
kp/0zIX4Jmz2MHvUkRGK2+DH5RvfQdahQ3/kCJYaYLNOrdhIMcpk9WgjXzrCztU8pivKpsgmdaZf
Q0DauJBVts40kVKZxnNOmOZ1bdVDa4ZNXVWEv35XQ2xM26pr89ZgBVdpxwvFn090ADmdx2HDRy0e
sugnzkRm9vlkYis514D9t54YTxKD/YD3IYyTKeqPg3K8vZU0J2n8KRE+4vgygWohBrdjuWxwu+6s
oKYbIxoMfVJKEYhZTAvHLMyhUvYqWQPkqrz7tjhqORXTGE5f5noLrH45yFOHUTPJZFC0nFeEEomP
YFEFUrkxDJPrx44n33DELHeJPzcLS/UrqwROJR0HVoDzIlPsOqFyMYX4gNVighQ6w90038yqJng6
fmgMixGnBR4afTb2oxCnlMkQk5ooOiVFRnDcNoew5bE4Zkam5nrQn8+GiosUw3XAyv6SXldXIw+z
Ux9LWD/0vsQFMLHsYSlroj0UmsW27KUqJ2rztZZuxz39wh1s7gFVJbrhu/PPyBaxpBN1A2f/k7PA
BlmJ7DnBvG9xZyVeGq6St364MQHmzDZDJL9/exfJgTa0SNZVKwPbSxlOfGDkM0Qf9+n9IiBlCM2n
j8N9tn9YGdBazO4N5T+wWISebdTWPFufTjr4yR1jeMz5hfK8mcjxKdUdW351/tppQCAzVCo0F47K
OeDk9h+X6CHdtMon3prV512jtYaGXfq43fGshgWbyX59hT2tbQicU/ljEvJr05ynCym4n7pLaBjf
0TjD56gaLwAfNG+Y85lZawwg5aTrEQZ3J8EIQWvnEQY6oAH9Dt1TkYQueuwl7t7LKW0xOPo8gvyM
InGzAruzEUgb5n1oeu/dJSFsspglZxrefawkP1XaVSdV0b0xtfOWfF66oMW8fJkzt1EP59UWgxBI
lMEDJ/XYiLq7qQcdPMo1NCOw7snBISApiYnYAIN/YmzdVBnukhyN9RZWI/8ADcR7D/cENcMvhW5v
vUBc6BoNtsQPsV9gqIRVWLjcdw8ly0PfYsAypgn3tEIqy4XRJst5i77f6LOWqboOq0LcffzK+WPy
aX18wd1ww+OtsNjichHdPpgh2igb4z90XSxVFdMLXl0xywAYEhmJnsJMB8Cv02aqUSUTRPkn+RYx
34Nhe5BlJbzm+NeE/q1KK7bIM9Xuspx6uYowwM8ve0enHn+pEeky+rJjueUaz6tNonSxxhHzsS28
R7oLzFk65+4iLBFNGNngkib0/ecsFMflAsGloN8vQvRRk467bh/E1cdQ54k9hfZLCVz6Ga+49QXn
4JXjTSptWWTJspg+ouvjTlsylmGR+Dqlv3v2jyUhHb1+hAW503U2T31LACM6ZcNPFAFwo7+oTHNH
47DZPi1OB8MewQ0aBoGojN2CHDfQsUj6K/92nHpXTzTmaNbEvbKFXwtI7wgTBur1pKYFtj6RkKKD
rT0U3qDiHw5i3Nk5A3t9mDMg1hEeFM2Re1f/QvhOfl0OCgyi6gqXnF/+E47bjZ0zr1eOOfqVSa8X
zjK9ZqdFpOEa4OVSC/3P6RgvU7UeLyp8Fgb8Ek192opvMcKhdNtF9I9HRMlAzaf/7ga0BvKRuhXN
wW5DzSaPSnSmLAWLC8LT3jaG0trsf2UObUg7e9Y96veaSYw4RMikyC1mmwFyUZqStjGlXNMnq01y
Ku2zFc3gZ381iD9Eh5uSzSoke9TTiLn+ktevKeep9wXQrNYdPN/JlvDsQWsYQzXKPhASAmkkgEX+
1RpJchmvtRk8WFkvCoqUmCbSPOdyH+WhR2xTO8Wwcb9ALE06V+gBgNfIDv2iBeVhtlhG8VkeuKxB
sIPGj2YGavimJA9DOdQHzBxldXSRHPmHjs2dTNFQmBbobzXsUbWEVJ3GOuwtYTbP9j/bqSBfpVIt
LRX2pmCtFEGXP5f8myMnVpCH5z2f2rKjFXAXqf7m3fHmJGpGqNMVymA2RUuM0+RThEgcYvm4Ylqc
AwHgJ8MaASFI6Z9VklNYDLqQ/f1zXueIToBlexAUcKbVXgIdLDilRQ2n3djGEmWMpXYr6ApZo/pX
pYWf0/RwUzfRvhJfJIc3BTBYonOi+8Ksv6fRewa+X0BmwngZJnP3KOgasy50JiuzCP+v1suMQ6+w
JDnyf2e+ttiiSrcYepbDtcXf0uXT34QafpMusesw7+LMznu8ZcTPzujOM24NftWVOJz3dicSOOWu
5TExf7qmhKtFRSeoyYfNYd6QA+O2eC65Ii6BCvdIDQYhTM2W0fOwsMIJIQOVMHFvkoJPnMrhBDg2
8YqSrfX2OUQvbnDwvnURsQdCDVEQ4QWMhr3p9tu3AbcMcDrhnqo53dQ9L2M4UtXIZPNmvoiexs/C
bDNdtY13hb49f+G10ZG+xlLoxO06BOZSn7WGqsKJNTrGzOpPM9q7EUK9Wn6S42M+7qs0QpS3p3mN
JK5UzNH/mro8/zqYssKZtb2GKE9Z40JQfTJKJeAlMXoLPmbyhrbdzuSFrcKEoY9IXOOjcY73s4R+
uYp0HBW7qExx4wNTis39Igw+i/cto3tKq8Z3y8SlKuIJ5+SUgq1HSQzY2YXup6rSXvFwCdoShw4h
DJPKIJWTVkgcAT+5gTvsSPod/M3ceI63jjIvI6aSKWYhBT6eX/6IY3Kgox4nI8brkb3tkwQF+d15
phvOtOZ3bjn7+VbCJNXzKacCQxHKgQRrVz/IK7urMhZpExFEetpRvGZRk7NQX5Mo85Jq0rQpfp5c
h/IX7KCcuwi3WpdLHu43wb/QyvFA79RshKXG+h5BLXg2Tyn3kv3bJzKMsBo57qVgbFGGwnvL4ZQi
gdCpPPB5wQVv/Oowez01MPu226LItBgnhLpS7oIxPMMHs7fonUny0OXZUbcpbx/e+BqnWq1NyN60
5eCUAIUPHoUo0rhphkC3Oo6LecYwNquQgFe7y8GdtCk8y4bD3BpI4EEuLQ/oLWr5oHr4J9bxYxga
UnBjnplSun5pIEi/KzigjdopcqujMbys6RhqUMW4wX0UrKSTAcgHoX73CWG924w+5djMW0Yn/wb4
Yz3mDX6texLuuXfQVVAWdQf+arUxDHZpRKE5wrqSJBqHvvCs3iGa1Yk4fT+DmY/jrVAhvug7nIUS
XJGtkIjlDZTDEG/fk0vQphNQPJfapE8N4UcuY+D5WsxOCoiT0RxZcd8IeNPFQ4HZSBBNTbnRrh89
bGeVyjflj6ArklQACBf5KPnNm4erPFKWTbf0428WsKKuyJgBo/9LTBZJHLv7jKSgILYMSmhXR0qV
eWvvImEaeE+LpUxkUkJ1CHk//HHBypdALM7X9Xz6FnFpMz5dz1DnxOrzlGymS6anyvig5rCbKsWw
CgK5vXdEkf7snU9dOJyC7u86zdWY8eI11R3j/ta0n2XlGQ7RH/pTPSs8OLJGR7O9IgxcQ7VBr9ZI
hOt5soh05Mx63tdug+KSkM7QLedmRgIBaPfxW7AbXI5NiMVEWo8JRSPj+JHNvRuaDr7iC02zMU/f
aL7KpJf+whCYk47VBObQAffUkhaNJKkEr+r/wmnl+Fii7Hwhq09Eqh1FnJlQRPoFHaqDN63RnRnD
WzeqzZR+ydbFEjn+aM4SlzBSuLe84iayJll6SUxnV9FlK+PuIH6WzqZaZUKOA2anfeNnZhMOg80T
C3VEBWW77xfOGIKNT+M88wkJeVFPhAAe3w/mhgAqy1XwVUOk18j0g/kJWCS9YHm0NJ3mxqFh9En7
4LpIfEuGkXdkPi8xXmNIw69fHAfakHpnjMY0SYJcgBxCPBbbrlf70/2rM7Te9eYIYa3MzjVVnynp
lyzeAtgW0JSerNDTUF/e77JJdWC4z1tzqfiEt60nhXFZ83WhbxOMnI44Q4WQZqJorLVj5FohXF0R
5McHbegncjkwAXdXJ+ame9iV0FQkC8egSrRFMSp7rzwk+dHRYUMxAp9WbDoXakxmIPFKLVx8jMMv
a2WcZ+kLvqB+Q7eXuNbdfYr/a+bwkHXRG/pmUDo7c+CsEvyGxCB4pUKX9Ouu92dip4fNZ099eE6X
ayrfW3z2FFlQrH+1QaCOESgVEhD8xBFvm2HmfkgasGqM0Ks4eWAiyhzOBwFq7BNc6ioZI1461hzX
xlz+76p0wYSGnw1vlDk2dCleOX3tRFZbPFrX2vTCekWxaB5VHL3Gp8LgJbDIc6Qya477LTOi6DAw
PlYrTANWgpf9Cjm1WBxidhOYPMWd95MOoeW2u0Xmm/TwdPTROLdwGEOAmjvE+bAp5tciJA/Nccpq
Em29i14ZiQVRp3Eq69c2Qr7PtgzjgBJ8O2RzAv/c6KAYmATBxmhd+CRtiRglOLMaqXv5SpY+CPDy
v8N+rOxICDI/YW98gTPmBtqgKuzj5kPa/r6PvpIoFoYRSm0o6X6XYl+mTflyfRrCNlSKlo0+YCNt
VOS2k5yKtbNdgbEPYKg/0DFo5TEP/omsbQ6gSsy6z9ffTJ5qUUxZ/jjp47z3PgOSt7UvyF+g1bzY
sp3m3bP+enTavCEjtt699ycAkTMR0VXjwZLqI93+U3wW8gG8Tp/d2cmmO8fZKi/ksKx9137OvemF
sqMhmT/tgujV5Q1Od0DrTc4P/mQusgqcOypoiRwS9a/YxOGkZ0E05OIMJ7pb607s3zGmm8MgzGjZ
xt3R8GtcaJ8FndV9gRuPMMNPJfUFgAAZJU3NNiMCgt2PcdpRF2RV78jik1Nj1jwmAfisZa5hEbNX
xhrwREgII/EMi7C04Mce57s7OyvsNP57RxmDYEH4Oj7FcFyVGwXgJFc4UI0t/uluzMtCFKbT4mTB
N2FecNHQKAuCu0/Uk5L+oKJe4+QvNID+Rh2FVwkP4Chu9S4Ujm1XCgTMhgI82l6uwa9LL9nf0DIH
VtiXnL4uEqc+qjSg/DG0D/0hmSl7rwtuktt+535h/4/YcCa8cJcO/OkjlYpedA/HcGNnITlTaJcI
aoDPCiBAWAp5fE/hY2H3WJf9LyYrkjL9U93iu73fGCNPJMsZ/c9W7D1fBals4Z5O1RGGjXkzcage
Mzxj8RtUOlWVIhBZzO2TmTCITOGsnuaPcmyaj7MKYkQZC3Jz/N2U/xBPz3fEO7Pyqu9o6lfLGtxf
AXDq1vUvxu6kAM1OH5CfnpHR5ah5ju/gvxcm4BT4U8wwy5iUCMQt0GWjIuT2ADQTY+gJGHCIHPuX
RGouzcRuMsCkX30f5d+OUKluQjVUHadmXiEsEoLGPT3VZmO46HO0wh2huQB0mpnCGVeBnmSSxifu
LCVIm7/Jkseyzr3GlIvtK8HnfedKDBiORYvmpe/1UX+ESglq072w7cv2htMyxV5SKtEmSh/DVbZA
AW9ArttJyIhu9JXX2hDXQoW+CZDIGr6LcvZfMWLmJWXV3FRKHj2pRKdZDiReBJG5gv2Ppo0V4b84
Bdo19L+ZTA1YqjD/evQPYqCE9+tcUlQabe1nwFIQDGrKYCkK4jpTGImWPtyyJkSejshnV9M6sqIX
dA/aEYP9xXR7d0P0l+zIpMle+MpA9QgKPYG00+3Y4wPW3XPfXfz3qVGFj22y0j23igW56mk0Vugk
8kxwjLu+Qeur0rM4QoYxX14t+lKTpxNDYI1v3vdKbCrFxouSlghGKeBWJZQOAYTJs2D3oJbP/ZqB
eNTE4EVZzlOL23bObtiCeTHvghglAPUmO4j6C3moOrzGpjXzPSpc2PhWVx93dFADPWy6AV5WK4OJ
PIcpJwAWoOS89BrQcOGaA8SgFWUEgUYb5F3ez5GV/Pl1F7EQB4DpeyX4XRXGbNeL8HXeARztuitE
pW8zbIC6Px/6IGRyipmyK1aW2ee474wU9ihsIU6IgvVzvdsgG+mQzYkSmaUdGJ16DxbAKG9y7Iie
YmDZArUUZNmsxYMj1BX5qvMMPpaXEllfDIuJjtNsoAZTxAunUxWi2/EzrBzU91/fqVvsIzi6uNAz
pzsyJIGGF4CL82n+hCvLySH7W7SPVmhox72vVrIRwRaewIINwbVQcKlLgsuIf+tIkare880VU/V1
OZbg9wHLqmeWusYhSxXMA62u+lwkGL/wVKKH3enyTMy6IQBMJuz+UFAoa52e0lVGaIxrPyhUz9K/
w+n6RUriD0mFtekTanUBqdGjHunJOjO5BsSvUSdRvIrCKCn+RB1XcWVe55TCUFd5PU5W/fktZlqY
JLw5EekhKfq9bL9wUW9wumaqX3YcoXBdFsTIN1omup5gXKQQ64d1UheXZvlEPZv+XifLnJKv+tbz
7upS1UlVvCNnqBr80RilXzmXCeu9HeOEYeRnsJWWGad56maAoVSVk8+AdSfPLAR/GlOGS4onxwOZ
CIs5Hf6nDgRlS7EGJx4WK3iSagGfZgGqdFuKhiPIPJ6mfG6tXK5schOZNtY78cLqiNz7Mne0Erbx
KIHhxtfRKqkfuF7yRJjVzoPDpa+ws7Bj7CLEgxBQCpuHSztbXbJPoWlaRFaKtGEdApgaGxbxfuqI
L273rKDB5vr79BLcUEfbk4HlTCnyyL6wdRVnZNs2HzYx+y8W/GtkU9j5LAkBUt4ufEg8Cvyj0taf
VkwgNvYelmRxTl95rj+agEBqtmqhEtJrACbG7NnApBwfLn2Ej3LZ3tU+ZzNwDy7YbpADq1jXdqcP
sLMeUqLULK5w5pOo2dUqiDuxBFhrESio+LCdO9N1tOXArPiDPJY4seakaZGgBpT3WdUpJW3kN1tg
KFCzLTjjeAISSXagVT0/6FxOSieMKDEEqfrttd+IxWXbPw86or/MMKPibqcyzNwYia+PVWxpFQvM
d+CidLvACkub99UBAY3Fq2FHl5KXgiphqa1gM3Ka5WYot/T0EshouzZ6lhL0Ebp5BlF3aP7dWQgk
UPYRqajT5/bocQd7OHM34V/pdksPZJzSdzPUefqnEs4feO8liEFhAIDvKBsToI1BYlGWZRdXtyr1
93L5i93HHMUDwpms/x4m221h5koSO/DTFTiLlswASm/9ugN7tx8ysO0V9CU8Xd5bnGGBl62TWKQj
+mHIO3tIAALDghnOK5IU3LcwhpxI/rq/QSuOhK5topEFcsdaF1uJS/jsbCIwHZTUvQwVhpcBOvC1
4Nwog84+kYw+ukkhfesj+xLl6oPSFLqjC80/5Pk3NUju59bWDheA92Y+49SN8wgX/tjzi3XM3ZYO
xF8eepTR0H/4z/XFZtfwN/u5glBN0+FFb5yKLZlJeZDV8CSUonlfv1l9C+eke/QYPghrgT2tDh9b
NnxoGc2VOBY23M8rVzFFfHCS+GPKehkwnKobXeYkrVuCgSQooRDK+x2Cyh1c5/QwYqA9IABGOff3
ZOiqmKWsaQR1VbL8CKKVrXBv99bl/sZR++hfZrWgT7cWJwCmwvxXzIWq5ZatYwgq/wrsBt2Nly9z
FSfTed+ZLG39GU11/n5MYf+XSBUwHLNvueGNFC7bTUr3gm2p8kPJTHqd0c2qDDZ0Dh5rbu8X0hbr
qtKLyOQ7GufXwNhks9VIJMvSyTufHfTWs45NLBoOC+tD6HLcqPuPGjNTf28kJdeOsRYlFil8uJwR
QwaVuSYo+eF5GZUgJmGYLMuoSCmw8+dvHsVA4wT04ZPWBnkH60lf8D/zxRx0qRsqfI7XplzJsDAZ
5GLuCom67wLLB6HIV5LfHqcKIZid3Lm9ZccWHmPqiekaBSz/dh0KUnsdV2mxbkbhOidh2/X2VxSp
StryxwDAA+kBi3DpiGgAHKzlyRCMkjydmBjespSZz8mTvesfZmsBYH4jU4KmjMuEUStrKUl4+t81
EC2aiCjD+gcGRTfeQWmv9WtiadA/5jMuRgglWKRGspWFWZYaF4IJfXdIb5l24sVf+AL4uNyDfZVK
yLeRYH6L+lHj6ZAR68L/osggLBcJ4iBcQ0A2DcwvqViPj1XAZhOWskabjoeFWInQ0xVHByOacTgu
/LL3dDQUdmYiHczqrC+EL0WbDXx1xLqgZwIGvY7kHCA4hDFYJyboh4YxFCvRdPAGk6+HU4pnOiwS
XVCZRPF0IyXqEVG5N6hiKIXPmWKosLX41ZQk78gnMP9yyarBJ5+uy7oLRufQKxCI++7BNKFtu9PO
HUPqccmHxGEW2RcQK2vb03qa+3iQlSJ/3Si7epk3N3aq7MhJF/wd8mFQHGne7chUPhhPUwH/o0n/
ocnUKTTTlUtuIfilIoVJZJkNAUcazJ4Pc19ldUcbRlaN4U+IsgGzRa5B3KxqnFuuOKmOM6azH3Zq
4NtD7lmLFQIir1WbzwW/5Wd5Skl+CEmXrVaZxs78Hya+DXej/ANE8nHKz6XMd+Y1279CDfiY7LYU
3Ufl3lJgJW/1aLWXWyt+8XDbWCs9GKTjpH12qt/E1lXUcgleyvHoTSYTbfuMt35yVHDoA1xE/1H2
A/GaUI3WenaqLKM+a/nArEtNTc1B7T/gLMa37RS63qOzJm56uz2O0omqtKwNu35YJjO9LNrIvwha
RB7XQVSIVfnz8IGUEeTc0svMSQ2zbE+qSf3NJtIZxTxlrmB092wm63mws63DKg3oX4OIoW4nIiSc
7uZIl3yTZ1x+4lb6LfYzfaLXVbeLUrJDAs98AvPE3+4rOjePd11pgvHhbq5fUPfbATvDQ8q0Fe8N
oAnTxXc/d/Kfu6uYiKt5eKqHXNzyq5nPztmwpjKLRFs5dLgVG2OGmCizW70tVSmkdIEmK3JAMOma
RsSYqqEIAMULqVjyLVK8BS56BE/1Qycxw7zga0AfpwmLC49adDDocmz7oBIOh+np0wbKGe5j1MFN
u1riMfMVSIfpFzrPb9BkfVDbwrc/wFoZlSf3vPWYsOXLd+YkvmbDnav0vaKg8vN+lBHesphpOT+o
SuOLdnxK7J7jXehyl8SKDh/UxEwzKcnn/uJplWeo3kT46zaYEwSNYZ2U6V/hUMehSeT6G7xk5JfV
hGUN6w77VHnbcP/vwPFDTQn6oiwbj1zGQNNljlOcZmHJSXp44ZXlcDJif2c+NH0epU/o0sPnf9ap
5sJiQsF0EXDLjxcdX/k+C6KqM2ZoXmEmqZm4v0TwlEDEkMTo+z6P8+mPZjR4NdAIfK6d4FKLowxD
/ZHdR7VHxBmw+mYVI6zZ7+YkRGKK/0L1CiO2dHEaXYIrfdwMxchCCR65DRWm0VxVTwJNcX2X4gVl
UDFsj+ykRJEYl0IVpVHLCAP/PVvnzFjUwJFvdG7aeGz1xY5G7e5Arij0ZTrBKa9dH1h9mzsYljFm
b9uvcJ+vmbPEV3R2SGM3HbniG/z4Hir9sqv2Ay+UBNgxRt9eg8B5IZzhLfff3BhNcfban8uvKzp2
Fi/E1ipKB7n7T/HjKPpBfGtnxnt82vAy5xp8D3RERTNQ3h9E+07Ou9Y6OAQd2CINg+HogPnOU9Sx
WUXEwyGKBvphuoh69V3KEGfw4BGLeAmN9lxObxrEB2YSW/dC6JXhpLjjkTXihnlheckLnfAlD/xf
+qGDAvbAlNn/WgKmH71fDrip4Oj0y+UqplKf6dm2yE1X+3TJS/nZ5RDVrY/pQQBWjZKNxm9D6Mku
XmZUAf8WrgDbhhvV6uvlKQuaRPJbNL4wJOnRs9SEoDVmDrcSAQ+6JLnV4PcQ8EeE3qQBS4AGXsZB
dv+DJoZGGqedtBU7mLXPAO1cm3mEMu3TNY1TVOCeOpZy9Rl2IS2hl7KTUPiLbe4HvXQHBC5i/LZs
ZRo1n+ZV6p0rH39PDRmwdl0yRoe0JD6a3LsLdJ12nq2obVQ4AXRxGIQyYZh81kYqAsYSTdDm9t2U
IzMrjLAIb+n1K+KkAXp1njUKbiUyM/s9fMFY8mwvN1U+hSMElmbIhRXG65UIpv+u4oIqOCgoOkdP
sBeryQDVkWq8QUzx8htxVDn5XDrIBymOdIYTnQAVt3/ZxCqMMuZ+/tUnkpi9tmT4QvtILwmJy/9+
l6/AR0j6Trsd/jiAQTUFsK3ZuElk9++Chml6QmMYcXeQK8sDS+iyfHeIPzektE6/j4kZujvcNIwx
yFSA9P2MICwye8aGe5oulyB73KiVAgRLUws9TU75947fzB03sib8ONSlIreE1rqmSjo1nzzO55jI
VHuFDm0J804pNBeigl6jkat7ysJMF1ZzJiIDnpfROIHT1BKg+xJDYZgc2T2/g3qvZetLMKrh6Nzu
Qw4M/PDxT6JKX7VyzuqkUjBicRwFL+phuBOryZ6qNGTTnVthn90kwx7ayONRX9PDpL0Dq0gG7hzr
teLlXf8c+q8NZ0jWBsk5pbKJnoGknqWDjbKPw2dQPSN4/CeKn8Yqkpoi1lg9so6FCoaAYxnBAxdH
QSrlJW9aJXb8zWyc6AyrikmTRgLuS9TJBbB9uAPBHHl9onjqBaATHyQJp3ygzzqe8+ezAE/+l1F8
VsHFr5NUIvZN7yKFlTP4ek2FNM3WmX8247znO6SnN6Fado8x/XYxSGgD5vfEXk+lm5P2xwIBRqkK
dU1nYaS7eyTk1ZvwWzCOxMSJ3sizuJoLkkQkUL5iunLN3goSRcYuA4lZZPbH8XXUdvJb8DnPErbI
R+FR5FYH56lGrzwlq5jS89mhkevBdIT1icOsDgls0FNH51N16pxO/8nEQcZOy7B6Lv3T7fvaqPuo
yeK3nt35j8PVdPjLCvln6j6ILfoZyT6qpat7tRBPUQN3nBjA/QKblvJFcqosNnrf6CILDi4aZNTF
nrsuG/Wn8mD3OHIqUT3+luQlkaFmU5asmCwVuBLAoczFFQlihdyatcyolnhgLRFcBy1XiG/DH/Cw
4ElpVIP0XepZXxtvZqbS1ah0m/ubHk3MQ1gfh08WC/mLsxTAt5GC5FisybR4ws/jqFsPjUzPDJJA
n6VPzqR3XG/dYXd3r5TPkkfW7vPYP2I8vcwCoj7QcwyXXzYwvfKoz9OgoCN97clZPK4GgdpTCp8a
klZblQDEFqgi88G2/G3veO2X/khhZuZiBChHJy9h5B1XfGpiTPelOMmBAMD8A3e+iPK6HwdU6xio
RAH3J7c0ewlSmhNLGmNmiI69UAnLiZE0SNNeIYq9Vf3+w+J6ZTLmIAAdsPOOWI99yKN8t9gSKQuh
4keM9QkvWz7k3kW0u2ljtishmEA44vBh9w+nhIpe9bVTAAc5YjlXsDuZ//4IJL+p1GJmUjmrJ9Qc
8ZtRSDOpIGM2bPBGqAgsLGy/zu+BK0IUYfLxE1qRn3ABJ0F73/hn9DQnczbPXuI6SyPSG9ZoZxlY
1Y1079YLGS41DlzV8XM4gn6T1+lJdSwQ1GfEb+A9Iggw/Rb2/ap4IP5s3Y443/j/0TnXezrjYZYk
ASybhBAOlOSfaS2YBGfkgkfRGDBpXi+/FJRJhtSfx+4mFAG0XB+dQjlHboohVSf310YvAT811eJA
D46yYFHef94Fk/tXbQTz/hGbTVJBByBChxNa8txrXTdQUe+OLWXB6p6bPEiTh+456NsS+j+67ISh
SVSHy2x9Hx9EKTBFnzPgkwVjghBdfxDGTi7Jc58uh9JQIQo/3VKybWGP0c9VoP8Z7Rc9/G1j+Hzb
FN2yyKN2jtvWseJjIDUtDeaERv2xRGJgENQbjVS/CVwvuD3lZHfTJMkJ3axhl3AFHzQqsufzxvOy
FXfYZaRHwydE5p1I0BkBE74veAUycZ1wcBOptaCsycrI7lDzKyX4rVfTrZyKqH9KghTG10UJK4QQ
+mP1vpjSXy6qzY5t6PIYJWlbW5B0ccdt5TzqF1bXGkOkpSOqsmeV8A60QdqpnSBS4aa5IGjt67fU
pQ8smcNDMAVjun868H5hPf6xKAVD2i7MBO4xHPgQkDHgKVsTq/bBGZODCQuCz2lPWVyYaTncj1GL
rmIyVFk1gVFDEa7P72CICl6va7CVJ7aVX8MD23iEikVVije8OJyQ7boCHhINuxgLoBaw/tnWzlge
CKFbR87fTIO0i/+Ugv7Bz5QPKKq2/WjRz+5aaGwGKdNGYR+g9eLIz3T4xQywAVlmy/DkxE9ksN0x
rSvl8rYtWDL76DiM/bRSZkBl7760UBJls+hftvNz4KBIOAjSKM7k/Y+jcRsPGoZRy9aSippF3V8P
apZDuW/ZyUdhqntoE/7Z6RPETKKfV1mQKGRC3IzCvzA5cn04z8O4GhY+oUKPpa2GBBW5gHW3YBic
aIGugbw28cSWywtuGdu9dR9OgHO1rQzUw8LpFqzxn+aRUCsU6JtTjO5hfj6UOI2dE32uotcwMOHv
XebqcbdnFEHj12xEuiI02+H1u5G5Gnc7mngq9bmFBgMdK8M9jP6v0scLTxY+9bmvJ03kcnLM5olQ
WCEzrMGct72ZdSetZL7j2JEyrAA0Y7R/2JKyVR+ChVEyIARulGevKKyuICtQLG8DvgW+H3MHdrBR
5q9bdibt/uKf1barUJTrcjXt4uAFNHl/TM49Cf9SX3PEf4uuFpTlO30YUN2FTupy32zz8rAa8YQZ
t1CGBlbtqKkBnsn3tnQRoMkwQScFqTopoy1fRTPImZgxYje2MVV8SEDGh34ZnkHuJFsqb4aZBLH9
QeoZTnSesgvD6o/4oWyJK5MvqqZz5QYIwNk2DNjZyUgeW3KiCPTb8bWlES8MXZ5om1zmPzmaTbf0
uMepPZtfu5vduxqhiAVsS0o66Dr90zKJFXhla5p/MwsBIj7bG6JwZXNuzhxHc8uJ4e05eXO+PCRd
8mS1S/VnVyljLdlJG5U1w3pJLanzlvdsxlCm7AXOvYpTbX4WJ5EEWOdc7vGcL/W5sKcDZBGZxvne
j1P0EI++H7yXFoCKUhCM8xo9N/wDqlpMKX6hx0uvxOvNZoM/QtCCTloJ9NZP8T2LjkEhrsEspRJa
5JOjvAfOPyEOCFEQSQ7ZhaaFzPIBpmi4aQy/UmBKiqHOnbsdH6DLJfyWrQNaS54ueDPcP5lSh1i/
L4WzE14nzeLj/Sz4SxFsvjResQ1zp+nxOdLzfRShKZEvy9S/FCN1mVOtKNGJouRBCESewN16OkMw
t1p7XxnWUaibs4AGAAcL5PXgIch94mX+sBPZzBiWgWhlnIQ8lowiVe616oKLICC+t9Tiuq57gTW8
aIP2+JvVxdQlL+LZOKcULfEyV1FTP2jT2Ajvw4v6tvkITRNyBZ2VaaNhrbo9f5bjWaovEQ80bc9/
j8ZQ+c8ZlpQg6RJLoBTKmS3z7sYXpLbrzoVKwSREgs0XZo0xTXw6vKsK01tj9Q1FyOGBUVXk41va
AMB09ya/uy+dUR0RJGRbu0M7hGdY/gNuwkuFueU1kb3iWYhL/YWt7dzg4sPAyXGXcsuMvSEhKB3z
koo1IAvvzvYKtSamTEecE7kLMcgj7gLTTJ1HIi/oYDI9OVZ4UVIM0MYkctQcKYXiaDZ7JNRI+St9
TPycaJgDkgq9Aa/fZr/CtS0MADj6sB3w3DOZnqCj04XzEC4xwnQrap2B/Yiyt7dPTKWDyGvLwOjq
zRwepyfiF5rirrlmlvO+brzWdeJx4qxqCiOrHyvNnFNZf+XkP8P7lCAG6ggJgiLsITp5P0IlKckX
HqfEHQuxgjz3765ojSYSjakpO9QyDX36ZdgUQk4ZTXO0jkx1LQVXfqilbyNKiJbVYzI4Awd4Yrm6
MwMklubHIsB8Fn5YMM0CGF35Z17fOh4N5SMW4zmWKTHPECPMjpP4dAh5JU6znd1/4J8GatpWvN41
77kxPTcFhYHTl5J0YlM88Qf/3rEPR18cdWyhh/qERWCAaWo30sstkhjEEHRGAqGAwX3ZJqm75hk/
5MGvjRhWS0nhCP+f5LS7Xjo+nguh96dzOwbO5u4FdlM6gbiVda1yb5O+gWlRpAqqqVQXArjeVp2U
7w2dqdI4wjWmZ9iafViYGQ+Cq5AIMwkqjAvjEO1MYF5+/ahwkQAjEuGJyY8wd8kgVxPC1uLI3a+E
4iN+Dfgzp3dwWA/pGrGH1SY8086VXv/1GmCzzxon5YMUSJy0xWjCZemzYcGv51XnxLDPqQLHFu0u
rgAZqI+2Gx7QDphQ5fFukEXLuZBHmUKAYeunzxXjqE9CHW5PGo3QX9mop0k+4qpfXdjWD3kEc8CT
A7BL+x8VT9fnBxap9iNaSs1rZcv2oUVmQRhsa/VjYcuDAKcvzsgLPZAlwvRDgYM4fqiUil9p8tZC
EtytavwBXYH7OUP7ueeNsvQIar0YlfI1IiiKxPk1XE9TM05tXiE4MdmmgKCeeY0c3SM6QKoqTkXr
uOd0jgeCxJdYmrdYsVEh55MxVXGFb5YSr9cJSAPT/pwVCpq4P9ehdHaiKxnW4JudsGj5MhIXpkkx
NhI6YfYVJT9EpuCoaqafObv82FWXI3TV1ZV5Z0pqfqbhwGP5hb6vm+aywByAOSN4zfjAXj8aGn2f
5r5lEftR0mIOsZ3xdfz848lcpxEhFvnpSt4iNv6L1ICfxOeCWSkvavBVr5kOtfn9CvPDpnORFL8n
SIJK/84ruHUnP6VmsbeUyvuBvdidOexebQV2MFaHQlcoCToLEBeVpPOzHp4RCBu7CpiEgxApcmgi
2VUKDVI4oKKhMCJUud1G7RUpRSNf9aqiAvWaeh7ZkbPvfOikRi5qFlA3yE/5VqgHEC28xGU7pdho
P4l+5/Me7nZtpn3cjbsYb8RFgADGWl7Wn5gXTobiYnxtxZR9jF0rKltPCsYLfdOT0wwitDd1l2w5
4T+F4KjCJRnqqUy4GXnW/QokSpLlpU/8ORIIvhit8djXtPGu09fOvLP8KVVwpW71NMKFgho9ls39
z0SbxXfQm4150fF9Ko10nmLV6mqCQB0I0rnXaGjnt4lt/PdsjhnjJ7LprNhLb3PCje6LbtBIkiUk
9IDR+st7HXNU7FNhBNpVSLDvTnv8CunbVifgVp5acQqVs0KuWUzJtVCEnmWwGoS1I5w+lJbL1P6U
r8gG47utSPBUBniPWdTRlbsS9Jce19KgC0yzOYl2oklHjO6O3y1jUkS9ppp8Uf1AaJU8x61jF0Dx
X/QjCawg8qMMIWxLyoumOVfeL4+EKyzm4XtVY57+j4KfqnXI9L7INWK3oTipm9KawsGKC+r4nhHp
Knv7vH1yEvJ2Ppf//7JLugBPQ5q9kkUQrFuJ7JKfAXPDsUB84jX5VRe4OFckSV6gub6nyw0RK68q
xgk8G2+SMDGuGroVw/UumceG3uBjLF+vkTrewnxJPL2Gv0mCCC0prC5241WQJ+acLkm+DpBfZQlA
a5NoTwPVFpssxda2Y6zAuOwZnwJuuiBiApWY8T2KHPb6wyf+aG4ospbaHSAsaYskzeWL2Yyv2UEu
nkvkadZlN5PV+8xMDGJTqB9CZErv7AVR/ubpLR/YoxQCedsHYW0gGWIAUimQ80X3EngjOkSCaxG1
xg2/0aVrkvWSGMB9HBVjY3x5jwqr2ieizFlEcOQTUd2Xhfl32pvdTC6iGxwWSBmi6YG/lfQk+rCn
pP4YPyQ9Zu+QATVFgPM+9clhK4rGobXcbN8iRQQdozboUme82rx7ljP1rCBVFCyKZC+j4ItbLHJ+
vvHX8ruma8hvGc2g0Jhjh0FvLwdbHdjbsGe1tFl2UpTU3gRycgQLBESSmspBRg+DVevB0mfvLZdP
CCixZc/vggAmo7sA82eqUK39IhP8w+yotYsn7g8a0DQGmfkBgO7AaXKB58oMKFZM3wceQG28qGC5
Vgt09+8YtqVcQ+8LlRcEg68gMIdOftRxjLJ7NtNAfQ43T5PHhdv4v7lVm1/rwA3yUqHlPNd6lv3I
Rk8RZxpKqQ4NDBF+7bVMlnvmfP4bsIKdY0ZeisV6gvc5zKMeOexr7gVrZoBCA2LkUrODJeGGhG9j
1T8q6O8/bh1gBOWoXlxbMzDR9R+e8O/cf8DFryyYHhMVQ3ybJhY6qMQYUZ1P3zmqFvjsJMlmFZyZ
CQ8Dvmj5z5s/2sGYt7cHQol3dtiSg2TGJzvNsdM0wwBpenxGJ4l+VO1deTspsFoSJhY5XI32IiUM
/Qa9ZWQb0bdkrQwdDJNmkx2lzbszjlfKQ6c76k/mb+gimpzjAUSs0pm942T6GKSJU02Ck2g74KLU
x5JO3ZF+GwQranWtjY13Khis5FRmPpi7WA8WYFhHyhI5bGllGiAB0M3zRTRslBLrTnNrNpJAIdXe
Z1qm9AAxF6P8aO2XGsH8xs3kw5Q8xGa+JdVn8cGUSMKSNezK2OF1pk4OhnZl7qUIFYTjq5cPIm8z
IUFu/q9fL5Z7qqVFMDGjGlw2cFtmtpOnC4CSlFlbYDyAvmnPJzQw6nPyIvSWxOpw9SrwY3FYqwps
iNaKFU8DR7CTLlPr6CdO1JeJd1uOVaqhg3vVNDKQJpc8SkQxaYFi+hhrGJoPaf7iibFvi3UVKphP
Q9a0lsB5ArYiXFCHtBeG40LbW8rGj8IFCEAqtPPcOjULBuoFOuKg8omVoS38qp8dfliyA1Kxgta6
a/jgkG242wVGTrK4J6xkYbR4SJYFc4OLBwgT5O2OV5ysDRHpeXdFunHyA3eeD6l64OHzswXqK7vd
JA4dkYWK/SSvOgV3ORvCNOgES9l5//VM2Lynkfv1S1PUJfhGbxqVyLxY3l0SUZGADOE3OLclwLG2
GtXR89LdKW7aOmLtDztdbT04TQdxpqgQ/FR/Edh2oMcUPlegKe/BrRoTgHXUO9dgdYnuHdF+kN6o
GsB8f1wOs6wPdmoQ0u1NUZoJroA19Ir34vRqsXUmE4l4GuTXs611LdUp69eTZFCO3QdhG4NC/rVM
BJRYSdtSYkaQJMUqL8cjHfu7EgTOCxA01is11Yx6/9tXImi7qnCfvZLEXohOmRf1qwidDA6AGI5h
hW7enupU2yOMoPHwFF46M9pvTssb+iKpGzS2o0hGB7uqALJhJCUPnB2dL5q7cGvAIPQJgYCFxyyj
pr/J/dhL4Ji2zswgSaSXwhgVmqp15q+rui5iKg0nvV5uNlBO8Ds83JNQqDMg13mervkxoHUO7qX+
v0KkFX8DBWlQEjcNfgEpuw+rQHX6LiojnubHfoETb7tNfKPIGaj9/dW5cwomr5T4U7yWh9weJwN/
iTx+flRxQHA3OHjXRMhymU+ckss/Ml7cI5Scg39+uk34w2RVwW9F3HxxAGlu50RIm/xMkPj2p1iD
QVtBnBNzHDNEMlO/5gHNZChY0gpZLEB0jsnk26EmYLX1RIvGior5SghnBtk9Z0g5/QSM2EN0tHro
0aQZL1yJV9EIC2qEQqO41ntvC9362Hj8BMEoTx35m9TbUdd2HdIh8hJMqQHsXxJBUf/cf56aqjWR
iXb0zrOmpp8vlI+0iIh4Yr65JkevrNbtTz0hDRzl0XnymoCWUV5v2DohSUQVqK1U4AtensA95UUr
mvTzLNQ51Sd14psRlkl9MvLkIg40sYagphkB64HtzR9nCl1yNKTiiV904SZizDZ8282pzCl8rPbE
AgDp83YsmjcBy38cWhcOVxbT3W/s+02TeRk4ThWTysDHsPB0FMMrX51ecxSHMIsWn7Mls5Kf09C8
NpOOdAMjj0TerX/t8RwmFU6i+NP2fImmCym+kr2xAFpaBdI197w/aFn6V0DCSWDdifAmK6QPtxXi
3oLjfnP70n9kNSewytz0iAJChmgmPgZPK34KyUMLnT6xfJWVXteJLk+zqs/NEG8EWBQE89mUo3T6
pfau7PpKGAmIuEp1MbxK3rLY25t0F492UzV+Pk/I1dm2TYoHHiyTw4S/cfEuK5HSM7+S12py1qvD
+n44yUP0RJmK0hyAPyctnRWhTRWxL063TUUPcSw4SyicpprAJSX/Zp5G0LX2KXxpeRqD9Z26QCRW
KzG5Lygb9Onzj/LDJifvo5OMyxxLoWALOtSFBWvLThu7pOhHe2D2jc0eCCAOeuTcHGQO9gwyA5gG
M8EJaBQEf6kU9IMqjjzgmEl/4B9A4EGemWo5uqgNZeU/nWMJ/iHL8xRqY/4puateL0WmBQtEALsH
E5vUTlZgQItXcWntrAM1kN11yzWUUk89/ZOIp4p2oTnzLCNX/fudfRbXkQtPmTQa4WGlFSqnFzGn
N4C9pb19fy/T2YW3AUyofo1eVkBk1O/YCq2T8kDnZmEyWO1mKUMeEtlYHAIeZ2aQgWYtoev0XMis
MNXYlMc3IyzXcH3MBSf6sMkVoDccFwholdcMK5Fm7Ustrf1QU+fTncAiBETLU2s19KGBbdGCmQNv
kxVh6Ts19D6qhEMenXP4pkriknVdX4KYW9gXP+F1yStZ1pTZZtgxQ3kkxT9MaiUq7RKoCnJhjWLh
yIWiYPNLfow0N5DfaQqE8TprAetBF/tcyPtEX/aN7WDV4+/FcXrpayNRMuPJ9sUukfqqqdvAC2TL
+mLUm0OX7wChjKXpISkTZZblktkK/yzmsvRkCd2xypQHHvDcWnDg7V5fkcCV2v4O1KtGHwjr6eHG
EVC1f0bNRIufz2V6L3WtsnVaiLcq7/MSugI/Dqziu1/NGzcdQSs9m1ijXSX/gqTI8ULDpzDb2zA2
zyLu9YX+2EqVuLfVmUIeipKtgtyqU7if2VFRC4P8FJ/lxtvcCTo0gre+aToaUyUCwwwo9gMFEqhL
n5iKOfz7NkPZ2EYMnBCmJ+g7vxKofLy0NNNWvPeZ7L76smALXeytabKqDfu4EI3rCImXGu0lD7G8
fHRzQsX0pqFMCxPDR81OSmht7VhH0/VrjJeIA6xXl5Ular6/oESspQgRmxJFCE2LnzCy1rr8ANWh
IrRHgz3Rku5DCUZgJsBZjwzfELjmrDZmPX7Iy/Ew1omXVSvNXOC4UOABHWFUtQc164n4ktPUfYwZ
0VfxwZbFIcmqUOQI+47uw8irFH2xAbe1sf/T8AK1+HzfsKADVUlWVnEQxONtlGOR4zvN4460a/1C
N4YCNbcC8J36YPOtAT9G2LUyeKzEH3Sd+YYVSYW88EGiXBI8X2FUi6Vqzp5rHWPNzTF3eDl8pyqi
G/jH5iPLRAfjrr400CA0sRBa+zf0sWwWwAuiD753M8ppKd7NxtlBnmt2lRoGKEn11LPuwy8azuP5
FV+2kdOF4JR3uP7aVRkT8XDDlHhZrIQ0ipB78mFKoOq3bOmw03Di0daKwnYR5kiWqDThfQADJ9zc
vOn9Hh14qz2oxPPVbFHQlpAEmHsW2V4qmXEVjHMZUxYpTXaYkfo78npsBCl9By+cwDWEg3LYoB/b
XOC8SUEb9ETawipk5VE6K0CukAFj9yk2dB/CDjZN2E6U5+kbUjRxnm3vdqRTTwuc2kX78AYrB5yD
Yroah+3pUCwxyotGpoWXu56OKn6WKM3UX8sIvzcLjAWqAqBKoAfJAI3ZLqgXlVewQGmb+e4gGE5e
60PuUAiVPhvY2cDQX3K4COHfi9Rwow4FrIyhyAYYPvfkcEjQaPiNahiVS8BsQpEj6d6pf6PiFmlg
3lPxynLFDPU42xpXNz5AReJ1B0EQXx1uRCKvaH5W4j2H/mTOpwu5bIy6X6R/3LiUxaRkVvG3ujW2
53vqCDHlxn0O5pLUgPwxBGpCCVEu1MoRlas92wUL3oFrPX/0Y3lG/BKCWruifKjyHkNsznEoAySN
kEb/Lnj5ttG4tPYbrcABIIfppobkAJnKR2LbkRNfnqp5rKMOGjVlteV2A87lcO8CxTvgk87yCDrT
QARkvjK+JQMMcSI7UrJkggN+VuTK+gXvBuNrXWuDZmOCFkZCHFyfMBHRphgTYnXaQUYZPmAc3w6u
S2LlNs5Kbb/UkKZAImcWJ9zeFULb3Ehxw0nHWdqjrhD64i/YAMtAKzk4D6ewm14jpxSn/wBz9ePh
YUD3DAJbtnZYJIzd7xwjD1ak61yHSIh4H7GZDYDtrlM/TpUjyI7opCq4U8rjNjXvAkBTW5lGUAvE
mgfVzYIM9nPmcva90MS7Q9kPXM/kalrdPder6IvREGqNZC07FQs4Sij8UKCwUdRHNMkZsvAIPVAL
JUMZYougyAl5+XXKqZonMGEUTUsCXBKL92HVhaTrKMEGlVuqOVjoTDy5WZMyNl1IkCZxLSsUh7qu
9JLqWP+en5u/oY/pO2oj04Pciu6g6VwPqnWvZ1SHegIM/98sw+nCQLdPf3Vj2cvyafc4TtqjqxGj
BRICqWg4vWkryHu9QwWn4MGbQ0LHSz/u8kTFWYx2k3T72n6jmhonAMQdojENkthJ/4ezYj2uZN6I
YTVIx2zCiRtoIXnA3VEotKJuf7Kx4I45jRfdI2i+f3AyGpjFVFMJ832U/OYFotveuCqmt/tAzC/+
7WviY4SI1GiJN5ErNvzPQYFvO+9HWjH2hgiBBrmg0beJpMezR4l8q9MOHAVjZQKH4OuO+WYLwBVl
yrcOE27yhkGEdsSZUqZSy0J99daFBSwpDHQvD6xKGBd9NDfnp65YJOv7R0AtXSqo7+GR3e4HqHDU
un5jYc0m2C5p5LAfKERquMo5PLw/WVXCbETNN62Z/KzVLHoaf2ANRqIcF5LrXS3W2yi5jQynqmZ8
+I5Dlu5mb6V+7LThj9QrKM/oLxFrwzJUMnURV9tPL5Hb2hfTCtKeHngwVh8hEZIFDD0l+twF1D7h
dkqLLFT18s/vKQOdiRxEf1CzpCU5tzhiBTCdeoTkezTtRQxC7rnFFoOLdcqE2ePz5X6pBXRiu6Y+
LJ64V3SaBjBz2x2Pnt8LJJONE1GY2O0APmV3s/DqFKLIYuag6LbCNXB9K0mWUcpjLON5MUzIl0WG
uQu8Co8xAdkcopPdDetZd/pejWQvyNzcgvTW731lArqQt7TpGh/DQ9kveeQ0uvQzU/TDljzhJ9cg
i4vlJ4OQpqzy/pvLo1PpDhF+9nPpXo+YQEUCApf7jHK0aBD0wo0AdlTVu5MCgUFuD16X1p1un9CK
BHbGuRKlu3UU3OXKe3uBx81ithg38JzGQnN3jfJp1chK2Z7iu1xq+m7wl1pASgVU+QCqRJag2CqN
yFMZ+vq3SlKvB8ofqkHPfj/J8GSZCd8PkO2RnP5VHSpAg0k0NM+E2rad+EwCCk/5QgFi2n4i4nKn
iGd48eQDfel/ySlRJ5G8tVGM5a7ri44/HFW8d/7tCUeNnAsda4ThTZcjt3MFlGmNMSkHYXBB3ArJ
anenyWB4wTzCCS6yf/H6SS4bwf6E3n6F91YPaSt1tT7Dm8avZ8Vhc12OhZT7N4Rqs3Q59DcNL7cI
X8csSXQcNXeBQCRCekqTXxJv08wATI18pYABHyHFw+nI+Q4rUrvh6zgf+KQF9gC4WgR/W92qvkeM
7/yP7UZNq2pNLjXPAdqxoyIlEjxmI7APngjmWIq7XmLnkCARCrQ1O+7/zUxjvlr7+K2TYBHG0ssF
jUoClLPtm4HxuJJBMhxL+KSbG3XF8CzP5Jc2BudjpUtlv/cwQu9b3pDzAm9tUfWz080MEgazeh4v
Mhf+0LRYpP52xuXv+rQh7Z/EkSUoqY4iq2hiQr6KnxxbqSAjh3vIhuw/6N1yAGOe3AKKXka0v0V9
9kZu7SU7uf8w0s3p9XNfoRmqM/DvkkpbugQtRKsx/gKZfCIOf1FHrQg07HB0/lT1+iFIXpomMZaT
xmNzX2k4Plub9+2XhXmSI1aSjSk2HWeWBjfxNesE5ShyyiWE/OIqKmXzoEorUAawMbxaeLbCpaQJ
My8IUah+tG61KQ6/ENH8m7QED4S7RQGOYldU4dseL7mC4s+QxVjdoQGml1p8CtFsFVybtzdDnlQS
rJGnemX73x8hDjnnCUIGqQCrWctplJ7i7tf3wDjzFe7ndyjdzTZavVA8KougpPiUjsZjvJQeBQVK
uhe3QLZsYvnSmB8SjVi9iKKV/IHLy06g5HIvSBsDVfCecmdeHNmWwwnk+G2e06rX2SB546pIa2+D
hJ4gjNflxnqWYqfSGKx2e1G3tT3Uq/WpGJWSDJPsv+oyAzE8OI8d6XNHC2jCGVqmR62pRi6nkaEI
cb/LIsabwwyviZnSza/JMVNXSD6Y6o1RFd7IgIHLazTZHyEiPSvqLfAPn9FsCH8/cfzj3sHVBDeV
2Ft56zZf6SmMs8kw5J1bb4pm1QNups23t5DAfK4NULGERtzgXaWO0iA72fZ27Cjdm9XmTsLL8PDO
N8xCCE1yGBdXjFT/zVw0MYi/d0J4pabdK8s0B5N+qcLNyFhsE4JicT+C+/5IMPt6KThbtYHrhUvy
ZJC9czyvr+1c4xUKsdQ7Xpv7h2RcGIxx+DGqHBFudHvrK7wL3d+DAwir/6rcqAvoQnUzcSHJ411L
AJvnvUzj/mg9+sXxZnOdiaNb2RDyUpjwTnoADr5/jQ5gz3Sl6QNoSZOkBdHC/DE64Ka/yBDwSnL0
KwO+VLeDpG9wK4+Ivqdtvws7lypU0wMdhKKNX1YDgdJPVRpAD4BmZuI8rx6sEj5Hd4aNabDC1Vxz
nqJOPqLXuhZ2wHE0VBTtlHiF6L80oFIM4FPMn27pVWY7/OvAx7FxrI1DAxWQNVmDXcsseQobS8Sp
LY9nYaBCwk7YMdZ0UYjzHuB4r8Vy1tR5ujEmwvcBujBmTBxAf5tszxkWmWxBvnx8rV2NaehD23JC
LenqIlSu/qYtPXU4mS5WfuCAoB39dJR1FZw6DXJ+DxooiZPrwmepnUKr//D6XPekhkugGno+UC+y
b+3Dcp6kjLfEVU6KwRMPRm6PO+BM3B7RJxJg2ZamvdIFxPaJX3vmxeG4SgEPRIe5QSHOIrFZNqjt
PJ0rOjqNCGZZgb8A4W7u7d2PdDzhSMA27+cYTswHzQBLig8Hl3cOW9RWN2ZLDWNa1AlXJ7wuDHDv
Yqj4QzF6ySuHeeKqBQaUw7e1K37Y3oHoeBS/TJ00gC6jCHH220OIZ80ZKysEbInd0cdpQujuH/qV
f2GeFhz1IAJQhzkPbqoNbGuJ4whmUr7fYh2/yKqf9DZsmWTrc7M6PPLmbJVmedthuJvNX4AW7gKW
uFQ2xcCzg8uHAyn+RxdGgxspHIR4Kzet/0CT7gFcvrgBGTSxIM+s5/UeCLAXO/DynCHSJoIvmQae
x5hqarx/wlp4ZlZTUW3czVK7ShkYcB6pQyC+iHCyeDxeDiekXiY1GACbeEzzNThby6oqpScsGir0
Qynr1cgRUnmWK4igHaEVGte7Dih3w8gJPay2fuMEK0rOTy+k6z1uaYNLaHBRLWUrR3lVI7VEJUGh
7mhuuJCIkYuZbreMxj9zzu+749aOaAMAAfrD73eaUTUN75BK0y23pauEG+sR83W5RAqg2nBv0U11
cg457N8N8JlwmG8lfxavI47G5ptUSmQClJChFqG4Ii1vLgpd7u2xsIPHRgWZ74FbDSDe6Ak4XKyg
J+bgx+8yiDJW93ozZZj8WkYAEc/22hYd9pgo9ncB5A/rgUWQOEwsvIyjmfrQoz8Xt3MlzEPqvrkD
nasYSXMG0tlpBZOciIq5masyXDHyFu8Dm8pysFNb2Z3hDTxAGDoE8leVdxST1tIhqnBi+IGRcCHa
ZJiDQxuktc676ct5O/JmiBF9WNCjCtufmOBncDA0wOLr2pogfiXccHBGmzWcBCDho4nFXuMkxW11
EnHl6Z6COnsFz8qao7PKSeIo8i80oQHSJa3IjJDsWjJSncqV4w9RwHx6LMCtY4PU4XsPG45CRE5W
bRzPqfBf+xHn35Nzpxg47M9VPjFVdBGdrajbTAE9Nvp5NAhMYKFQUpVSnsAaTE9JQInK1kX1YIDB
4/+2sWlUAc3RzEECEaMlIecpS1p0irpU5N2scuvpxvQTAKvkD5Hw0ILu6huqs4uiwYYGr5QaWjBq
72TiiC7yKJOohvi9a9120I+wKeCI6mY8RItE2csoVMevVjPBLWKatu7WQc41js63cbzrgbacndie
2zucGOZ39q30AbmaaXV0keaL50NBBY22kowPhlxnVXUi976lzjQ0C7zwCvbgaWVg6R5kneb9P4YT
rCymaqL63rsLBDbdeuJo4DWSNH9qdsBRSUBJHuAE2M+LJ5FBq/vuuacZJdXkMdjUTgrBsnNfnac/
0NYN5aaMBV7dO9T7GoMECCYiB7fqUjZItCfDQEZpSS+b4HV0xPgwFFWchaKIV8HCVeJE6moIoyb1
u/DawC43cEeRT56k2jBZgdU7v5n4oMzO11tFIrP/JlWXOYEPzfXk6yI07W3a9FmdfaJ0nRJiHJKF
VnbeypdaV+JH09Zm8FGbSQe4L4QJyRlDE30uqm8QebdywAKcSHbMLIDB69Ca8IOymF+IKgrDuKEJ
eumLd0Ri9W/04bbmzgSo4crhCThpWVLNuHwvcav319Cz90+jV1PztNLsA//jO3WYkGf4LSRA2cPC
4UDQeRhxvfMscQXhWvl47VOKsqyK2MFvcfEfIf/7ESEU/L6wSzV9rI+E3m1/eMap2VDoDN6rjZ1C
g6JWUqZzjvhXhX3Fi6iwxKogYKat6UVpO9ZGwt7yrZp8UIU7HgbhowtCjmzBFJ0CUCoBNQFfp2kq
V427mm+ZIFvT3z/YLHPnrIbN6irujl5qaUBoaS1ZohfPS8t7yeQLJfexII2w6VIqsDSJYVgjKNQW
/cfb8FEXS2JI05v5DFBKOohQzo8cvKLjoMAkapznypbxqkIXiQkoliNR9DpSpG/akAHDhf7nhk1+
RiXmzaEXlwKHmAoZrysEPJcjFpyc1c+el3fROpCO/PtZKfH5KEg3XVXG16YR4lP23Cm0KT46f8Z5
PlkU6Mx83HY94KKVWxZG3X9ZFHn43e1dRgErXsa/S36DI2vft36lajpvE216lKV3YgbBdG2JDknL
4hRxZUTzI8KHKrNWGY6c32gx16K3PEL8HQ36F5PDgzwrP+8MBXF90lhI6f9pU//leiw19DZ+vSuS
4Mp3SHjV5GxKmP5SYqgmz2JGipxgOJwnJI2gulhuwHhtwINZAM1Sjm37j7JEJoNVaRjtQNd57cGW
5LTR2IsG+TRQ+iPaF5jFK+XyjrETxH3TTypjqIUG1VMscF/JctuMnbcLIZxJ1G9lMslX49skGJir
Bei7wVg0lmNJ+UXWhi6+yRGWjLRHsRC7CtQUq3GHVTwctbGJwy3bNcR2V2uxksIeqGnBgZiXoVVn
97ZqtC4GVChlWb5idEb3dGzvHcjH1wjPxS++ckKDH516ppjkcJTW55AF1jxp1oHnx4HhPKrLjZ8s
qv+oxKoCETYC7sr66yooFIUmXgMV5MrCJvVm+Vv/oadSLcp1qNqAjaaSBtkZLB/vDU94zE/bG4A+
wWhpH+dVh3fqTEQchF79gpKsx0k4va7VEc5DrUg/4+hy/4HGhe7V7iocLEsWzoiF8mYEqaXZw7/d
tgXbFcPOzDAh1NajqllNYsOHg7a4GgtrdkrmNYNtkJT0ONrLKmJVKOrTcD9XcYsHHCsSQSSZJjpk
yODZnNxQoQXCdLrWlai19lfzwCUG61U5ixfNW62Gk27CQSRYumV76Im9EcRV9OesqlOgwGOzmWfx
k1rP+oPNy40hqlZj1BcG3rv8VxkphCwC8JX5IA1IU3am7lIPbO4d0lr9DkjuFutClCpPTt8lqb2w
tqGx/r/FerRZrmU10h/lFvs23f0J9seLOznMk/bg2hq1Cs7IqiI4TKKb9NuW2tt1gF/ZkUqzBOmZ
98BuLqNSUmu48DG6njnoKvF/56uW6NTbZ4PYzOwaRlnLt1bX/n1iW5bt6Pnd15ksK9xbYrvaj1Q4
EKiOFu0z/QvRBpMDnl/Q2BfjRuahcfK6N++UMB5phXaT9Kd5UM77Vl+PxR+fZTHftG+0cmxefDqJ
VuAJFnoSQYwQLsa4f2dAoVoqf+u5oEXL1YFvnVBdmGcv6ac4oECMqL7V/X6mWNuY/V2MDquL6vN1
qZlHIP/N9P9ZBbRLLq9WKpKbLM65JqGw+/+Jbmn69xlAipLc9fchba4xS7x/uCVkAaqpSQdNCiIo
ddemvgyJh3ugX3UzGB/fshjUWltw9UPqylFBaqgfjEHSQQe7d7A5sOZOW7itLhI/Pt1GR1Vpy28K
VC4hbD5AiuUAh8k+aGjIlCK3ypyVjTjQDkX7XqMDVz1VcCR+dcXP7nolPLHzuAeo4SaTb/ssISXL
hD6NKG3pls1BQWwgenTj6990FpuYQ3jjELE7pfeuXgdbCATlhhY+t8OV0Yknl0jcdCreEO8C3vHl
y/DiMP3zlKZfIZ940eo9BsLXN2W0XkW4Yxc8VqtjckQ8D5Mokl3s2SyubJmG5uEbraGDXr27sTrE
dO5npY/HW3lnAb4BRJXk9o1JEBC0fQoKcjogDxYO5hMEAcE/vs/O1YQRYQNIpe/gMwjbFn0+sXMm
QBzw8daJsevc7Ohrr3wO7R9laR4/fl6R0VdPbY2vLGU4gF4sN/3n01aBBnpBK9MDXX1yJ1xNnU5k
slKJPKbGpxN0DLFNKmTqD94KQ+iq0VeFJ57Vhd+yXmoVVrBgkcTqcgjQMbiTT/ngb4Dq4vF8wjjo
eNyd51FTMakkKIzaHJSEW1u2J8oAIIC4DLPCcYpmyhoK/E5E8H/UTRsOHP484nUXnHwVMjjkYqbp
NPM1Xw512Ehqs2ve4ekT4IGkf6opkM1GAycvn58GNLVFdFc+jNCn8VnemxSvdMdDxfsDgF4xYv1M
z69iiOkdxkZ1GB50NScpLbOnhm7rxT4tudJz4SxNHf7ELDMfI/fmCWCj2tfvu3LIFzTp1YmkHmye
mAFT/cqSi06v3Sk4ivs4ZsWjGrbLOyDei204MJd44ReGP8rzoHzwzHsD95+zMEFIA3smw4BUOo7J
ktfHb/Y9+NDpwWYBeIeh+mejrXS/62oR5LPkkoGUO9EyNm+R8tioB18YBQSL1D1EOsa/VjTxB8LC
wpGhwLou0PT1M6mkoywXE4t8Eyx25cEZVdPA5jtxtJrUIzeD4GroxzSp60ZT5Qsywn3dXgbtH/+G
yiyE88lI149WZF7QN4EWal3RVNR6lJdkJDvneXFr6Wwjke/XXCscc/NG14P2K/YxujpU9iA1heve
SCNat5cJmx8hFZMqxUO+fGgEt3/8q8ZMjbDbHTwNj7uPa8zwpZubCVX4JKqoJhRjfPQI3TZJzmjB
ThRpqtvV3zA3DRNtQzcMazfed7L/0nXjNTNreH32+571D8gTraz0CyqHBF5EKReik4/bXb1hCC/1
tJ76ZvMHxrdIgUrrZdE7TA/1qZguvG3p/QP6C5JfxGAWaqt+aIMJN2L4/v8d7GblVVw4YD8y4B3a
qJx/SZ/MqC7+l5P7VQVNVsvTHKN/4NZGREvvx+VTckrlI2GlyGAkLH5lNu8fn5Z/g0OJXcCvAvHF
MTX9ox2cjBh55XzHVH7uSLK22qYZRsQFfJ/zswtWI4WjiJtdQkFY1JVkjXg8AEAxcW6iadBxShVm
f1kD6JRaJt2mba2CYL+diy3LBLyFXGf8YDB93h0HWaCIslGESjaAMcIkSqsYn6pexizkrB5Jj2NX
S2D3btpjrHtWLKOQkt9SClo37Zr4cp5l/WCr5J6/PMxGEHp5f7DvBgsWw+hzYM1Km/r+ov4urVYu
DYFmOy/rs03ryD5aebE8+uNIXEu0ITeqhTVVxvVuo+dGNpmJ5b1zOT8LrHMw4Vf/fBL3FhEAumbl
kwmnLLhHKwST+dpvKuWGtPdKkcOrmhIo9sJ/Ii0acOwomxnG59EMailPv/2K5YBDlnjKH+A5zyM+
WXts/TzqznRZwzoCS831GURXO2vQ0dInxuW/nbfkcMpmaB/6DP8HRdcK3Tair3ANKG8zsG8JJuDt
f6rrCHcHUeXxd7IfRJSYb4j+iiX9fh0nbUa59zUdqef2PsS5ac1QJ2IQUcAXfo7JN6tDP5Q5XVu5
EmhtV10KbxMtzffQqZe+Bv4t1e7w0KKNaAfs9vfRx1Z+k6hjl6ZAkfm0WZcS6f4g7gDJIhV2UQa9
MfiAEMpS/xc3XZh4xieGfdjKGcCRve1Xcf04vZMSmV2o5rX8/Auf2/mCaYr5Ez1m5k+KGeoYuNrj
HP7PVu2wWYF7H3gxqUdP9mKcS3FAunrurkjwQS+VhEnnYk19mAJltCYV7jSnmKdhZ89S4O2WAKzR
3P98fvdri9Sigl/1w/AyC1A7qn6fksfifysETETwvt/NMyZzs8xAntq/T+pi5S1USXJKMag8OLGm
ngTWd1V13jP23vIQ/9wTbsDr4UH0rOihGruGrja4PwGiVRlkhtIeMf2R7yfuanQ5wL2de8ZRipEu
Xx19ux5BAXu6413m8w/CjK0M+9ADR3LqPXlVVt4Og9EBgdI0SOs3g/FuCEaWKhYZ62+Fz76Sv6t1
6qu2bJAwVhoNBlfzzRV1NRBQ6tMUC3V0sXCbA62JSrSQUylwDo00TwALAaRvYGwkaNLHCda7PmIp
MqeIP6cYg5Aynf8sIPkzvH+w9J7N26f6LFznbfDYbgYWiTAWKvGvd4O7wPFicQfSkBEajkfZrasU
yVUqMbxNciqEHpPBBVhOSkQMasSfhUfDReOxGP/d/+gxZfeRWxj/9iYYO9NQpd/8uyJpb15p6je0
wHK0uHzfEdJFcchj/EsGvPtBHgrjlSSPwyeiQJOFEwvXX+yQSKXKi/S0UMEjc+sbBgrqT5sBtykV
qHpxNkCk95T8Ud9Tck+cushQTtyR8TOUVcP6VKG4mGGFHqmcsX/rNxfbQtSNgfwHlQkFgR1fC+d5
d6p5Z+10lsBEdK/oipvcsiFeTBTVjwi0CY55jThkFloVXVN5NTqiCowH8dWc1dWKeJd7NX8vt1U/
ztFSOrHa7qF+iYQBRltHKzIH5C7MJovrgJcQkNgO0eW0ASL5mvEoPTFdS7cctmB6FUFaVQurUTQw
+lMcCxqcVluw1cawbmicOX2KYY2fZ42xU4DPEVKQ7RwK8VaYl4mwQ+HdgGg/isT8hW++1kgfCj7U
a7OhKhPFRH9gYlpxvhdimoqhGIpdX3KEUZPVp3s8MBD7/Aw7NtDJQoDHlFCBMQxzRYSjcPaNDHSH
6E5tCzP1qHQJwKDsuvo5Quyaf59k3xy8l6NbbOe8WSje8ojGb7pyf0B8PKeUXkSdYDs789TJihZv
5vzUqJdJBpm4/MpMkRFTrtmwss6zYEj85y67BYfVDnjqXVPJj3OmTDNEjtwRWCHKyH/Apf76Cws3
U4BWPVZreszFyTG6k6uJoFnb9DunGZkAnYxZGdDguE05hfxv1v7DNCU91qiF4uOqlczfkrkXByaZ
THSKq9O2LazncAD98zKJGO6TW8mNjDOpZ4fYF54Y+Lv/ncfqdJm+OGy3fGb8ahkQ5ER68kYQQ4PL
9p8fCm+Txbh/CJsaiqC5Ywpdj5g3iXyWo9tLnyPuWXeMxaChhJ2lgAZpXjRX7jHiojJAprv/ihJN
0hvghytG8zdDV8Nd2DKXxqRoYcUWunRtWUD1c0XFfvvMbOWlcZ9SaCKaoYVGZBVMLUxoca8yJJr7
hooB3xvTdxJGQJlB+sCnyjpHrD0YJB+MBkLeEvfw4HLr2teTFQ/NE4tJcv5P4l0HrPmysYCrkZow
+QpCR6ga9iKzvHyScGvvej6gfEYaqYC5WJjB1PSj5B6P/s1tPA94L/wO9xxUxrJp/0wkzjp/3UQE
x0pvTr4ACBPtIfZvFDOtWDrveR57uR/+tfhtjZruGuqfqbbN1ZllUNbZE1tVZyy7GQgQTBtR8lQB
IbLLE30h5KDfYIjcNs9WpQl/oAann0Z0704zNCMMPNxzpVi5Bluq9dTbgMKp6JQWfQmCYBj3Ku0r
pc6py8B3lwo6eXn06n33f0FVxPGN4HA3pqJakJUeRg+0C0j4dWfRsVobrI9ukScuMwMO/emqO6Zx
ADbGrQNnuJWClTQV3hISbgF4WQOP0Mg0RQqSmkTIkNZ0YzHn+sL5Bp6UGTEKlyGS22WjDzC6r3Bw
EJQwpSjrhaxSnBFjdS9RaXIAQ5iQPUy7mnlbzapaisu/J/SKdq0yTTnnSIbEdrAjrJZTJ5boet3F
Y7E+eKhMR6lQtz6k0oS47gYrCe+mBOSciY2eyurtNZoEznOJnis/gOJabKtl2YuO9WZhEf3JJCiE
+4r+2J1APzB3QmNXH/EAQ5EvCXLL715potJg/y1cFVXWTWsdjVzTDl2F493DPbnhHzZunQxE/IHh
8H4Zc47S0joJ76g99cAFrJN/CGMTGCFWANO47ClXkhi+/5bv8YW0izMGTRgWuApIB7XlrC364kdl
JZo1Yq+fPCkJq8y/tBe5GkUGhTV5FPI+wY3ZnlhL5/j2IJtFctpkiPk5rmo6pD9Fl7JNy21pyrzO
n0rUizDjVv2AC6oA6KDDXZ0BrCCibH3c8RMpGn2CHHEyLEfjZxEOnHwNHOzqq41d0chUdKs3+sIC
FaxfpW7Mjd5hRDEjDAbn2OPFhOM8Lc7t+Ofzu9CHVzSzKevUL2cBoqlqaKdHExbCHHT1E94oWOjh
/pFZXqucxOGEYjfCwMTDHK/5awmA27nHh4Z7RSxcKOEHJwJ7VE0dBLe8SYdEtbMwGPwYflhLmGmD
5PBYC8EHWezz8nXWv5iDQVp1MYeex8m6Inze4RfkiGNAbthgxm3JNy2xU/uots/87CLcoliAlBTO
PYgy29/y4Rti8CL8owQxQSyFj2anwnii8AiIDi+V+2BZbFRT3jo0RL/1sgx8RpXPv+m2t9eo9GYR
zFmToyM6/7j25NdNCi3M2nTE/cjXzDjNRtHmkk1MPV56SEO7EvuwyMPdRrXNmTaIvXTdBK8DkwhI
t/VvJ4NMB6gIUgOWvb8Jb1akDH99a32NKvvKuuQSLn4smDYn4JAIvVoC3RxEVBo+TOCNJkFLDBcI
dW4LA/YOxca1RXe6y8SMinRn5dcJhxzeXVNWNOgjl6eKXvQJ3PVJMEJSj921H35XEqABwrpIFDcJ
/Tz96U1rkmIvmE+RA3Tt8w5jPQhH1bzPlWvw0LJPGhQaSc05WFZQSs2R2KKdIw3odpNg7kI/w5lL
sdXy2ZIO7bA7Wa3qQHM+3ts9Itm8dyjF5wGCBN+g70uXSrMYIK3CyAQlvsKUvEk44JvdgyZw4nUc
mMnH1lsZKk8JjwIrzi/nVrGBMF8m5HyNlH765G3opmj9JEU9dWUwGxmljLIc/q04jcbZ3bgiSATv
fGNiXcJtJ+Voh+6dtarw6PYGNRZVL4Uofoa29gE4hu5OAmGgdPjCrBQ/ZOreydGlhGDJgS0ixPCm
5UegURFnB2N2Qbfr9Fd75ZeBQcQ4MgJf4AzI7srCwo5n8cpUFYBhNCvoakaJ6B1dUk37xUpbKeb7
FzxIIgczlrW/SqkuVxjgbtbgC01CEDWpXdSEcukqFsx+xl333Rmn+UcLSAB9+5+KsYAI50VhIdgv
D3lsSAycjtnTVeIG192yBx7IoQRl+a8P0Wdd9tVrQix8PtfYBapT30xvDqATQta9vgSr3zYFr5Wy
pH5VY/w6QiacGgXVWL0lCaxZ6kBMBPhi1gQPhsKFajwS0DnsyMVGKhkNP15n2dj3QQXHIWn0LXuD
AjSJWBxXwgFOxZLKu34xmuPs41vaNpzAEQG66L2bCUa1NMYRsjn36SXLb/WAYtIHomVWVavuQX5z
I54tUknve03u5pQ9Nv4pm22ykldvaHb0cb+7h1uEdntrsUlnuH57elMU26ypFT+H4poOYYizttqA
EKl/q87irDpC4XHOHDAJ/3wOwFBnbnnEoqcXPta80y/jGDG+5dRt4MNxyrCCyMJ3wARSWJ/B1RRe
/vXu7WDVijU2BPnCLajrxjXvgPIKzFcQReobxM323UlIHl7vK9P3oOq+3h9Nag6J+ULJuHrrIJYM
x4GgSo+lEvPxKHNm3AmpnerNN4CvhtdZsfBTxzwQeyl83JNFGOpkSZPtidg0WyM6p0SNyKjZqy2Z
5o8+Jcalmmm14vobZdRcbiPe+46vhuqS9f6GTuStzhgFVZ+AC4gpuSZRTG/RQHcpQyacDq7k190T
p4a9OIUC2hzZnq5koe9FPUWh9sb2A05I8Vv1pGiPIwPEt4E18dfjuf4D1434SwUp4OyvEVDhdEzp
Ui1zAZjJHRywoXA/Q9p84Pmec/K+D/AIajogI1pqo9M0N2OcW/ciqkLErgZ/NvfrT7QT5QzUmbPg
xM7dm129c5NXAJgP62/RQD/HuZ4HvPc3sLq3Mri5OmJSnmhg/M3ZLkyPEDLdDZN4Kt83YYFtyvI6
KvKpdkOkXwQPndB5d5YlUrjV27svl3wj/Tz1CCgbQpq/0svLOQnRBMsZ4+0zy0LUnn5iSluQjZEr
rdpic93xhbgj21MAb5NKHLoAvXFtlyyP35AeKbr1u0yt9vQrZ9+8JJzoniiq6jxvyGm6AASAzj6e
rzJN1F3pJwqow6KroxgqC6hoc+FBlozK1cN3It3mKlGhKudbnYbaej15tXqsT7FPn/4Sfhv9p3mL
6lvUsGbdBL2Mvg/xqe/Fyl8Q9KzMwmbaeUZqvsjQ70L7H8ZWyLJvUGsu0EXcvPofY6EryzWq5/ni
u5TmfWZ9W8luwH9Q8xlXL6n8yHHRovyGsIaB4F0PVjOktJvl/lIADc3IFER/UVOne/XAHRZKWkMT
Pf2l5mPto/6GpPOqZuc857LjEMJ33OJyuaZ1m3pulh6ROPcFULGDV2MdUvJ4nkXZaXzEYpNr8GUt
1e/+bC2fs5dwj+/g/Mnz/3xLxG18o6vSEJM80IJpCzKVV4OveoMAGfY3N5wegN/EZtOUn+BCKvS8
9tKmopTdW6vuO5y4Kq4qMqToVSJiPjLikntbnOM6GgWZLFLARyy5SY8x1iOwedbIEzKeTjVfb+aX
B3vxbZPRgx7Lwtq3NRoPdxv6qipKFS/2Pg75GdqXXFNtJSnXAiNgdq9mc9zOTXLp1k8FoitLkUUy
CcHPIVBNyEAliVCEdnKVoOkvUCfBB2d4d6Y8pAKk44oKarEtV85riUBOcryvi7GTNFmhp2GmYhRV
BBq3JxfzpkMV5Jd25vu/FyVTEEU0k5OtQw7Np4FY19XDdl5SHFivugqWjgzJkEQhWpngNztfrHMa
7f/yM7pRTw7UBo4ipFyZZm8tNDPR+sKJjM6vED/HToxkSs/BWidNs1Fn1bJa9QXaScf9MKwj35wz
sNOzDb+Aq6iBkqRpVC+WRhFgRvhckX+we901NZ0OYCwcH26PQfuw2iMFSW4d3+Zh0V0a4zimG28N
nwo11A4q6vLG3mZOHUohE3QkFJd69toTzOnqdR/nIyBL5vPVQNxS0O2u2lq41PRFsNPuYW9aY3XW
tR8Izjl1AsXOYUKTqsuIzoSdQqfQFjqtDwCqM0dyqu+o09UAC4/ILgZ8UJ8CgRRqJ9XK6QAgEyk0
izMtLw2Fci2qaiUQIhI0N2EUmXFRyXk1vvfb9IoxzAADPBVyVa8ed/tPGspa6gYC8Wtk6Di8h2Re
KBMj1Bq6WyD6MiysjkME4fg8hQqjjFeWC2BJlEwRE7kYai/4RLLVCjqTA27SI5aq1mDIT2mCjRXX
vBI4cmDKpHSOTyQqWiTL97T4uhMiTHDdS4PwXnbq5ZOY5XgvCRtSOhQBT0QSLFJLckpWYtPcddpo
8J1dHKYRrAzpND7qafngWHqa3wMTo5AcRubRhF3V4jYnx3cQln5+u9en7JlquPtipGaNuYusaIgL
jqiz3S4X2F55M6L99l9+GFJmuCZeefs+Xtze1qodd44AAyjSp6WusOGKfTsx5S3OeuggwGpwk2iJ
tQ7s7EVoTxyt46DxGWRHXA1Oy+NigCoCPF65Dh5oKu8hgwexb3xmvJKg8/+pripm5xfe9D9iUe16
fTwgwrFFwwqGKlL0HzfjYdQnfgjvWqP7WZQQ01XLIA/5Mf4/Cdt28y1K/MALSPTqo1C7jAKkqdN0
yzz1kQxmGaEzOFoOgdP2o2Pyv/WcXZxqVSifV4YUm2fPyTezPn1nU343+DskJ8RHRCRSGE3m9MF4
ZKUJLacjNq3+XuyqZkbtEzpaFtBDdM5/Qwb5uUHgf0XJso1bBjGSlRAq68khJ1jJYOX8FFia78aO
k2cMA6lKdJXR2xWkZhfw/uoEbU8OkU1tiH+BtmCNJvNnj5B3XOAjVZRtE9EnZRaOjJ+4L+Fu0nln
3t0UsswCiPR+zEG1SpIZLhsoddx1tgMGpiXTv7qy9BAx5I+8xcU2+9oUtGV0ARwFPxNIli3VZSVn
PMHMQPz0Zks8NWyWJpHXjX+BfCVSPiHo5H0lTbuEr9rBVP5foHa8g6rQj3qwnnvcPygcc5+3M3dt
mcRvxJAVEm83nMd9PxiK4VQDJ2TCtHnXCNfnRim1IfPMUL9cCFN7bffzPNktVEWsQ5EzKFSfkFq/
8e7+DfZ3LoOs1+O+Rd1l6+WFPcxN/+XJNVlUvwynrmr0wL21oRA4AVECZ8WbqC72TgiuRqhik4fL
Ih68A6qleJqdA2LCnMTfrLbJRfKTEZT2LqTsCSIT5jEHaaK3r0T8Moz8HK14zWkNV54cxtTK1N4p
ZWlllHAlWVnyPsoNPOfsiZK/UVmQjiLAr5uMpurok26vq/wa+640P9R+RlTBnlDza5tAzO3n3bFo
eUWJUMEuu6FrxUpqHfJHO31SHVlXwXzbJnrlWI7PAWAmsdWaSWlqie54t0+nb30CKAgbaPyUDB+y
EMDMaPxTC1tA7vuSeP6Espblf1NtS3Xrz+iy6AL9rikT7O+EuVlFrsa2ONoxzJM7uq7srkzUSObh
3rj87uPH+jzW8TJjU5f5uh64EDRF/KuyIt9uB4ZgOnh+iDXL2sNmAH3POVTy3yWzWJi3Axcu1gRc
YzC2XVj6bxkGL4HogzUdLCZElY96mycpcrkDnbC3o/UZ/ohbVegUgHO5Bpt8rpcdWxsU65d2dke7
3ZSp90t06veE8XGogOpbPrgBV/L0ymUZlRUL60SNu2t00RigUKqBm+ZIJrg9fjAvVZbDGcoGGSxj
XNkpaJg4cz7/LFmihO/eLH4aX8DFQ48CC4jcZhvQTW15H3LtLYMiAFzHLHX6F0jvcXn6wmtM2h7J
zLE+ZmBBm2TmgAyilPdyOfjtooIkHdvcHcduozcRtS3VQVrodSFoQ4OMTpeyCgv9wa/fCDKDX7q4
G1/ixpT7gaDa2ABVQmRbdwA1b5K9FKZ9RwKZhPP0hniGumC3WgCrEPrxb3Lz9xqZYkvf6W8xcWoj
8BGVbhk78CDdm4Pwdy3kmJkUj1CwVTM68UQJnbCA78rDUnHB2IuJ572vMbSjEvhU1mqp7mrAQZNz
nOa75q6aAP3py11valURE/BFYvYiRmYvp6Z9nPaEid4Bn1rIXvCkKRF6Jv/ahor3pJMm8h5Ydcal
NQjzIxjl5c1uNywpevwRYDFgnAZwSUuaGMM0dtkpMPuRPmae4XB32/Zl3+XXnsEzhDxJnq2cwzWs
MwIYT4KNPEybyeuk8BpUtGsOsPgrbJ13qIgvClCYbD6+2lzp0CKR+czw0/v2R+ODphyxmu5ncIQQ
VFE2DjRnS5hCBQMEZCiR3tHVlkHi7b9EcEX/Zq7MUgbNG8F/SUvkply0uV1CwYPRSA0dv3fXc4yY
jCRFpk/hVZ4R1Uhy39AKRIrotRy5IoCZ6LbKgwmzT1Sof5VNRn2tjIpI9VSLwvdEkqABD56arkRR
x3e6ZRUTO/JvHFs8KcrhfFmDtIBHxm1vGkAvHlBWcrSZNNnWsR00uzEs0hJbasvV539DCcW2XmLJ
7K7bA7QQbKUuUPdQ8t4Z8JcT4zFV46r2CRi39YQ+NMBXo4elHY2TJkF42G4QuGHobBWrjCSQY4gf
jTlwBb4zXUhYO4I3L4zvRMUOn3cxj5fafE8jUz9du5L+zMCizsSdpazof9SxxbXcf031L0f+r0FI
WtlNcFEMFI2B/UncexlVLsb09ZmAHP+t6s+dMs+SvcLsG3mZYaGZYoKio/6iJ99wTWML/lT8Qfwo
P2iGXjKh9gtm2xMGhFyR1HsEfyORW5JK29r39kPsFiCpoTmSPs5vJryvXqdCSsUGADLIZRd+5hZa
4Hbz/IiXu/PLJWLeQuC78tC7cTVhQvki+EoDJ2UoVYb8Ty+CSTvWVQkzuU+7jQD7fpaC5buqHxVn
VwhEGvtte1c0iX0xzhmRP5XbyFaHDOIl7HeulIR/P98SzrcJxnPLPAGmN8b2cUSwwkM+GlXLHaZD
p6JH3i+j2bbyXG4K+S2UDv4hDUjpUApyUmg2rFsGnVjYqtcfLtycoyoTRMb3ykXJLqj4fV2e9LbL
3bRtX3endTRwojyesaAuSU50p/YtpDy6Qow9hWFlhUaj3Vo10FR9ER1W3Dd+xJrQ3ChttwEMPafS
YcLw9J7ThreAWvndXn6RjoAB+W0XousFL47muSTijpC6tVX8OdD4rbBzHjK5C3TKepnI1/fdlnlz
UKyWHK8fWoFanRf0DQphiJeif3DbKZGEH6GhGbV+PHh12vKTzjM8dZxBC20OQCNCf/uzhnPYAcMD
fqJwNO/ETTua9ytk75UUbD/UfuTrGpMMA3zpF61U8Jfv7kjMK29Lb9se04CZQPbtotZOCSnZEfre
HF0jxOyNMWh4k2Pxw1mcI8xO1LQNUk3JRZ69lTw9dcYWiAsVyDep1LaUYWfxJNy0VrnW/sut5i6Z
lG6KfzQtTXqTNfMCQlSmu1TiNzqU/MO2Jcg+jErUCcwZsSyJITnC4YZ17ZmeCzFFcsmqp23YW29v
fB2xKOttAaK2TBHQFqRrjLM9imxRifC4HKfO6sDhEaWfKyv1Re+DyF3r1ISNauSIwZmTJIE5CNTn
663hkD6rW+yxMgmxvqiEUmCX27QBBNJSKAPKoq3p9zOZRC1BHXoL6BCl9WR38izWEHaAXusMIE1p
Oc1WBCc7mZk16120WGYQaN1zz5FP9gFGwrnnUtZOLM7iKTE92xF6oC6OGiQmOSEYz8NRo9SFoD0k
XP24KHR3iSwhWJNwdayPmrZCxuNBFnoSnqbA8XHZxbyjqCmFFxZRrnqCem9mPFzEIJ2xW04aYuM3
3Z47B5lKqDDIPVpPs2vzD19jkDJSWPffNYjFZsGl/HN0UdZHiG+oq0TdrF3Qo40PMCNuplCA/Viv
0yPpP+Y7RhIc42JocZlwlk3DfPmHA2xErw/glWebUlHn4rJIYPbTMNJgDNlydlqIXT94AUn+8PT+
U9RC0lBYBgIUOr3Hls1l4ep8lCHvCVxDH0bxNhS9BlMqQ0b7VF3S/bAOvVTh2V35SMpYE4+90h7P
AgyAnhUmS2hVpoGZOWte2y5C8OYq+3dojUgCWTifNnOeX1gNZr0VZHy8PpfGNHgIH3k6uPyT9VQY
dCS9Idf38HaP/mLowIDxSXRUnycQ9sNdx/iZytJqgRuALtC3vW89GNtaq9oQLgzIrcfYA+PL9/xs
lPUwGyYgHPsrTSymQsxcOq4CeYT+jxTwlLi2OBuW9sDHmJ/PWCaIMRwmFm+47RDLQd7vmaOiarTK
UEkmDgKoSR56cg7/8O8MHEM3Z08gyZTVKFWwXR+xlLez5vuNix7M8RSL0OFVn1ELY+ja3ZrEtOx1
WmvWoRyj1LLmgxKEbAQmNKCsAvF7zKbl/m4pwk1MkhWRblwoKjduRaZbp8I1/G06okfqHaPiAmNI
qtN9kIN7AmrrqipRw2WLgPtv7dL0LgL/pvz00jS0KvhdWp+af16wMzRKEl4kXjeMWr+ri1sC3IQ7
WtnH+RqZSY1JL95bsUrAuY2+qrCDkcOFGng9zlb9cNBVXynzug3sBn73YGCZDMo95pGOpG+mIizQ
MS+kzzWswkm9EEl63WitgIUrDgnYavJdlWFiJXlPXgdB2fypeMiR/9iRX+1jOsUOhQ3/tPI6YfHe
zS8yYtIuayN4+BqOsm1yrl0vuRhy32RCtwyZ0g1FOGgnNivG3ObW/hwrcJVhFKftu/iiLOixYm1k
lNmMPPUjm+puPoHhxcZHd6i9jqg5djVMERXdfWDEbaNmKsIvERqObR7THDu+WcjbQEgR+HSQjdcz
XWTlSjsdHUAN8XL+HULMYpDNt5GHv6JMbwhZDHP0WWiepXZ0DpbBtQt3+8PLhIDLC2R1t9W/p8dd
Y5Eierv30sqpCMf8OqUcOa0MwojsmasILfvx+vxopOLAaqvVE5wTryDu5LOM+biXApDChx7iPHXF
HalwZ0ygU5MTDkmjRl+U2KRdJRl+tYjix4hIeCubswuaqCSUZYQl8rP7pwL55n9Ti9MMjxViVW6R
3o8D4WNsD9WrpRouc2N1jjn071fBmL3PRCWuljq8HqRJb0B/IYN80shpsBr048rMBRScSu7f4G8r
uI7vS0rY1HiT4+vsGXnfDcVGJbzK7XvTVtjoHjExQMamDAt1qtOjwnkj9OBPLN5JMb1DTVUgtGJf
mYd7nQVzO3tuKD9aqyRR9R/QnLrjedovg0Md7IZ+gcpua9NsFXBaRd6menahm3D2E9xcuAlAJV4I
v/8KTl6ObBQcmcTs4Dqb+WtJtJYGwN4mb+t4E+Xp0VPCbZD65bdJtPflBsXjjxZ/zS6HY11mBbdW
9z0YD3d8fKFS+Jijtn63XGbh3AnIg3OGX5ZTDcHvfQxYtSZivJDjTnx1WPukwjdpPCo1SWTcRM2I
CPm46sN8L/nr1KpAjjDUfcffx3ylwMnPGvTFH1ltBNQK+jMEpVhxz2slycWy/zW8SZjzaUpUS+0a
SFwP968+w4MQJN9E6sooAQ9tez/zYx7j2l9xoil1JHba0bY+Pts2mdP5xrjBV8qqvhYDOxZ8SOI0
qiVLdb/dr68X1f8rfjJmWp9gdFmXXknu44EP3wkad9YGknVpIyVkCGSfJsUGH38qmtLXIamRxsO5
cLv5IfPPJ86p/21kMz9KsaSFZj1O5GaA74g+ceCVJA7wGhRyEdleq9KTlqyyTkkkJVySvcnJjRtC
Czdm98lDFREB/aC+y47dLz2S20QlVKtG2vcUjiwWtIYkIEnenLDVPVn3y7pnb6GM5xh7xn/h7GxN
66AFH/SAB4oMky0DQZyjDfMLiJ3ZxzQLeiShcMxmd/l3GNZvQJQWz/bGT7sts9AtiUaspfqQIlU5
8ii9eqC7RaY2yNTffGT0aj6+0AgJXs+95/aPfyZOVFdFXcHv0JZ2FlPqALBswkbFj+VAfP50Y58D
Sj/Gcmr08inIGAa5SiBOi7auU7AKFxoEmiFkvvw3YAU9uHoteHjOvOHvBquVPkd2Ve4JWUSXxBhy
34FTNR2tIaio0oVCdBDO1+6AzgE37bJcficlfvg1HfNE+9Lb4nrfbnmF1Ulzwj8sSSPss8s8SLmX
V0a4VZNjFG3woWhoc7Mc8RvPlNbHDz/IHdbNdwASfd4vXszE9LPpgkpnzN1YEK5SQecmusNqc7/o
QxoNulciCzBEiYRG1cxomj5LRpkEadPEpqbgb3Cu6HFo2VtBDzVyNfUUzhKpGsSArGHP97UOkN7d
bynogj+6GxI0P4ArHmMNWp73sRt9WrRkT3WmeNitEPBlYYw6Rs78oDuBVXmEpC+QP+hrKWrhu8LF
qxd7GMeUfUMb3Dh258b1/x0YkiTsoiYmUfPs6GFDxX2GYTkyII81dBA5974weumauWln8Vc5jngi
VZup/EkZEhEaW6FBLZYj4Hcg5JM6IyeQXg/IyXrsahM4m8jJPz6iQyDnzph6PIDEATbfG0Jp1vON
j/EUW6UmCdluYflG4olAPDnun41IngNPim/R6aey0McpM+mR5aFJLqNPtisXFyrJETPl+jwapYIa
2E5Zb4A6ESjDB3Swp//9S2FnSiCxzP5Rgnhx5T4lQV0leoCf42RCo0DoECGjetgwxM0uicmyDE6Z
dJtQhoOxsykPvpJ7Gvp1VZtqlGIp15nLmnDogLeHBvPYsBl+hCRXvpsVUneUFe5x+tTqsN2tB8Nj
myKs2+xrMKALS0IeDMH2lU1Pwz0sH36n7idkCyILenf2S96gNO84rjilgeY57SgPahoqNuklpYdT
vNtFl/Gb63pix8eszplDoEyWpSdFj5Xe1Gl3JT5MeD8zwlOkEoTucOtL79IqT9zu1eB7mRpeCsyd
oH4FfxaHpOW72MmfBY/wnU6ZYKj+jXhPD292Nl3WnpsyqRqHMJK3wKQwlFU+R/x9WwLd1M/g3hT7
2JZbL4hS6mEebpitTKZCMxk+QX9pEDRT3f75G9MjRjhoQjujiv9mrDCL108ruKl0gJzEuxccZSul
LS2+uX2uFR2YEWBQQI+n3vI8mlTBioU3Sb7U5gslUDaRECbjtXih7VMBYgWJcNIClhse7w93j78i
tKECn5c5Y6QD2lXZc4Irn0yE+RNrf8iZrOV0CXiuiljzitG79riBY5zOAomeT2q1SePUL1gG488j
mNaUjJJnH6i2CrC+Ye/B6B5x4A5QHNA8uUJ+qVPuXX9ve4Dc75MwnyPq7W2m+N1dB6uiZ3M6hoRT
6Jbl0zu76j4xK+ZLeyNvhQkXcbN1PcsD2qYRtB8Epo91KpYgly6Cw1NcacQcezhjUGqVcsL2qf5R
p8/tqBTk9Edc5gMd5NbVo+ee/DsmekizDcZacGOZU+kquOou78Cg6Adraq/hqzGQS+YcbF0jCVvj
CLv/J62YroGafJUTJi3CR16midK1CbxpR6x0JLDQCM0L5WYOIjiVy+l/w1X/S45IEdude0QTyPGf
v6yfYG9awdH9hBlRhtARyp9gfRnm/88L80KPFDDciAZb/q4sFESMAdiaheOcu9FA3VAfOxarLNBD
hsNcBM2CDtmKXheFRlm22uf358ZZvw9uz0MMjD9p0DJAPkxG6IIm66Gb3pQEHDozb7OrSc0OgnEY
mvd2RAxq+gwizDjpwpcL6FRrduHTqOHbAAHSgPc+WCbxWgHJBKwFM8mMyTCVTRgfupCp5vOhTPqE
Pg+zjESIskf3NuvJsLQM1VJ1cbQ4Ow9i/Ok8oj2RmgrYSslU6gOtMQx0hUOXRO/pnwZ/ZOor873K
twB4I+LQBZlXJIQXasZcem4VJ//dO2C87jymf1/Qu7MdFw38xBLg17X3T7mCR/Cjl2Ifk3QVJMAy
O728qllAAaHcu60z7dVrpGJnaheTcVUj1Epx6yaAhfyHKilQiJ2cKxTpl/W+iilBaU7fKUZH2yj4
/cXOHgwj3kZSuSx0SpMoe/B0g1V/lJ9qmrkT65/RD9KkNajg4gXEzRTtn4Ez8DRl68VAR+RXE+Mn
euWrZNgg2BjSpi1bAZ0xWO8A+9+y5UPM3W2fBaLbsUCyn6+1pFJN8Tmmw5wKEVzV/bvmvbRUVS5m
GCMQNwRf1heV4UhPHUpi9Aud5CD3YXMj4ntBGkK6VPY/8JORitR99H+Ul9fHcjUr1Jthmur6zPWK
6icuNBG0YwQ3xajz4BkMqLEqcw1ackrHDUp/Z0925DLl0UJoZbvzNdfbh3bYwqLYtT8iP3SrUxCo
MfrWaan2ZhIdRAwWV2U6r/XKij3NBsHRSppkGxbjF+xOC5DHMq3QjCelv4oqRZDbT0XEpOHCf9pV
WQ7tqnkmMkGSfCX57Q8NTpErH5NK4kvayMxlqsustGzxETWlHdwYk1KK3TNmDFXtnEniFcEn3hGP
c15P2l4qWYkBVJaTr61+96+It1/O9yUgKTc6esq1nL+Z3iIoRjq4fZzulqZ40gC2EmQdDlsZNFPn
paSMMJQ5GG3NVlB90Ins7ZGUy8+rBEGrH5xyVBgMYVWYn6FQ1VXmA9QGcASXCvK/Edc6Dmp0wZQ1
+YsoYj5UNGd6ITxGVDlGsfuVIAE6UH2T1wLABblDNmwjnNhe62dPr9N1Ud529UkDDdClM5Y0jkUX
wpB9+iwXb1KEjhUIuVxXv9JbEGCNASaGopYg8M7djmcwII00srKrfKY9KcqsnyhlpQ6H6S1wSPKO
Ujlj8Iq54aWu/XVNlP+1x3RK9hhbty9utCAtIo0hx8ZWm0pKl33ocQcrPPjCe6SP7R426SUvbGBH
+mz5vWZwBJUpwWpa8U4eP3zznkv+Wb+J7WTb+cW2TGfoTMq0JcGeY+GwtIuUR0l4efoddWegCVaM
TVEl3keZ8Vytxsss7+2RGk6D3pKqdVFe3hJa4cZyDWPmOwVTkO/Aumaxc+kHUNrZiPJ29GTBwMNY
PobXsj1XpIIlEHnfsIPmiWM8qszcIrm7jAdV1RywvBwyC4wCCMpcleEbgP9v+pfOPtaM9fOAAj+9
EHt/URvUPztL1vxvFUo9aVgXyz4Vm7qe5jjuTcQLfU/YzbU8hhjjbLieNXKwfOpr0UOJp11p2Ryc
vynjEAOo0oKDqaSBLvBrKhdaqZoH4ooQsuZhl6RQjg1ULNjOYr+wTTmOyVnmblFfZYa6MaREwxkw
qqhJ/Rp3xhOSW7NEjhZwI2egbS7nVJD+sUsGoltnkv4zSJwA+ghonmbT38ll8nOPQcLAv1gcsakE
tKKtqxQpQ0awcpMxmwDbWjb1faNywo8hXZ5imvK/Lv+FtioIv8PEmEinrTXdCcmOjlz+jeeFO/Nw
oXXTuM+wSSE6OvHTgfVqNZsu2nmIW3IzjT8BCX/lQZazVFc573a+VSNhK8jbPDuOTiYTvtrlpht3
Gc71XLw26ioSjqUEpRU6p+6ENVPoI8iRHoROE2DWClGYJihZeobC3rrFN4x8Mojz+jIczFl0rmGX
J7fJa+O7fJoSyxQ5JQ6sGYCgMQmtrPiEXeKmfZlvZfU2+eKvpRQSGZEqNcVS8sYiqK+FV34NDYx1
PPh2rmjhI1Vuxaw48VJ0HrW1A5pWkyrxAzLC261+MEvPSoXXSLagxYcrecu4iEXu8r3efp0RIw1j
fPbutAT0Y6YtSJjFzWK4F6tCfe1828mQ0FLvkDdkuKesBuDfnzddd6B0+DGg1tyxdOn93JutL8zA
r/hmmCBsNqxKQDWVRTYKvzYPATWM+QdaoyZqwa9CcqcZGGLo4JND9T0aBmcjFHIcxWMkholESZXs
dYHcpHf8pxDmrzUz3bjosZmEmF3u4Z6fEDQZ4hQXSdEi8Cfl3fQxUxPrClpahSpfxIuk0Y19G/A0
9Bdiusjb4+T1gx65M/ISj2FoOrdRyBXK+XepcIyeTDZdreMEjKIaNkwtC0W95c7lmbS6sm2AntJp
8rP+KhD8M/4rgOsbFOw8IYCAKUJfO/60WfscMclJqlDOe6CSot9zTauBO+YO8kOpmaSsLJqB+4hO
y6jo8p/Fp7gH4wcXrd9/fZpxqlAeFtX4i/0d2r1nQyhNYNODro4CKdyYxeVHaNDTCp0rs4aEHA2F
X/9iq3Zlxc+NXbuJ++9wYNOYffek7CLEAJVu2q1KHyHJZE4jgNzfkkatwD2bDRtWJ0GZMmrdTF8T
pFUL8Y5/2kTLjzLf3X40puf9P5KvK3O0r5BIBH38Ul5vwjrI1vwgEIXLcCmk6CysX7+UcUKBu3n6
/BF4ZdAnZrORpg/XTdTo/fBh99Qnw/5s9bJfoq6DO9X9f4VLFz8unuyGi4np62sP1s/z5f8q1RAE
ZImZ0ybB3qyTY1PFY6fGULzPYzwUNFnomA0y/3AZW3XGnNblBrANvNbYj/NafSFBQD8jh/MgnEk/
/NtPezV8O2YNO46IAd2NGw17OQtmp4l/SiQBIu2r+zv4/GQIfSq91T5udAfMZzYCCsQVz7wfYjAn
XvNSa3JKI1/lP1hzXZhOxGDyR4B+yJCpfkiN2oCSCufVUR1YuCV+RyimIDzyc24iqCft+c8uqOEM
x6CszJqplublfMCpPGARBs9A2ZdP6uaf4MLGCI7r6UEDvvBk1xVBuyt0Af3BL6mR/R0mcJng7DjI
5ElS6JQMoT9cEjEB8Ya5EDpIDqziPGw34wVhy4HvL1NuS3esC8IlVOwA1VtRt90jCWbY0Q0oro73
pL7ncs7dvKIiBPj33+OjenQj2LgIzFJ6hBI2bqfFKsDOFP7rcHHM1e2f3omi/kj+CvzUO+yvKHb5
geryJoeWm/RTY4akO/6HVDKznXzWw0t/oDc8mA+kI0Dbq1Wc/sJF96yOSIuf3GiE9rZ/cAlTe/lI
ly0GdUQwc/yAx6IbJ+GLgWwqYXX6UBeXJ2j1OiFxWI/B8Cjp7n67CurlBH1abOxAgkNeHrzofgNv
uiS8/cXQNgW6nwFAmd4Ax5tOF/l4/BAsd7aFz5Hqopklbsr5bYAl9umS+ce3uU8CND2wsitAkwOT
/Yrjsox8srJKHW8kLgUFpYI54h0Qq4M3yQrXVM7bOosne7TPu5vvM1VGmDmGGSXytvkxXjHYyjto
ZDjpYPXzeR3aiCTP3qFLxHQze1IpZcInTjFhUCJBB+AmCtnTnRvMax+Ob+SVus6ysL9lZPx97pep
Ftd+vnZ2GRy82eRx+rSXQ2tG3mRaK9Mo06wmL3GcgIdPknodcJZ7EpDm5X0JOLaAKAxHGeoI3R+V
VwC8vmimEkxOYM0j54TF228q7ytJEr4IP7dtDWH42PD1ngNIYESwg2G8NGxpp/A30Db+B7DjLzx5
bo8Id7eaZUQyeL/Y6h7eJyL+Q6W8zawAk4VdKIj2LsAHrF8RTlJYMVn1/R+JzKClSnWYH/wtfrKS
dJ+ur6Qdvz0AfaJ1QsK7dyji/lExsn+Gn2fey5xG8f5UG/zTSP+7tk3hencpRvx33ttvyN5HnNEe
nGBnGN7xogjAHRN0vj2CxUJprr3C9i8Bjoik7GEhqWZ1W8XSNFIC0O9YQgDbNyaiYOwdVZDSmYvV
JS0AETPh/EJaysLy3b0FqaWb+Kwc4d3hVSSwl6w64qmWyIzeiBqDlLWDJHxnYTx4wbuyIeEl4rlA
RfOR6QYwgbLwsT13vTz44tTcPI+mYR/kNxcghzI0cXtBRiQRjtWZL73OKe8ZALvjexms/AYSSMMB
GVWzGWIXtEz2nVsK65bu22lS6w/sNfwu7B6P1+62MohKZgOOi6xrLVFbpBXg4+VDM4CojC41SqZF
xIbWcgey8QQ/c54ZbgGkW+VuzP108iLMVjgEbJWTe0Eu8wlY523i1+qGv7Vu17u+h3aJzLe59PcT
xAeAIvCUXHRuBhLHqgSPAVY43HsOwP8SUGDFGTnLQ2lD3TSrB0Es/gCFQoLFrSyO1hs5LY8u+36x
zA3XEyQte7oMOfV94Il97NqZ33sKSMz0dPMjymq8HNgHTJyBwk6eewA4463opiQt96+L96wl/yiW
f/G7P/JTdJ4stp/zTuC/jlzbvFOTCEKVmYHNNMbBnek+PJqQtJiOVL2mvTy8y1L0Jj0/mcxp0xy1
pr3xfd9FIp3z7GVJhiDW+dcpifQ3NUZEHFVJwOAhVejI373GCfetgmJnCOQhUIXdHYp3jQNci4a0
/Khil1SeaCJmLLw/QrQfDFekuUfTO6m4wOJiIQq7DwWo8VeeosA0B0kiogs3Kl4yP+AiZ7CWu8TY
40A+9/qtcavlpyukbvTDNZynN9WsZQpfdneEZHH3MGN3Pl6xqIG78mrsWUpkzoEDzetoz49TfYZM
xHSavXlHwB21YubnoGUJerYEJoeyH0TeLNh3NnZtNDkbomTfJ8wyif2QKpdY3kX2/q8683uI2dYu
oT5bLC5bPt55EkDmb8W3GcuiRCmIIV2dhZz4THY9i3glNHWxBxdfWUm8+FLXAe8w5Mm//MKUZo6r
BRc/gR61PeHWpUQGwXbh8myQTf1T5CqIgl6aDz6usnN2TvCxYM2c7KlCQcUHHYl5//rNmY2RSWj6
UoAACyo8r4t1zv55w9vP11kJdz3Ru7XmH5PPxZ6Fh3cczx+ragpz2wMnl7jET80cI0LaLMw=
`protect end_protected

