

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
F6vZD7oP7yEsXSGX9Bj8IlGmCHNHZTxr0EqFLtf/pZfkGGh13rIajlApy8+H+IUMAvi2SjrfWhM+
rbpo0EDpgg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
C6AvHnapQTJq96+XRFLqWPzjjTOUc2Ch++roETe7nfPsKK/Q1vK31kjZiTRBIoLF27YloaNJtyGN
5tb8dYgAKEyoeYhXOUsZ6VUjZWDgCclwj3wPZDV82XF618ynfs+seL/pkqyIm2lTvesQlcQI1wFH
/OouOB2XhRvRvj9fHCE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TLg9x/mjN5uehk+g4R0sirOXK4prtzQScs4Wl7zD4dOmtc48pHBzEpo6gak5NVR/J/qbmLHIyKJN
jOUBEPPdf2wAEMPgrzYx0ip60YimIXynLpLSqJQ2anjmR+ZH62WsSkOZWnbN6ji6UZyh77ut9tId
5DKEd/rDiSasPVyA1aoDwwgYLdWLXQfp2gP/r+OsO86Ly6vMvnFbHwFuqEhhwlokry5J6n7pZUId
1BNGIIGdg5NF2/pVBAyc5oY9sXL2mp+nUqo5ioese6LS1WxfScxYkvWS6A7W/eRSA+Q+0uDwO4QY
GUmYaxD5CDTqkGr8Gi6Pfa4Nqh2G1ovw5LkxBA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rzJnGBzniOXYMgWZQhUgwFsF3/Ftf4OdJdLxelm8+Z648E5Pts6ATZ7lgb2rnAtDE89/7CV+B491
XNnnrNB8L9QtpC3GwrIN5QRyoO+dvkdY2d1gypiWErN2kjNuoRWhHnaWJ4sERUtCR79UYo/wPTLC
Id4h+KNFxRbvY4xN3yqpzEZFL4eGkx9H0wRG3UHKgmWVrW5y7PNzWRRs2CYVoIkrshHAsgHzaCOE
mXlrER1zuex9CrQ/kPrp3o1sBLWNOobbDAvzi92/n9yg3YPASs0COd8zbC2Si5LklvC9zE1z7hOZ
h+gtRFatxmR2vIstGfhYnxcIeL9SiWFVtrZJ1w==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iYSfhRf8uN2NTpFWL3iQ28bDKhCVfXblEBICf8NzPpBEhA+WxeGVqKUIkI5y6xEegexfeqQi5NSk
0F0u7adkWJA90Ms2lZifpMaTtX4Itjl1Q9gk0vpGdaJeHwbwPJwfwAnni1xlES+czyWgXo/3pbHa
7WbdFKr/Mys1aIAHzATlVBdMvEVU7y633Z1A7stVnx8D51x/7xkBNn8sQMsi7jA5I8XlQLqVKRk8
ru+L7R9//ydhyCRZCgy7QEfvF395OlAL6byLhkomRETmktIlOsfBUU6Ff0qKxNqLnM6fyzQMBkVq
JvEQhRBjn5+uZ2bYVRGzlY5OPN9VLj2UMqZXeQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QAF5a/Yra7Rn5EnGGubHg/HcKhsF9ZLpk5ZLxiNBw4pHoD39IbG2IffecZBxNt0oKTQk4jhNLXnm
yyCWEVxX52C2fN4Xmn4WdTHcYUemMdx84dtXH+l6fdzswTUdWOSznMaiR1YadgGVRObcGMy3aARM
yyR1t8doiG60oEesyIU=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
brBQUuW2YAZU+kuTuwMybjF9u3nQmOP9axVkBY7fn+Cn+4ByMT/xR2U/NtIGMFOlR97LaKmcPsxo
+OtdgoRW3h6R3LXPnwPlCxhtWXv1la0SVi0+nqEdXXZZu9MFtjXIMxQg7Aq4AfXFVPPeyFtudlzP
qJgw6kQqRB6vidxRdFG+2MgsX3682zAgf7Oj8l2F7KYKQXDXwWSPm0fla0na6dz9iWt7q1lkJB+C
jQvtgpeeS7LQPUs6FbYT1ig3ujK7MGU8s5yAdmatc7LUaNGbsW0hDu1vweXKpORr/JlNLWZDWrzX
V3kjGV/LoTmexyNf6aKk7VHVpBekpbD1+GeRZw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 506768)
`protect data_block
BmXTD4Tib0rOWAdHSuLPDqbdaIpvDBTsSu82ZNFtnwHh/PUdT5afo8JiYNU/NwUMiuaS21XZ86vo
cipPpgmETSfQ0fphvcpnAvT9IBvf8RnXzmFJKe0LOWe5akYFYZ1Sele1w9zB2gwtJX8dDUcve6iE
jY1ygo7GfeXh1gUxW9MwVRatwBH6SPL1WkwW1FEaL1vK9PXVlh9aQj9GZc5cTjZ0bFbrBvGX2Cc5
mgTID0UScNqOfhpMFvlwqVhCy0pTfIGTfU+Qbyc8YWCyQ+TkFgf3Luv3yjVDoydushtanmkof5Ie
oX7jQZxYxg9/ftSyd8vo6LKpJ2lsJH6A87lPzzKtChGCsP7xvCuGqhIJfxQ7hsVnhlttJNr0gMs7
FYkCc5Le9qFAIwaTo7ThIhEQNNai+PQ0BOuzHaHZMm2DIyemEjUPLLbvccIR/fvehY5kiFYnBAoT
TTQNBUvPPN9btsbbu8+rsAXWtVeVY3c8vVrdxyVvosFfxh07W+vyDOdKAzuQviSMcuNt4KQ0KWLy
/B+k9bsa8wLi4++MIIacTdi5Ue63X2BVHzSut7q7i8OM5eT6KVauK0jQ3WeGFmxoPBQcelmdk+u5
yE9+uYR60YUukr//Lk7jKla135JT+A7vD61Fvf0Oo5t2ZatgBrqw9Yks6NdVestN2V37+ucNRS8s
K4J6jZsGTXqfJJCKNzCk62qtG5WIINPVyu1K26fbqkuzVHYQK/LeFXucbhVw+MPYzjbeMZHJISPz
ClXw/n9kAndrfvvZJ4B1vkHpWAk7JOglsWe8W9FVHZNB14pUVcKUY7TeU3f8kPz4kCx7HWemw7mT
4Y5kr7Xri8ZlVSwdvZrM4VFYM6OCnS1f2DERV2XO4y1czzHYMzcQ5579/4rjmAZaP/xhmp53IuHP
hYwoltXLDwUDW1QPw3tQ+Szw+v3x9ulD9QtaXsULai61t3RyVCyDVbF3tN5K5gtB1A6KuUhqh7vX
dWjMQi5z9ugpzFFFXOhEbv5LUW0ykIUHWN6TPVqrQ6Zr4z24l1WHvNmik2LTEukawct6zrXHoAjy
R116PyoPfj28nQJ1zyB4fhU0WBmPP7RRcX/0f+3DJbZzNxFK4Fs7G+TkpMomDKvocL1gIa3bD+mc
/owvAWkMoL3bTjYMCaQIsMoX4KnZq6w1a3+KL2U8mpo0L4jyRpgSO3HzPZzWH4RKrWCW7h1u0zkD
Z96OK8aJuBnVUXUO2ASuDdcopgh9/zmWuXf2CCEOARx28lVU5OpPsZp4tuwxu37Q/v/Qywdsr6qg
6hOAJVqx8f7al2uzM4+qmMvBHHNvvwgK4aIyMZqbQkXgXX5V+Bj5SGDSKZ+TA/o2dV4hIToK5w5W
IiWHAfAaX66DVexH2Iiyx1HZXxsjBmnoMFZ0fp7GkG/YgO/3k8EY6HBmjcXMTe+cyUuRvCxFzuDq
g2HKX4NzjNIwAztSokEIOjrTLV3h07rO3aY3WBAooptFwC6AL/rMLyVHHRBsK/9d5DijDwzZsTNF
52e8Y2v66DU/RURUdzv0qrMGh/TUFixatkEfA7TNf3mEZJHaqGrlGJ9eO1wh9Rp/ry+g29uKJU5x
UpJtRQrrjr5axD3EB5uYoc/KgNWYSq3LdeYXGNC5UKl4a7gKcxWPr7PJvNoV1nhtXf91DxoWNAK2
/BEgARui7qXmFMgJr0bGwrVAp65BOnotBRrKpi7iW3lI5wSj+8UhuAz0TBQC13Jx4FaD+fnYTDP7
fiNrPizwczggaDRa2uAl8IKJ4DisJxqneSkJcHUb0ek6xUs9vBXEedlgTKplY8myHRqXYv8OVtvx
JEMTRdJo9kgoCLJBNnSiyrNOmdvUQIZsQI/GOxEFTK8b51uFOGm9GZnA45PhlN0xYRGjMLesFH+4
y34Lv3D5eN2xw152Vw1U/L0DH4JbmhvFadNIAcA+QNuAL+CgXlrb7R+uFrqFJQI7zvofOpD43krc
iipCImZ+UQORZEiE1hJpL7OtsUaf6f/J9sR+lXn7xjtPxezukcxEKK1TN/m9rULMvKg4EfehiOzA
R5hgib3XjE42wVCcgeMmSMXHfRJwbYYALBpBE8zrQIW9QuyWP6a3NO0FxsV09xJ8Olp75kWXXDaE
qjOAPxzbYPb+lRKXm4c46jpIOmM/Ht1pfL/dmlm3QvFBW1JduYC+/QS8NWMwi082TK27U/G/vu93
z3Hq7SsSbDM9NbosPc5ZaN8cLItxZtaJKpymWHrWxmb4h6NZI6GvWjraz3geWFyJzNyV906OvUzx
MG9429Sa82eghap+vn75iwLTmdDs7nEL5ehSHEMbTaqRrm0eT4K74WUINUEZyMNoytWAk2UtqMoE
P3wIVCizPm3r/i4NqCi90U1dSiXY/i1MqAIdYUcUa5QQtz2g4AQ+CzmRQVXbOt/H8XOfHPlI4l50
qeER5a57DVGWi9kPEQJJb0+D+j3UfBn+GReGGWZ+25WFo4bYidrWrOKj57QOhjr8jdKBl+87z5oL
VcSMpfaUsY8u+6NuVi7YFzBJIWUCgD6xw8Z3KJPXvSSYj0ki08WbDYRsljTRL2NBqtub6xepMY4/
52XQo488K4l3dlZAaUZj2aJ8eslb2m63dq3f2tqvMxPl6462IIctr7r6Mn2vIIkWOPD1ZAQdB+jn
uI2LqR4ij6uhvZo4/JdzI0xx0iCke26kjTHxuC6k/y5VzuzeiV5PAP50GgxlHztMimhrCLjJq1SU
1yo9/K+gd78paGxk11G5uzXgDl54rIyDeh7SgwFuXULDcfM8vr3RV0b5nJ4SXUYqwKjjwBWpiSWe
n1LM/w2FTl1rv7LR0mYl2i7ioPA6rWKBbfFjJkDZDBEGKNDESBwsxKvBbVeRaYlBUK3NQlUtzgJ/
NX4lt58vTK+MWCUxbcC37dn3BX+c6Ghmb74QFMwvidJxAvN+/B3U+RtjPzi1F35UfgqRciQRsPBb
8jhhiGlZjDtUGnQ4Xz+7gMtUrCVuqZYqroFEWbrXtbKNC2Yuknwbcj2ud2QrLCPkqMx8X/5o5tXG
dwMwZsvgkVNCVKUxISL3uSDaYulyHnfPS5C9Sgo44NO1ZfnTFD12+Z2rc5KamacolUycpBRBTuih
nl+z/pDamOTXsY2NID20V/nPSveuWxzJjafD8h9YmIlXpJW9xeasJmqKOkSM+EWDAePOF0YZAYsU
IcJL5i1/SVRYvFMdEC0WyBPOr57455ud21rB63Tsd7U6oOBvnt6LSHM7pZnw1wYin1VClZPuXesg
wdKv07qOg8VL0CdrAvD8Ria18YQlgmuQrkCFL38Z2K9IjEZ/pKVAQYwHweKXMnGP617BYhNm7Tnu
RUEgUVgOQYH911HlC4KX1ZDbM0YIDSshRm99t8CnSl1g/Rxi6Ertntu8sjo8a0rJUld49cHkbr4f
A5Prj2XBE7Qpe1zXmyKu6X6kTrCgSBA7GSSZT/3G/b6pQBAeYTDHAOlHvJFEot6v5/X6X28F8peH
PIvHpf/AqfFVoi4GHRAGHHUlogECI6Q1fOVsaRFIYY2esAmbhvrdOv8ucRIdJZ64JsbDGa5jgtrl
shsfniw5asRkNL1KZxPW+nGJpfjH+51moBYydfD2H9MhsX0KEu03nl+wGRxIybAqZhsx2FT4rre4
i91TKUDAnsTsviQYLNJxzmojVfJW185pxTJtSxoeq/w5k/owSIQ3fIwdjfjmt3vJCaNmDdckH7MO
9PhTNmwJ+2Zq2u+civS/3wOsLMeRAsbJyl9yH1szFQ/i0uJfdklc0UApejseDAF6pcYgYP8O1pRl
841a4ZaRJhRIeDM5tDjPvL+YRF0x1rfGKsFYWlUqgoDy9IAKWOQIZ+Ej0+gmx5htDBdWa0l6BOW1
6xkzrYuZYSCe0jrhR88dKuPsKjVAae4T9mkxBEoAighwnZdYIalb6Qdeby/zwaMIju7VvCrUCv4b
mXc0kKRa39DvIrutId6FEtCT7JNBDJnq0oKwqZzzkR+MUp7mMHl+yNJo8rwPsJ7LeAlJM3TVdSib
O18lVMC4AIDTQyLHARm4ELzBzkHN6YPN0s8tp9uQ+jQ01aiLe2X0nZPLg6GTJ9ffhGqYdLHokv4M
jijuD1uWEXQ6QgOBk3gXs3ow+1GnN8/1Nifm5s5d2knLmp6zPcJX2NvdS/Go2yIvqDgx9ypn1RQk
uWqQn1TmN7eCUyfXnzkUNTiI42zY9Q1/KKwJjNjaEOyuwL7Yazu5zMOl/0zzhh5apC+WdUArDz9K
hDFS9VTz5tCRTPa01h+/U+35QNe5tE8S4uNfQG37Y8ldnntHulfF4EfHXI6wqS5W0s2LT7QoUVqK
UtZEfRDGZlDo1mLCajKz6rOXwDvG6/La52OCl6I81PmsMjSUKTp+Bb+L3DQibllk49/eW1wh9jHH
5h1B9FLZ84hMTLZAjjeQP68BQfMhs5BB/1WxPeFRUk2s5/2w+iW1kfdr1jIiPL4o/r2O2FzYSobU
PFOEeSI6x/M3Sg8xbT3Q7BEgu5KKV0FaguDlavwjl8+gVw2fSBTa7xnRElv7diOBr9fIMkN3QqQw
70J5Ww3AeM8n39DLehpsY+liFzlrtbiIzxcU+1ES2U+Yu22EpUBBEJMhvX/dtm1Lrpr/VBn0xKcn
dalEkRI1pEV3tKCgAijpU2tV1l2y7VTH0fRWiqj26OIY78GqdhFsv16l10igFoYyi2Etv6qe3M75
lhmiP0Mk1f+uTe1deHoY8pA9KFqasXtzgTvd4mmTgKpgIJMjqsQJhyvhTCLvnRhvLUjX9P7j3LZo
Qs/gi0v+OUgvq+kBOdfaE2VfBIEgY4h/hYHoyOeD1lX9zPebBNZAyncvboTwV+y5vOSO8xSiaFDu
qdBgKseYWNI/AdfoD20BjhWD7BYyYfCyML1mTARg2ZFfhk4Ozv78ZNxJxkLk2rkrAC6HDZreljKT
oe16HGbq5Zak2ohMNww9PDYAZ1eypZx/fxCQtLhwyKVPW4Yjho2mf5DRYi7+LyUm362/ZIDRJUKq
je5Bn9wQ+B6PCaTjdjOC8LMNPMgWDQNXEyeP7WfjuIkTTlMsmOGLnyNQ1GzJ4tC81xx+kj4jxTJS
9jqzNPlzSAiZ4LuB+WMQap6h6Jw3rWzQxgaJHd522TDfDLRIqPS89wEd5Q/g5oGFZ7uwXIt3ob2u
W108hgLSMxY6QfItXDF//H5j+1sMAq4tDGQQwbD8+0gz3aZ4TQ7anl7PyMcnisnbHpfFe0V0eS9p
+aqPeDwybP2QfyaGb1pX6G/B6Xxv5S3HEb5P0MwhEZOrkgNwwz86IKghO0LRUFj+aHG6rPTuDqgr
C0kBbHqNYWogFB0M6JpwRmUS+FrzdyXP/aUbIUKpTJPvuzO98mLPfJdge/znea+RxnwbA33mGlLR
SPp/fs0+gK3X/20cUv7/gBawNj4bP68nRnShFZaMc5u21yqrsC4tzBQcoXHzut6DsGAmdXNg8N4A
up3vs04Jf4ZWt6dciI99lSTECYQLgBqD6ieATKK+QFug7vAnadta9AnVHQaSF0RwOyqLAHXMJWog
IoDSQO6ugj0P+peGAMVTN7Efge0oOjBlGM1UlNYNDz1DlSTea6IS/FY8SIwAXl+yW0FZwW3LdE4W
O13XQgQCfGiia9fSytxPlJSrkLCJYv2BKaTfWUbNatuerQBPdcUD73A4j2sioBICr0at3TFNEw+y
SI6NXmH26UozznoCD2IR481EvKcB+b++ATC6mPXo+KxaSs6Ix/E/nItyZqduqEaWK9jhMmmF4w1W
/EEa+/RJ/7NpG0lPNuDRYqI8qlOOL+K+ZY+/IjkK4VoISXFLRFVApUFCa+Wu1gk13pdGuc4mw5yh
4PiByuJkjW1i3Z7hUBtvuVSWNEBDpf9BGx1dHVZm9vatDnnPVUnNSJ3R2ZzTzD/qJX8M23gjZtNm
279jV4CkxdjXDzrk3QytT8ezGkpLuHYDzNAJBNlet2j51oQ07BhIU/hBEA+5ft3E1se4SwogkClX
5sEhYox7A4+59TGjMKC5Xu3WWckJRqVaibd3i4zNFTwYbmqWCCQcM2bnqrRSS+cX36v/kvBg68fB
Cda1IAImwa5K7GZyANUi+p1K+5FwnJoeii7KOYd9N4jGmYSdLCas8eM0lipzm8gqisO1uCsVGa2k
afBnjZ5t1pXyvI7DtdK5fRiiL0NYOsP6ecquwwtfSMr8cw2JKMuRkJzT0Xq/DBM9ju73PVftAux5
2x56bO3FXL2r3FvnYGLTXcYeDeQ8Too/VgIJckPCSw+PAxuWjYRNRDWaLg02/fnl3m7gu4M5+sgo
6A9ilCakKmZfgPux+7YM3dsZ87MSMQEUg0z8Yhyg+KfgpBBwvDY4rjAAEIXw/F6NwW7+OP5gp3R1
tupInaY4BQH4exeNhq5YP6RUMnuc+yQyTaiCIa+l+QBBR54YnGfPW71auZFWV59wNaL5YleHRVCp
m3z8jTmyHZ0noBm9okx9AMKVa+FSNQ2pkIeLb6dlJW7rV253rftz+k0YmzE2nOgGnZ2he6jDQZiM
aDRfNDsVnD6SxeY404ey79kRedsExWofXIfBNdWm+hAauG7/U9Mha42tVn64zo5q02CEHjiYNRCz
Xbq7MkJqOKkyc4eIIUd5EeSe4PUUXh/o+Fv2Ly1LG+bKWu5VoP/dpx1hgLrB/Kl4hDtWuTQsOmok
1jqjve4Buxn4sdJ50NaelZvokI8WWbto+aHYWNsR7iM/lQrelmEr2JmQLdcfRP5/k3qHL4wreF4B
Xo32gjaE1lATRuQdya4d5YQHPLLi3eiqvCyPi+uDAiauBP6OoAKuZuu11hhqNsykCqNEgCSfkviK
59JmFrHI8rKGugzI+e8vMJkv0jA5e2VHjgDpllVvvdLuU3rv+fFYyF6d4iUBJsGJE6UAu7otnZOo
fCReh+GLO+nUzYUIxteow835I+c+9O5BhkKCboGru/ZUl9eESqzaAG0kdB5v4VXKx1sa8VDwR5y0
dxB3hKMABiVfN/yzE6OOK4pb7QitjzmYGhhmM3etcjv9zQeHk65Ma15e/X4LfFPY4nNKDWFfyvKM
Wo4A1OdoicfNWeEMmAUn9WG59IzW0LEyBY8Dypm31Dk9X8ZT4lOVrSVYQYgfsVRCng2IoMqDkMIE
Exj3hXesKB/K+dD2PWb6VlG4MAxSBRuO8fy2evP67Ia/5YAClYEyJyjOwBhCkpKB3G8yug68Unpr
2ZgPEEVrGVjke6hBc6JhgB5SnvLcVjvM6Rx+CShDFJy9eZcsAxcaoDzHCie/xN7RtKpILcomMYLr
mmIBKVWk3ZMMPfYH4ZMlM/05nBfcLBZs1q0h8zh1tfLjmhgJgq2oU4I0PY5FgD0bBZjVzkzNPS3O
Jy8Hg4KMbc3EH9vTG5ecbbWsANX/a199bWyZvhpHLxYd6Bfoyz0t7gyLZss/qH+cOu7cyP8AA/tx
cSauhCYPIXlsbUWspVKvu+ggNhOjWytFYtTdLXK61IZfy8o+0bZRMhfIA8Dljt7zfaITtuWVjTQo
eOp8LVmHu0Iw5hjKxWGoFnUPIELxdrlbiqLQcixI9ssuWX1Wh1UWFs4mJK5r/0ydZbrtjAlF4BeQ
GeUNONihfUXMBPIaciZSm2GaxhzUMeAvUtEgyEyak0yqmYFvl2LUD4ePbaWCgyGcKaftqcqmaCz8
Gmy7S465mj7MgZHrQKg1l4Wkumt4ADoWYmEaSpbMouJNfD51tCVWe74qr2w6HkHR4ZOKhuLXaG/Q
Jj6/tcBxmvfClGjBYEvo0KZI/z47EAP8viXQ3M/s+yvSjobZyjUk4QYjcmtyoa1W3NWVJxLGeycj
jZtnkl9tSZbzMr08UM7PVcqN98zuZlsN5dHNJIcyyQEKK7AOvPbEKlNITwJJ5OeiFynz6h83G+G1
xc1HyuX1OxmAeo9SK+XghTxRFRNWGzmz8602GsMWZpgtpupyamMelct7LVatJyJPf/RgAuWto4Ye
r1RGIbC79cScD436N4OvtRN2UhfX3KMieO2rfuzSbq8MYzKAie5oz+zGeJ5UCcyZR5JEeZKrdDWw
KE9voP8q73v7jQYxPYOVDMY/x7qmX5/Cc+Gu5qiHR4NzfKBotktMymIDRwIpTJzrHb34aI9i3J59
ZDipgwjIT1RHelm1wZwm6aBWdMGk6ajMYQjt7qboyoSbA8mwDwm5p8DbxXLEmh3/l/QwxveqUI22
Sv3rfOH3/ibV+Lb/PnraG39yi9dFV22bqqlGGKMlYI2FDcb99+irBRmEe2EweCgbI5krv+CB6iqa
yt+glqn/GUwUInihBAKaN/L9MXHevPSw6op0bnAcbQGB+ynDxg8gMpGTO6LKeaDEdmKkl0mxD/q+
VpEwDQS+jJVt71MYOn8NRgc5ZHI7iFPWpcS5yof7HIxz9MhsezzcRji2CyDXTOe+2kQOkTVGJ1yh
HtcxYjG+9SwswpVqhFGUnC7UP0w37mRS1kc25kXiQcOMi3y9BYj0wL9eHiOvBM/LjMhrD5gLWedy
FlTav3cN33O2f1JBuGfKLwm/nM1F8XderJYXBoIuifkkNhhi/LHs0fH9JjjER6i6IEdhhjXKsa0d
QZkvFNYDvYYzJEJLxVc5vxE8qaxbcAIa29vmTuKvWduI6NYxv0FZuGv4ZXAYRkLtbUh5dx3wHTo8
aTHvXDNFVQaG4broHmFxZJza8QL35CwAMvIJM0gako+q7B5iKu51eGTPXYRFoGO5rRbC6NgON43s
+PEDLLNO2CDs8E0pdt3H/dQ7pKq46yeoxblPNAl2hhD5HAqSglOWFhFCJV6xIE7/Y5QmGIyg6Chn
LsfOOCVxhcYXVwnJAW3fBRCoOTog05uDVWbeZ97ATmqZztYOQm7wjaD9uT2HeTg/Eukt/lQtkv0g
J7ljBWFHITEHEe8Mb4BWFAGn45ELRaVNgETiR3DKWfEeJHn8G1a1cmG9URPseu1n20QQuWOvjTJi
vVY7BMkNo6v0AXonDLUv7yeHPBDUY3RJvCCNzZhEeA5zuODjdCF07Jd8xSIBixZxbpO6XYdwID4q
v6lQanGQiYzfcAmgGNwPC603AcrQgA6gjqWzzm4JZOFHNrZO5BdyHTYWPd0J3JbmW4IQqcrnsArI
GLIDKEGMgXGtj+ajKlUF4LyFyb7xND/LV0aNJ554gfYwx1Gcd5aw8ETArXIKuVu/BgHu0pOCyDJj
o8SUhYYnEifCIqyiF+LFnu4CTNJFpv03AIdDrlpfd58wM85mWQaXOvshzHO7+oyhEGoJSQDz/nuo
zFySpd3biXviOHEBfl/8A+IWZkXQ2E0sjGtng+dWmY9THZdnWsFOuxBKr+ugUQvXnGbMy+SAvNJ6
DGNFOPpOLsKkedsI7SxLjmjsdt+9vhtnLFett5Gr4dWjeMiihQ+fgqpU1/7qvNvT2w1jRRtfc673
0FL0I9TuvA9p5yqlNgPBZSAtzZW3BZh8zicnq/aWXjb+0t4yo5V8UnJBCY+c67dCz8q8PcVGrwI+
CgsI+g4TTSAm5aZW1BRH//vy8JUfmUUIAL9BgJWi5NxVzOo2KCK7JkRb8FdByAG5jGwkArME1ASB
79ODnYfo6WE3O9tpoYQlJDIgvgB7E6e+MWx51THFkhKSXCEaz2RqCHRDVwWVoPYIYQnaBj9rxbhQ
GMaiRjnqqfcPbymuu2dup+pCrpDT0RBqD2jdwQMcBzqL5C2RJwh+FzWGEUQvgzDLOSe3peGqmmke
zC3kgt3krNzsV7Zvk+nujIuT5GG/xh9ygLXCRNUJnF1E6n8PFT/KaNj5rdaatrA4A5Fq7Rkh6Ft1
clxH5IqD4iXG5xq2fAmqncVP8zs4VBKcJg8zJ3+AETSU6myq5aYdwSUlnsPBMSnwhPJCDZoxF8GB
dQtHJQUz/D7Iqw1bjMFTYtqKZZvQ/eQMPGuvK2pbEBBn/6kBaOM8f+Y1rftIf9hK94jegEjh9BnI
tOIO7LIILHpgmtEOPfLK+kqfAlXQHt0lGW634xUFWD4fMEhzTlZWHRPsc45CgCBJe84CQ6h4G6+n
0RmkrObl5kh1iz3glKJuq+F9qesOBjB8hv4/FvTXHEB1YFR2cJwRp9xJJZMpsV5aPPcw5X6Gpj+P
fT906OvUkPk9Iqw4KQ4xy8IpbzTlmMgW6eR7yyrNINPNEWL2orswGRpjadg5DiBDgKaRvj4/3AyA
WkvtYCSSQJuqtc8xcF3Csg18muiuD4OXAphz6m59owOkUuxUscITs2Cto0aR80JXJlTzP2UiwfQ8
fxPT5QS3N/TC0xEWN1HjMQUmafmd6jl8TRDDq/lWbA9TE+3EnSrqzZk7fZCI9CE7NItLYMB8JFLt
Q5dWFdUvx2J0LtATQ8XokgIWT/LNa3cHMTO/dnVksqsyutaF6nDsTa6gE7DkVtO92bmQVYesAnbZ
5NgqOmn6syfdrnQX5/f45Z+dpAbrHdF13q8csPv4EvF0pSr+yWqd+xFKvwnGGYDTXWLbl8SsPfcC
OGZyZW177JJIwYIFwVLyw0QKOZSd6zadVE0+yNjnWSHvktceV+FvsrQYlu9QyH3Ts4VkrMFxL1V3
wsNOLIfoY4FstVilQoBUFTsv6KjwB8IfzwVes7AWpcmpeDXkXvq06UbK12BTjqzkj1jbyamzlOAb
zbAwzBPvZ2CzQyqQfJeb0J4Bd/A0RTG05g+aT8ktcQ8f0zi54eBUvYgbOmWtxzL/MX+8r52938mC
7wUEElcsTtzMeLY8/kSpnVTgjfSLgrJS+gYqHooXPvXY7bRnDzN+n4FKou/WkLtJR2XVw4yKd1EV
vl8S6b69jHsTpZMXurCpuLSgYJ58bV9b9J6alVDYRZMO3RCDPfU6sAvn+DspEVdvqXO8PR6cwQ1o
TDgvAF3kH2G4UIi74dHm1zeb2xm1Sx9owIfIfmwWSTnRK3kOzcyUdw/DAPxfG1BUCjoQOqJFRlYM
fUs+P7Zbmv3LbJI7YR/P3KSrLQuW8U5QmHMWmhdd/f+8qmqPQrB/24WNthSEUqjvLaU/AtLvI/oK
+ugGTGdwGNMthnc0gfsFnBWpyPVn5J1e+WbqSMMQxsxiW1uaoPz9LGs+LAHqo8lDpvw2b9COhFXg
rcA+dOYX8woeMxdQERdpR5eo4UTdv36ES9b4mhDpkIHB36AD4FW+EoFfY7zMgSkn549N8YLWaWfY
ORtwYV5sOzNt5hAKQUPp9Q/bqTdtLNECFPpP1idSNzuq+NAnSwU1u5zHWw9a7WHy14l2nXEG9a1t
+6Ju1pIcb0r/uEkoJobiMOAKKXACbl3MEM6L0y2QYAZqulaI/BMSBP3L5xCG4pXDK56qMhmoxu1g
PIJZUTySOjcabxeNByhLNaAqxiCSmTrJoqMASolhBxYo/dbt3te3YT4AVnN2x6+jPqM/7Rk1XkQv
k4NX1iU8Uaxz0wLFpu91wXTpjxhp/cXw1zcojkk7tz5dppKrGcG4kIdGdC+uiQClbcZqlhXKm1/V
RTtcajtxB7Jf7WZRWc+fcYXVp6bsLDgVzRHn8K7cK723KR3ppxRAUgBj+ZnwMwE66Zs0JM+TX9vU
enQBbOs5i41239E0yY3UQcSpZOGd9uqmoXIqvtWZcj6uSLTFJ0y2DgPPnveVaTbUoE1AyI5tijBy
zE7yX7MARFeZVvYjNRUAdtrNL4VPXRJmUWUwV5jiGkwrZqoNkhyLil9P9SKMhIS1vXFE8PiWUKHO
sKsrQQt9OGiujb/eSKwMU+M//jUj4uQVGmyM4otjVzC+d8i8VcLBbNp1GjFjnZK6Gsw1yOjkUzIU
+2t71y4Olmbt0lZQLI68/J/TGn9EdNCkkxPO5BbiPrY1Ewn3FXOccJJk03FP0dFrPb5kRqtpBfSn
3w7lS47JFbWfk/dLC7KA8GLdwmdjSH9baZbkoU5D7i/AowlPWtQ3ZPIH1stH8raHSXwVDqPhjaJS
Ase2NF6x2U6wncfxCBn0MiN2rEIhQS16wfZXTxJgwWThpVM6mLlhwVPFJNGlcBpPhoK72+K25hGu
U+Ag1ZmpQ6XjT17if0eZhizOfLTdn4MxcLRCkzuvfn9SLycv/3V2xP0gbDB4Z47goeKqEhZfYeSk
bYgx4MmeNxZnb5cTZhByqwxlc3xRKPU6zTbpvNxqhFbxCezeIVW5ADDioMcEVdI3mpqRfeCHbT/G
QQkLLwrPjj0pwbiVJZ21dDcTgfFFhxK/kQadGcBIL80ZohjE1ck+WpJClv390DzQgrgNJga9ON0y
usD/LImhe4BmX3QasbeBP046V8KttXQkyIK0v+0DPn/1MlOEGXHUrsqg6RHYS3UV+nl2YiqUZIrY
oJKVIcaoj1ll8wx7K9bIy3t1p68vc6KS9uDN2QQDOwvuNLw/7SIJyTfF4qA0p7rGML3vCJvqjQrk
Y8Q848QdYNELcsQpB2Rq/ZrCgrUlkdqkL6wP2S3WHKZVQ1S84LfWjQbIWxoZSwi07HYHh1cbaIWQ
0+eeETstsJUG+lc0zor4CY3rniVq+5oQKGftAgNrZw+jhwRWDwfGIVjnCp/ZIifb68j1DzjwDJwp
7+tKTqmuDp5Dc/MPE3+pDjF62ZQFK8be7m2FFo0ZQqcV14qdUOLiC5/ESqNGlbd0JFirzZqKSLMG
c0YU34d+dlE+Q3ooaJJZPqPgwBUWTEZM4jk6MLBNx4Oh2MyH7SkdAKZuaiTbk18uzuswc8Fmcg7Y
CklozYuwiJWFzXL0n1MLqWOgRQpZ8dOIY1RWwfi7UrBjuAXIcPm76xYLh3N8sIwImr7BNRIykt7h
tweI5PwLGF+YpgFjfXKcfT2grbGImd5qf7DjeGuAc5A1iCy/eJeGwe1d8L3pXfgrZhiJifZOK7y6
O0hNADnWkTnPHHc40IBmwjUnsL1lhc1O6RuovW6b8fW1qMibf9J361gGndHZOK5bfg4I57+rNFDv
474MdeRDO6JdXAhqe8p87MHfb/VC1IGkLn0V9zoGQ2v2zHlOfeo64Ae3T3qYof2q6ik2fM8xCIE5
1ybZQbYzJ0+S8OOF0Fg1NifgU02+U1UR+QdfHuom8HKm7EEQwRcsOyZNcdPGxjRVQP8LD7VQmx8p
iRJYbzmJk6+DMi5RnOcT0eBIw3jgdQ9DVimcrVwa2JalES8cGNRcAs0BFs8gQe0YaLrjkQwHjD0D
yBI5FM/imHhIPszlhRfPWpRnMa5blqASfLFW1Y+mic+Yt00QqYrPhymVsswVWVwTx/n5V+u2abjg
qPMufyYl7I8A0PPOCRYrz+IPJreXsByK2dEmXfgY7WYAoV3nmkjRtsQ3xlZ39HUQMRvtc6E7oEV+
bHvaZi7r+RW89ywjIlVcO4LISqU65CrK5kpWpLpJtsfz6fwXq0el0nb04Cud0DpSF3rbhE2UsE3N
Nbr1i/6/xGWrp0/bjKMBcDUjRIm2E7O8BiwQnjQAVvuI5wJ8+Rb1vifce+Y6PXAK5Y2SvG1xOlGB
1IRf52FVOhiC6UeOTbfWMsfnt+F9Fc95QRkUpKxyiHJXuo5NJ8+Fv2gNqxAjbH4exVY5thUToZIX
NGu/7PEbQE5PHIo0E1Ih6GY6xNmeMuLKVOBuMeqzcql6pS0JDQg+Mmlx1QaYd+smp/UEHRe2P4ia
7bs8MduYlZkfFI1irG+S6GrYbb3JI5gNjp5daRNejx9zPVCrA6CBeFxB17MC7iZpdKU32o5JAxAC
Yhfrak203tdlJH/z4Wd5dxETWXwSGtlw8m/dOLoyBrwc84SkZlehcN1klV/FSTCtBWikrDVEiCWS
8XZHis4GyhHvkOndyDtvDdjd2IxOT5D93SycyikD/UVKXkTUenSIiOXNa+tJTXzRvZptuvhoiyp5
IHY0rT1Ym9vWdKHShleS5K1oz9vSLWYelK3eajnlhGQO1jaBZGHJQjcbJPcX9ABDxB/t+4xugMRk
JPBjuYoDQ3qNXYMXY6ndfhqoLoTUfsrcYxQAL3Ny3PNUpDv8F32MLsF6MWf6pTeEJL/ObEl/fEdU
dN6MF9IJi4TTg5NnEP54QTa0SIWgu6MZE8uqvfOnC6k2NmvSM5n/617RkWKwqvZ9h+iTpCyuVvhZ
YSztAe4vCuxc4k5V3cL4uF1C2UCgU54rbD2GDer809H9QBTdtVh39FfjMGAAlBCVEwCoNVW9s6mY
fXjFTlLeTc0Im1834njHAcoJtHms+v4obqGV0NkfQPaN1fsr0J/AJohlGxHln3WGwGpVXzVSVvG4
3j5s2Bz8BtzqP1jPTYUdKZwcPuy7rod7WHviCod7GeGOIkN6mTE2Vv6G6wpWm9tIFcGnv4gBajbT
W8++S+7SroSVk/3VwgxnkASMGjCjZAye1jSrDVAj0WdNHGfyqlvndgPRPXp0NWxoOYoLY+QZ8rcd
LvCA+oC2An9gt/ePMQXqOG7WTdKVYJr7OZWZJqNjMgGukdQfSq/+GGODh0NZqyu7Ae0q640zt0IS
nYwBLXPwQgIgdc7UDlIjdxmMoUo7HFspE2wdQot+LQr4YNmat72VuDZvKESNJiItTqd1OOOx+AFP
V+qxTBrlz8PpCu1QT+RYFIVAmI86dpfpsRUmyIZu1KLVLpK5MB25aU8+Jw6w9iNvX8JunhCOMK8/
+KYE8vWt34T+1k9TCoWYd+VsFnc7sKjeZ9L6zC0ivhcTSV49nlfJ9w9uc9GdISIgESdk09CWLOJf
5Jks1iLHRVaxzRXEhIsO5bLXFtEhz3Nix5fOEqa11kWsFYcI31Dk690iMq3wF9VhnFIWml40PIU4
gpihCdV/PYzDgVn6A2QhFUuNtQMKQt7EnY7WdtMzdWurKtQAq2Kvi4x6ifNQ2wOjmszbLuoZKPBR
4youAAFLZjXj/06Pin4gSjLVzSQG/kStcuU8mwV5ngEycAXYdgppsk2oKxDIOX6zDdwwqdQSsvWn
K5tBj6rR53PP1LqxfaYbLZb2Tz6E26g5Mo4gkbOKdsO+sXbB9suzzfjo06Jt2iG7raCQQ94KFQ0V
qF+JoyNzTyz+Gv4ssQA2LvvPzyRUpiw6o4AzcENoBBcLmEX3EchbXsSoHtHSJPK6S0+BNG+9ll2r
2Gx0YVvfdlkUzCCS3mn29e9ZOusC9oNV6EjZa9qW9rgSY20TpRwdIY2MlhzIVOHKI1eyxokLTN+K
TZSytExwQ6Cc/ze5eQ53c7roRYTqbl7QjOQtr+a1eQVwogLOYMflhOkEebnsctFKJeP2yoRMVE/v
iGtma7MNVFetetUi25Aw+IbZ2T3NHk9E0k81teMy/m5RRMSqPfbKlfAMBLTVHjzGX7P01SpzR1zB
6m6YM1YizdBkXtse27gUl1gwamdO0qyAuB5xtADbU6YJuBDFooXtQJeshy/CxdNdIX9yMIweI4+y
QLvDJ6IpoV9YEYDmOPV4nlEBw1Gbn1oVWdD5/RqjZn8FJidIyZ4c9WOhOioiN1jc8UZ0AvYnkzr+
2kNVnjQHk9LXydwhtJSLH8zGDbHk0PS1CKsXdEvsApG1N1TUjiodHHLd+NunRRXU4MIX4BnhNCJv
km9tj8L9ubZgt4p8Ez9ESd019SJi53Y/hReGUiF2fVPi/q/hDYdV14b8MPqHBNx6wjO8syXB5wph
FDTFPKLPgC+4NE88zKN8+/pEkg5WAzvTEPsiLvWeXyNkGyHbyu3cSBQb5WECbQsXKlMCY2r9608U
m5OMvieoUcPKoJPMoSvKb0BxOZzSrkrGahN5Fy1tfeDb6ReWGDpbK7U6xEBL58MIgS+K5GHxHR2Y
9eg/O5WIUwaKVcgOtiWO/MkhKT1iDZAQHoX0tyBhKMN48kcN+V2YCe7NsVtu38q7uqkaboPxZJYK
mXdhz8gDxTste2Ary2FKz1Rju8J8mZOqWIpDj4rSUSY67jtCSSZLsOYFzyOx6og4luvGRoAxqChR
6iKzLeSPThu84vo2XumsAD0Q8G5K+YzjZhgZq4uTYxDr0AdCk1IQ6Ejnk5RhCS8ew9jAsLnA9miW
8nCHaYEVTWtTX8nZQhxgPxZKHYdHt2nuZUkacjVmM3s0e0U6fVzO2ZhewyrEHcFiNz2ECSadSxJM
WEM+M2/LbDhfellD1nnyOEl/Acq8tqQpDzpI9yQLv0rYi9ym3jU5RDKD6H6y+AY1lQPoREMoC4KR
jLpS6dvMWXfa6MtyV1swJ6Pm0gcLlGp8ab5Qfq1sdzxK0JZF86uPArv+wm2fbd9YVckUcKDEMbFB
UPlj2Vp5Aw//XXlVpIXHA4FTTEc2l+TRgILp2eNe340Gfzez6CM+I52UMmcN+tfuNeGf0mVZ5L7j
o2Kf2JtnS0qjX4DQVncFNbE9q9Ko8L3Vsk71kMgPETePAqUH0kly7veMrrS7hpVFSzTOLKXuNXYr
7wTYOA7u/AZT43sQhCClEMsn5J3Kq/tzblZ8zv5ATWSXtxqpEi/8+Cbv+K/sUOfsnhwI8FStcWj3
z6LltflgPhOzzwtcWCmPxM6kda55xo4yRdimNk5fXfgIXDo2mmMH/ShUuKETUdeuRdxLtPXECaYJ
Dywl0yuPgDvdCje4Qb8g244XLeHD9C5kXH5Ex8g+HY5Y64QcQj1knlj5udH9MBaNqpI2+gnoxCGF
NDGh2n3x1mayqcWx5wscR5Ew8DR81yjxdJCKO2ESKejCycpHP4bVELkM9oHg7vpYRmK9pPXwqFCm
q1n67m90HixL22BZ+uZZhhZoZx9M4x3Qo4K3g4gZ+2r6/bgse/ALRQSRQPetkSxvELSZ6SQuVl7C
2G2gogLpqdmjKOaqHgon7g78PdABoCiQA5qspVICvSdtUHie1Z8jGdCIBQM7HcmCN4mRlQvN1G2o
5lj1eGngajiQc3Z+GDPtNcxPLp2U40OAWodYmUJPJJDpAX3ksYd6H8VLbvS22iA7ux1xyZx2a6G7
M330A2r3WqqEWblG8T7sqKVBMhAqEDjzTCRM98JXWT3jlvcSwOiNllOHW473JpTIjjgb7JVTvKqF
XfogUzv9ejvEos2yriDDx0eEwkrOF/TPxYFbN6MqUxOnAxBGCgrPOJ2kO1Sbzks0vwLJ1nWXanLt
btPkuov7dLnOWt4j8s1X1eC60CoRUR8rOBaD6N3qo9Mpj7QzUJHUoPgqRVFuREffAi3XZeVmi7F8
L9p16jwbiRMZSZyIpaH4bBS1oZDbSOU7MS7t9Gc5OMhT4+gMQnjAqJpVO/N5IIgO29qZAUHTYe0f
8gHIBb86yZ33LbwpvZhzOVoJl9XkLwX9SXWMHmQELGvBSY5tQXoxBJO7q/h8tii+IHhS2jojop0/
fC2QvDVDjRqF9rrt7z7WaBw6eluZAyWT476A1R58aCCl/I+7DTp2CI0htJjslVHRffIEx+q+C+bi
5E0HVNQ6vYiat/0Zrx89qyWBF+uiE4BFneehgi5mZ7dfUdhuLZU6d8OLFOnIwM3RIISqQv7f9SvL
MadalQ6sGRY8Q9exUagG7Q4CyqKewLLUA3PdVIDGwiYpLOoqy0Em+NqRsps515nXdxD2CV7oMusV
S0UiO6gszZUos6aBe/9v8M8fZX+BW5SwqaBPgcfMr+V43nWYLAX2+CCcwxwJr690LWBOlJX1S7jT
VQ7lR1XAb4P/9cy8CloOKxN1i1UByUH11iInr+QWIZ4LV7p40Y4+WdyhEzTCufNNQntNBfXxEkAG
IcC6hQllUhnt5n0OmHRxoSgPxwqCjeX8elmXlJhpGcQ2eRcQxv8sw/PyTvsKWN+82uoQLavNUW9L
/F0uFg5cHeRAwAMGlRXHmTVIxy6Wm4qRJfK0yLNXTl8JjvrANSxAtmNVRt9OiU0e+hi7ze3+nHey
IIatUl1Wi7QTRMw6iDe6UJzF0TNDpdOAkT+G0w0AkYSrVOSJfP3rQfOI/QpauVrT0FdJSNthNU3j
0lEkuSb80fXKu2KwCJXNz4QiszVJ6ajXTsWazZTmcGFfie/NRWY7QLTvn0IrrOgXjyxp7phB4wNW
p0gaJiIBGs8on9/TTHS55aPctncZdY+ZwhBneC5MIOSYr94PxbXfGtSH7h0ZUtG5mrwi3GHQgLTj
UVkvfixupsPbuGolibWNmrs5BAbb6dnAsMLP0CEtEM+vHCsXNmUBZTYvcgIquh23rPc5crU9iG91
XgYQb2kP2PLHM0rTLb7RQsAN8v1rAB+kBQjjp9ARcGGWiIF+hLFMWGFyGf1qHzZFE+IqzdRDKfSb
HXMLORrKLgos6yNQHH1HxOl3cNV60JG3Qi0uLn1G8yeMBezWzSr648gDh1ZvN2DES4AdRSCTQh6L
DeRE2URtqc/3TBwksyDWOOJpLcvcnZAginqajPuaELyRIv148HfJTMfWalsT4UG86NpchPE3TvZj
mGLDd4FsFU9LSYP1rhCf3clkjwr5qxYtudNQv7kgtxDNG4mgl5oO5NcoawenG/gbrZQbiNo1sPmh
oAi5y8UOCGF8+dEowTZtNgik7BhnNeTiwAFT6Ar5TGP78EV+rNMfIe4aRZVMwK+nXgUSLZJ37RR3
CU8P0saMxvdOUgAzLrWb/gYvedsv+u8gUN679LPzImulRN1Jtwu1hFoKVEAAe5V+PfrCEU06T9ey
s1tU/CfvxrtRetKtImlhjALaPA6KURXzfjWBFQqsojWusk11Q8cDHMVHB5/POP1YlSXuRKX/yxi4
33LJ8hE0cC02QMG9BwIDo6UqM1E9kRb5CpgaTf9qVXiNzNyuE4gZYqoHREEzGml7Uu9+Tnl8/96B
aB1EBf6L4VJt1pMlNXyMdjr16vzjNEBIilv1fhMOM8jAFfIzT3GW3tKTNcypndzw+LJln66UiXgt
Nd3el2YIiQi8z0sRBGf8cyLy774BzFPpVa4aVUn0M9H5XhkXRAxvdJIWfdVjIdE7CHexOkimVT75
FCIBnmVpd+lWZ+oZ5VJcjzM/HapOMJuw0jFE/WDmDRUqFfftyOY8toRZXBdtMCH2bwDrGJNWD1Jw
dSKy6Bxn/LrBdeXIyGPDDIjsEtesdvHSjnyY9isW3SwS4pXT9aGziOOfx6F5ZohG+JainD+cmW6c
Gk+/Enfw2cbQTUJyAt2rLPEMrq8A/iL6hZInjD250Nrmt8f3f4PLTsr+JztW+NwTks/lETjk1F0y
EGuT2L3KdTNRs0cuGxBDL40sAPPLnNYJeZEo6Lwi+ULau5qLapjiygBVr9gIZtuVFP/3dTqAv13N
9l3WMIgcu0YKEcSAUdzh8l6FM+fP5ZIrOyc9QJASVapLNw+dAF+TNswAD3uz1EAbcR0HsEtnjfnT
YvMmiyEyO2NNdc/KF3qJVRcWF31ecp+2BmGlljrkWBjXYthaNPXQOXl7HhYdy6b9EpqCLuSNAblS
JGS+J7k/gdeZW9OQXRYOv97voewpBj1/8eQa5dKwUXVNg6pk66mKMqPGNKxwxFOQ1jD8/K/wgbMc
rEJiE+7uOnNNmbtXUUqKztoHuZDG/rdc+X7hS3ioauDHerI8ge/OUeLaOgf6IjdxQrPU8av+Pg/h
iEwV8Tk9t8XKjHwD8eBQnVrpx2UQNB2YG96Zm6FTUwXzhiXSzMpiKpn9mJhiUjuI/gTY+EP1rqBQ
8UY0trVAJ0HiIlNuCIZgjDUqyBBe6v3inTcyBqWmaBtzvRWZAWIvwfvX2EF2uGZZtYgQrSSazkSI
8pgo0WRRrEZHCoZtFfEXOcBFaaAXHYgc5kVkGzhvQOk2fOFgTW4ppvZlYvEi7FCl+EgUo1CyvOX2
xAggqppB705r3VBoZqMXjXEHFvepS/U3bJgak/35Umo0Esodc903iWN9NXim7yhwrAbdD3u+drth
8+RumH73jRAcv5+zuuV51/pSjdIACXzQgrz2roo1rIR3pOYeKg6zSxR//27b158zKZLbyJRCcXwS
ksvEFM5b9jWnnrsfTf3BAR9JCn1++yCpbFo4K4cSdY1kRksFpMqW12UdVmPlyTaWNP8pGzVj7sGH
OlSoWhb0zV+UZ4GFIMZrmbzDHhzzgBnP7g3eg1E4vAJazVADQaeRKlLgB2iRNw9SZyDDd2WEqt0v
oQPHI7hrp3wi1O5iwfgRqPXqp5CtEpG1AJBdgVGDH1iVQCQwAVYArTxv9HHXS4Y5iywoI6hhz/dB
ka10ZxDwnkxXb8MqDetOHy9jymK+uHnBO6H+5v4H4xLvXYcco3KpaKRvb1Wv9DbW0kr7rOuhsn/w
pdViQEQLYtXs4bJB1vIR+DGrpxbgZLsoGF9mR8Mcw5mI0ExdKx4coUfOsosME8lZuRVPy1s0sAk+
l6nFJWP+9iB72vHT7936BHNoXt3gYvcGAt/paOlG3siKeD+CzefLHEbUYLDxykddgad4B+CJ+R3u
JY/w8R8hK1QCvJxpUwX8ksPj4CNxf+svwRBYmI/xeJp5CtrbtXI9qHwNYGe44chGNSU4tvHFXrVx
tbb8/FYS/jtE0UUPrLrrzXOOwthvxkDks0dq+nQoT/zzmiPgpNJ9rWJWdkhCJ5yYE5f1PvuxZJBd
QQhY9eEhJO5jOLvQ7D+KEpazXiStpLl+ZIy+sG1/mWcQCexXAEipFXd/exnIWk6YUA59XtwnSf5L
9Rl2KpSXvrf+GnNma3bAR3UOqQtIswM/3eAh2WfCwjniIlg7hfUYa+a4G7JtehvSXNf58AWY/5v9
mjOdtMgkEoVAQG2H190mXu1tMd8oxRdKap0bwoScboOgGvVoxUN1PGS5G7Oz5Q1NkFoAQKJpyjx2
YA6Cdk5Kzsr7xxHnbALuUx29FHjy4KeYym1qeTdJSVuOcDnupXcFMrICiS/+qhyCNdv38n1EhkpF
/h0ojMVTkx6GtTmXnKmPMBCZuN6a965IHrofsUthceYXQ418Ere/hoC03GQoFRsjFIz/lO7gbHn9
vXNgdur7m8lSgwcWY3INBWXy5Bt6FkIYY9VKFEldgVHbdzGRoe4ZksfUcdI2JDY6X2LJVKGSHrvh
n3L54GYpQU3iDW7a70VjDVeFB00kXMzDGQ1KKBN7bTC1KqvILNaJ9A17suN8T3wchFygoaobXMpI
zewd32z6d/g0UzYsyjrzqCKBlPfgNLeDso3fsLYWsrFFpaHAGWkO0RrNa4bpaFXOdI/vYr0Cmd2u
0MixSxbbda8VYnnQCx5BlQOi+xmvfGlBEYoJQE7dEhIPXPMyH3KJKCkc+eqXcmZI9f31wVfKRVgy
nX3niPOB+e+bd91MHtPpJ/zqa35qGOOYxNMcYOirU0cbbuAYByYOLrdxg3QI7YPiKiMNrwmOLq4V
cbfXZYeu3NmkrIRfDJVi7A8pV0G49bYtc7vnfa1qXBWkM3RFzpcSewf6LAmBAvzWtlVwcfUnMpRH
g9SPR6A8Fv93KJdS45KtuuLP3XRpd8uRHr4hG+7shaFM4vJ94i4tZm4OmuHGEC3kBWbGi8qtS58U
lmfGFUd13tLb9MNYbZKAajTMb/KBfF8IG7nr/4IBFoSNQhzDl90N1E/E3v05PNx+GDbdhY2Gvrq4
/sbduBI2KTqI7Qzclh55KhbNxY7If7U1/Oet0nGUGqoo9QUEjIb91HbzmUpstCj6DlqXBh+7HtZ0
zsDhvwIHmhi9uebHKlRTPiZtZXmdDe/GdxFYrFBFIgjCr+JFgPe7RKm/IKWUz24vBlAui+IGc8hp
pkyx/v/p9rk+D6uOm0kA1MEWfzZ6cSMXUNFkJekg+YR5mMkJvRq4hztLzX5HkgdQYfHyaiYnZ/NY
KbGvpXhLiNn0neCL+5LPV80/5Moun0aIpoCSEppj6gMYQ+Q3Px5wxKOUl4T0xKYY/ssgHnJyEBg7
/jBTNDVey3InCsg4JkO4/Gz8bhIBwu3srYDUCtTjqwtbdrH7OGSn8PMhiQzN/pCbQ+Trx5rMPWMI
86eopfxlEVYXWZ69g+3z80WjIF6Opj6F2ITyUY40dkyGSvhn9URHgMmajdgvdOxUEOBNIU5SpwXM
V6JoQbZSr3IX5hVCBze5ouS+/fKkA9Eo5WlcXil9V96Blq9rsoPfvq41gURGxhmJBVmxN+ZDv9gC
NJdVQ97o/tM1/lPCCn3hoSFcEWBnObsJmMUQghfPhPINyK9FbnxST0HNInTo1fRXN68TG41WMDK3
CpIE2y5e3nVMPTzHu9zpdjErbbhzVYqR5fl1xbRoPsQC1jHQGK5vWPRgTctNehHprYckLqUCwJYK
8EsmgJt55ZhieLrEWpcFGauEumz09PwNYlT5MhocAdeeY7jqvLj5zwuZk9X8k4D+CuBrcwhCQ0CP
l+B8Ez7toxwV0IfsUBvMaR67eMkCVAADB+gy2EuBe5RLoHSwc+YUxlDDH7FYAW7nBH7lF3yJ57Hp
QhIFGbyWSmR/KhnakfmFDVqxuExnaOSdYMSs74hC5kWl16KMhEpvyi2KpeD936IY657zgitTu43b
5p9001OYsOmDtNBYZg7LNIVbnJn5UyqCD6f457KskA2kSIawCiU7Y8RLekVGzPCk6IG4CFubtFmF
i1kcIluBYulyrGcuuL5mPtP5IDhhrQ8dVG55Cb9Z4pD86WxvAYqqosKVyd48OIzTcNE5q6XkzWfD
bSq4js9R55xuwsImYD/ytTIaRjR3nbdOgedpJzR08ZtyzfMM0DIYZim9bTrNDNxRTsD4f3231AAp
d3emCr1xtkrQI2wZjQlPoh2fExTQG7Gq2as0piB1uMUVki18290UlYyHK48QI8YylsInK+CQn6nr
ep07CiMn5dA75WZnTZQGjRoJIQf3iUdnDoh+hTLdPWJrA4Ke6n3rgGBFzDd1Bdmv6OYrDIVYWrdN
xo9GlWQu9+d3r0fljvq309uQlNdQLfQFYyboiB/prCr88gLuxt0w0rYbG/v2FzgVAPSPSnYmQDFA
wmP3V7hzbLIz249HURzXxuuTqgg4/4iovawt+F8OiCrJJz8q5BQam+SRsszRq2SzLcDdCoPZSFb9
CLtY+AjFvaICs/31/KHEbzdDMfnK69WTS62u/OiSWa0/QDwwcf+/6KoY4/2J68INfyRR5/34csBZ
wdZGZaRtkVwIkHlux5ki9QSEHKa+Rj4WCqjgLlsFSIf7tTZdKeq0RrsDQOT4EAx7oG1Ja9VQNsdL
3nIcS50c522cFipfQtK3XmwTt7FpBnigstAB12UmYDTR2OOUfjLW1KIzOrsqivjS8R/NC01Bj6bE
u+duhYpvwDIlipvMf3PGWwG/fGvT44xVtHiu9KyKif5D6bDqwq25cWqKjHOCjfw9PWZ1+Gtw2IBN
l+iQ7J8QPTXEaIvOlr4jGCp2EpkHDvhSXGJwuC2FniWehn3e1+7HgHFPFZBuU3x2b92xJQqm3Pfd
bFmR7H3ZQx9v7VXc/iDgTwh5vjqUDfEWfDvju8tkpwFPC50aSOZUgSPRr9Tx9frJGjG1MPjftSsQ
CW1ugsANxWRUNxePYECeXIGaFwrhIJAhiDPVblgWRFJKlQvTc3/RDGZ2ReXHv/w2HWRDVk2XNkCF
T4Jv1xnWZ7fE3m3wX2+mzSZleTOtYTwXRl2T3cLN6GrVH2UesFkRxlpk+vromvxzzm50ZS7oVnDC
G0UZ+ek1hjV8/L2YcIWk2ieGwgKpvq+fQEe1IDAenTdJv23Cg+2fZYWSo6ZF5jeWmZC9qkEGRI7d
e171hm4euIdhPeJq/upMctlsFMXDoOmiJ2HNEHdtAqoin6YSIc1n6hKFdYTih+Is06ImwHCJUJMn
iS9azeVi+6CR6nIIEqx/aPIy0AXY+0LVqPSSqtsbh8T3JNl3YM/TeTgAA+EMSMTNiCd960P5ilBZ
NmkVf5KF5LTEXdVRQUwa93L/YsLvW+BS9rwYGOnHZaaiMk6Ph8DmWKfAH6KvQgT3o3EkDMuEgieG
aRI8f0sVJrMWWjGw8Iyu/OKpLI+pSwFhTeu3fum70Id5qB+0zlbzDfBGaC/oL8v95Tc9M7UPPZiK
AE043F6AxSJMMeWMsSHO8QLUgDr9qqR3mohNbEdkfCOJzFmrT51zNdL1r14Pwk4PreriONHP0dts
aKNzT5PJHyumBRpuw8A7OnosnqOdxxLubmybVryws3z7VwnhxxLqItx7X+ihH7V7z5Jx1iQxC3C+
gV3jGRSRSL/Kdu5skkIyBVhF8YLV/f+2ziVfjhy+9/mTvOlvjzbNdrHXzdxASRKUJ7rdKoZhF+zd
KabXq5GhPVyiqQOrZsB/V+IKWEUW7I4+Lc0m/5nMuAkH2J2/otVxKB2ecIolX0LrU+0efD4CuC6z
5c2t9tew5MSMwU5oJXaTdd9kRqyDGIEPRzgh0ELOzBZT0dkt5glCRMytFLp4ibYw2831xomLV8/a
VEGh5jziRl/GJrpfJV0+1+kiwp8Yk8Dn+yYstn728TRLITP3KDAVbBmDb+VOzE01Q2o28dLtm7/t
PMnuR7LtMbvcAK8X7Rz3Rel75DHlVbwFPBgqu/q5oD6bL+QhQ9L4sw9wVrBvX+i3uSm9Q2bQPqQ8
wS/veYdQZ5W86Ln7VUUdG8l0GOdJOi7MD1bGYjfyYYQWjQjRQE3AYjjlQUwznoSmCd+5nfYppwVF
fpwBcN4w4U8eq7tSReEeFf7OMU7umY2JzujNNzk/L/5BVZpoLnWoz5MMukXmDiIDNGVNDqF9B+/P
SHcP8t/oVQj2tZyyGJ8Hk1oCb77Gz7zVoRwa/7MCzVkBvl5xk4UC8x+KMnfe6VY9YpdbrQG9WCLl
Fj4svm3UyeWAK0ysE2971mWSJBs46tCCz3LzNO6I1uf5paBS5iLoQSdW35x1cuED79qFfNGyAxZJ
Zvd9BPSTK7CG1mVRihU7wZueuJZ6yCFI1XADyUs6M1sIhuVkfiIto87e2pQrBtK0sk4ipAMDFMGT
C1ncZzcUdWQxCAE8wGIHALGpUZNqKSU6b9xxMnqveFPf+w8CVG981EylrHm2wapTGMcHV3gPE+af
KRR4h9gJAkQBxH0RYQ8PvdkGpCT9Pbsq6bD3m6oylsRzICpCOksOOlw48CsIuPugFCXmN5ws1pba
eBJwUo4pLtF9GbVYwwy7YeBS5UYpczoVwZqklmOyC+MiVG1mQ7c0GzdzITqJaT9GSMTu0LN/X/Bm
SfLULiBoMktpPatr3xR9OSr37Y1RqNYaJrxvntAGcT9t+yOaRIHAiKHM2TUbPLkrp8CgPxmfoQIv
9P0+zg1JG10kz58Mc5XvoHNV2zJdZnn1+7PM9wqadOHKIKQKJ78KOURSBFQdFxrNNwhKyCed1LSA
6gxZ27RgOtVmC+7vTfuxR43ezdSU62UDTLJJoGbbUI9+gMT6y3XdFR/MxsCqAFFZy+NBGqR+RFnV
rjtkasgrpUZRc05gy2ZW0og4635pvfRVEss72ANQ359tjFln0o5jRNiBhAzSaqOuieSlyF2hX0XD
P7TnbUNO7pserdt+E0A1+/fyIixFPxL/0s1tQmZK4UOghgjS9ZDczxZIPPRaUU/YGE1/KFLY8nYm
zBBUZSGWq45MXbYRwVugwKSXBc6XlCC8woW/98KWK32Py2PSdZfbrPM/ZXoNXb/oRptVd0IWzjov
bepVk5nSKC/UZWKXeSrEIdiLzflorGJYA55RJPprlT5xDQjgpG5QGtIUwSZv8MkIhCscVFd9lotI
ePeVxG03+9kGW1iJlfo688Zh+KwTEH3WnASBSjbzDDAjRRSiA9EyY7tDGmETIEYTmGS+4Kf1qVF0
xNX91sHfg7F8QuPAZbVNi2ML8no5lt+hORX/isEQlG57KmhvX9MbV4Klb7RayIQj38Pwpvnb6G1S
hopRPKADpzkb4WFc3yyVSp1TgLysCUI4S5PS/q3gzD+geRepXfn0LM9SjruRFH21A2QKViaYgcH2
esWIduICX2jw80yWKFQI1n4Pa1A4n5WGtY8lSPcnU+/Ab5wZ8kf+88o6tVhUh7g5GvNGSjlSxjPB
MdDA9Izbat6P9LGZMzbK5cMeREOzdD0b7wIKx+FXtnj3yPGvHHsPO1k+2PGPjf0mA6eDfJmjjhKR
yJAI21GwSxCbDTx0ISPAX3Lyr0Q1X8L2scM4lX/GAyNiIcNd62xg0ZYYiGuripY2Yva3Bb24OJQV
WltKyYr5Nqpyh854eET7kI06DzSB93kKPJDd5uTAH8zP6Y4qWpvAVcUNx36oYnkYtPvhY1aae6MD
Liy+0lqYO5zrM8HAcQ7M9gk0e6nE4HD/IpFs1PKQdT9/zF4Vd9N4JInGIAfglFsRncg6CSgOKPti
tvGJfJ8ybGqq8DeczbE4BEXRUxnHv1oEetx9ZIR1Ld694//zaviegIXiB39Ab32zRvB3HFQWxRlm
rVArJjU+AOdlnT1tqxK7ON4jlmBxjIrlLHYfdiUqQZlD/ZDX8XTkgrGieyb3i45lTqAqdY6WC2IW
j2UyiHG7kEqE44dijjknRzRw4+BGO73K1yPF1NmW2M7LMvDr9coPVG8w76i9QvMRHdi1ZaBH4+fM
7/gbAz1H1YbHl+9FlxateBUlfPTiHCuk3/aknLA8dbfJT0IRbw1eRUXSqHidqpOahyBpjk3zZxV8
bDux8V/c1q0qjnIoDBrE2ts9NDHUz8sTz7QpjqywWd22Q3oIrRJyaqhWNpVl9HP23OWhqXhwzcjo
n0i8koAaomqsjq973Z2efVg/Cmy94Sa4s6qFhBmxXEKYPb0JYHLHK7jEq2ATm2gCdRWCphl8TYcD
g4ZdYbxlOXAbfimpNyeOSUdGAe+3sX73GdD7VBkAuELhw/46QUK1LbWwn6Jhuu/kX67wY+g8t6xz
U/40X0OagqJJKR/aB9ZHPi12XwtGB7PT2o0ma5PxwMK/wUH6xSsAhVpsF4fMgjyqqhQN951YUU5T
zHw5DANDLHLyOlxArdCINaOXX5c4am/87ecc9mYDQM9m30+ngB0UHA+TYeF7utRYkrU/nlHRpipy
oGaj5Oda/AxunzrDi0ctcrocTWsWVdSkEDnnl/xqohesntNax5YxpYZCZU1Mxqod0oelVyWJBIes
cCs927JsXzRu1U4NSUjQYSFpGbs2Vil/uv/sROWChEmcMwZGPFUSJIVOwaR8hnay7W6s3bX6/mzP
YAgKmJXt2Ex1WCa47q7W38m914y3S/EP+3hPj5bG/w7Pqa/cu+0yCl/p7rRHQgHQVQCR5atah8Wd
UxGJMC1gcIy064+sHTNKGVqjIUmClG1AzKobc9+gWY1A6lEV6dNTkl5n3zDNm76EL7hglE70JnFd
j/KsiGd6oA/+I4RSzqI0O2nVOkSSYpGMhNHginUgkMZiBbc1PByxe+8wgJJa2QqoAj7nAJcG7iNb
P9yxhJzZ2Dr09zWjfiMc4qv/TcoaA8OFNBpDWIa6o/LQrBWcfMj8DGZmtbbg86EAk35u8ndkZgrH
IH4LKHZLBqrTp/xJaAaWW5cZFXSl5gCU6uBSLFzuY5cl+rbxg5Ya19WOb8eAMGXrI17tX4/ec6WZ
7EiK1W/rTZfVjGdqOugVewnkkLGfrO19oyZ9h3veNyfsxdNaQgLBpoKh40mG7d4YegQeDLQzC8jx
sBdgN4f9lCWAtwGLc6Z5VmcyHWDLK5lcJv3Sgu0EmUYFdmyKZf3lf7JAgTFdIo6Q7EjzQCkLhyvv
fWlRLH4x1ItrRt3AxJqReCyN0fpV8sjyZ13Fng2zitnAr4fxnXxDXDazwynhng6P5tu+9+Xw63T1
hgeEdCLncSaSrlSz59qi7fuYo7Z73UG9FsT/9cn1iOZK31WEFzfYuHO89uAIiZD1nAt+vHRmvPMf
YNFwtt92zz07xOQM+R3ejoysv66Mt5db248DFm8ZxrxMcIbLZfhlLYR/bMxUFW/RmKVSHAbMgYcF
O4K4SiFaw0VWxahIfobuH49wxFrAvR33dPV5qar44vYO/d944s9LSZN/P/mU9/4fEQPYR0r6SxTZ
FTMZVT9JQ0X5eoKofA7DGjDjRi3MBdP/imKyU5kTADhI9YpYr4uZ6y7Rn28C8dUlpaH2MhBw+uc8
KBYkZ1Ezm//9uthHB9CbBMWygDBVnhTNdnBaEaLkgAhTsiaPpxDNHHUaWaD8ESKyZVZtFy2s5eMb
VLXFaMKoq9jUAKmcUS5d7A966ndVcJkcuoGhBUV8qQmjnwjA16YGNdPXHrerqt3xqL2/OnReVYFw
D4gm8fVXLa+YFfL4JJ0T9AjcFnVNsrElOteY+k9ls97f0ykcNuQlFbFcSNXsPXM6RpQ9+1W9I89g
vdrKz4uwNOgHY/oQqaOoxxlknT65oRc4uxKbv8bQhKaJCmyn4RTNEQoYvEI43izZ4pghEgIv3r+5
fXcN0wYsyoKDKw0PuGwhHc3X9VrvGTcubck4lbaW/fc0hZvjzZ21w1FtvKPRjao5m61LgKTnxcPk
+wlharqKrW7YC6Wt5Hr2JO2OyRqcUJe7WQNLeXLh+Uq6+SBrvmmWK0B/V7wsnR7de3P7/wl+hj7m
N2lyfvfeFCaL5fDjqJxGVGRGkdULAXamIO+s0OACJzIpBVZpcHxvISj8VUr2Qho5a/HIYOp61aC+
gen9nPT6pceMBN7YL1mFsRR+/Un4ky1MG+rtyO/oxn84U3lqMRWIFo7WL9+QOdiEHhCWNEVbqs45
5TFW4uf5UuPtldAVwrQvlYEnM1Nj8Bexr1UvOVCHrKnDrpK6So+/LptkhxGQxbnfms0ssQRusElU
BgmeVyguyiG4IjzI5IWdBt/9PdRUl2aVzNOoADzFoJoA/cTC797+liKG1uBdVOZp92J9ZbYNSdDV
RYVqHn9ANn4ZKZ4/2vsBjqENXXBbgP1pVL0brOkiKIADSIr7cczGV48hKz5o4M8FzeLwp9A8bScC
XfLzg5Utv+d40oHhiaENc8+LcfYab4aoshkTZfjNHzdQmugmeGf9u4ExGYBosLFLTQsknwL9k6HP
MCiyXr8EA84T+a09G0aHhrHJOBm2VPJ2qEycMqEELzM+YrKz6OeVHIFLFuE3IAecJpIsRh/kxEfg
eKl39tlL/rLfoyRH98q6mCMhJBAOBNuui1R1bQlGIS9zrm3kVl5IHud7ZKBfIx6Ql6GqMsyzSX8h
K0kjyb6N/J3flAIOnzGiRHzZ5fd2YRUqof1e85TxxPPbHTMPFinOYh2dlxqoiLW37cHjVekjlUYk
qoVA47YvVYxsqTt2G5NDGO0lzHiK3vQWwLvXLKzdLpxCyLMXOPF1nKE2wXyYpPulHoFJR4E/HtoN
OtaKpc9Pe0pOlBlpC2RUZcC6+428ASt/80CVejbzkGPs8lPgjm8GW8JO4xbsU+x3XsC4z9QvcTye
BSPgzgX9YA7brIWUEO7QMageH7rfzy1z8IE2gOOv165nCdfBSyNOAH3aJtWRYs7HlllvPTmmNhBU
U6mX6DFb3315RLz26PVfSar3xqHYjIWJD22d3JqP+pkf3Dn2FNyPRTs7t2lvuZdKdauXePTy7ZMp
SeDE5rUONqXZ/9YcIQFjdmPs6zMNfAByDgpnaZu3GpDSqKc2uA1+bGLEbShySjvrDS8H8E8oYdK3
af17eiL/lSAB3kUgjJGNW+tfu96NWrwmx0Y4rI1wcg/7NpxsfNWlui9F2hUdyUk3uT8dbGX/utMl
zt+5zxU/HD9MCvDk9uOdxHsgMakzEs08XDFfrtBo0UzGIpq4052GnNx1kofK4RMMWmOVcMN7aqfo
jSzIMxPMge0TZi0hDyQG89Ln0c9BD/f+uvpGH1Dhdyto1ok5wsX9Ue/MKiIv95aYPprJ70pgYmq1
Ayhz7P7Re0E5/dof4RowhvHZEwcVbI147rqbk1Zo8SUXRxI+1mymxiutwbXwEGXeVLZRqjMOhKSf
DhPrsDwSzRMTa8Cu0r8wGXb3d/CeADuEujTWLh46bNuCZri2iiy940qcqdNUNWtWCGTnQpn2m+HK
h4CdkEEheYd62iii29dF4IZ2lm8qabMa4s5g4+DYrd6KThqNRHfbeozGg77ilzR7CLjDjXEd3XgL
ttvLp1lD9i6jI4YC53DBmYV3MHE2kfcUty5r+s0Sp/bZjnFLRRXuWh5bNWjUG4bbH5wCWPA3rTIT
zKJbjUNOSxUTT/ZmfiW13CMQA3vBrqXts/VISmPFfvxpBsUVpc+8Ni0aN1uVl6FaaVqmAXdDoF5b
MRMKdnvoLEFuBr8pwwNAJOLJ9fT8+VKME36XdkS9X0ByP/RKtR0VX5y1sKlYQC2RN5E9cGERjLIW
tarl0pdpU0HIkTs1UqW3a81d1blbhrxV3XKd8tqTI/gyrLRtoZfcxYA9uPfmH0EYyeJK9piRokMd
rvRtI4qKjYTEeWxLc24u/RadzhglE+UK7FVVuukZjFtQzWZeyDstpWVLbiDwr1iOJQU7s3BAFBEn
GAGnl6ptB1oL5UUvdx75QPh+C+nR6uy/fkDwoStrX9qwN0o7QD1hwEzD62WKG/xNpVlwK+8L2Sw1
o48R9111z3IbGjeA4auqWJLd83z9JVMCQ5T3nHVov47FfdgT38Qf36HWv5DBCGgSyPZFSrUwPS50
UjLNbmT4vDMM41fiAN0ab05Yr03GccxZq/Us1CVgECR665m7wib2klpq5SVfwhiDGPddxR++n/ae
Myup0SOGByrHhrM95P86aRRhU1YVrv3LIS1JebmlKDeVH/I2B90HtDCxDhSaACFRPfojKRt1vN3L
vAhXD4eFpTdoWg6u668lAjhFq6SrHYfz4dgVQygFTXCUplBs2z28skcEFyyJs1GHVj4jTOmcVv/+
TH12bvLm4v86s5CS42ZecHUAFVpO0nY0n9pnwiF/12PalEMCbHBFmOlb9uGEP8xfwnMZ5Xkb5tQx
MJfpuIyFTPe7CVbdhRG3k6pZtyNQ9eLQrkeoklha8r7Aq+0Ox9D1qLKmH3do1OOJI3gg3UYi7zlZ
+jDDORLRruXKjchQ1kQMKxb8g/2qJiFmksfOGAffU4nguayU2o4MU+GUvU7bWBDPWcHR2kZkyW9S
i8kYfVNTt4QoSCFZbhuKLSTb68+j2W+9ACSs4q6OCk7kqMQg4Y7ovqnZsWgrRiKetsvZi0fB7ZeJ
xHK1RweK98Gh9zBNx6fgfE/V/8O9ai+L8QNYn/yxnLEncEBP6syet1LORw3zk5ZIepXLH1iiwWYW
yJ3qECT0qzeMZq2n1unCP1tWPrNvcIe4y/MXY2pi5S2p0M2gacrdbF1YNRNagmW8n2HvddqZhXcZ
n3cRM6OEYDVMYf8ag4rjuGe45XU6m/iH1wb9HKrvp5xEv+CrG9DvJ7vWasYgeFD1aM6sqsTtl3HO
lvYjRbFwyLTPUuvk6DtEFFyyZfFsCx3hI5XpjIqBoo5FQWnZH8uvlOvY16bCREpQME11XZbejQ2d
k5UFbNR1O3hr//aAk6ZpVA9BICAwwti8ylKUG39UdbyPip4VHsZWazXuIEj/QsYcx1LLcWoV6LrC
L9cmjEOYwTzQuM5qBA7ulvBc71xXQUijyLG6TUZ91leL6DQmHLNtX/LGoUimLH5gLrE8Xoy558Js
znskYlXZ4js/QtvyNqEbDXgOGU0XLH4Y2dcA3rg5X1evCoI8TEstKsrsjjJ7xNTwCnK57vQhOELm
rTzaPCQYEBbAn2eUjJFTIwKquGoXCJzhaskFV+6yWRvmpds+aNq3wxcch3s64WHEMYRsLtj23dk3
lgRMEBMcrOmgj5xVOjzPWEaze++rn8uIO7mokxmTjPpjn/pVS9ZL3LYjvjNklTH65KHwdZydPa4R
FfSgnELdnvetQD3kGD1DRz+Zh8PosupPA7NIF/P1M2isAcVc5NNaDHr9RpTlJb9+gxoyuF71JXqC
BGUTW/27c+SvOM1YyyRHcteoLzbLzMXB7Uhttlopnysl8lj3oaFeX38FE8kFPyQVkvRLZ6f9OGxg
3AAx/4CQ8dxtTDKIB1jSXhjmONtrxaRdCnM+wOoUCoSQQmN7xgtl7ckKOqbLjciRW7jFPOws8y68
4mnwmpCwaFia3vRE67+QZvJMcfxB08pEI+NjNJGFt0YMW5EDw5/nB43K42YKxA7xSLxIS3RgD441
7ifak1k3ZuoufveAlRyr1EBOyxhKFERtK0/FMucfza0OdgiXW3blo8LKBSWS1k1dEaUCkyZcJtwS
HIn36KinM8Pc6+tHc+BgzpLl71Jpyzu502iRrGSHZ30zP0CfJ9ebB3jt0/XJvlw7IuNn3E5AhbV/
4153CmAv0L33Iok9GJWNzGewf/FX/nOQQ7o2hnk7o+wJTayFq+YALdFW4WAOazd9QMKEFeC3M4SS
PV217a+ieIiaRg9AbDeNXV4wWaXO4zqisupRyiAxpZFykUjFEUvlIpdtbGpZ/5hxCsYy8ygdZaUy
uSvPLA72ZYcPeqfBdgJhF5k5V1PUHag4sBROtHGAq32piksDvPONU5eDkAckPmN2rcsaQOCcy+3R
u3KfNqzmyKAacjbPoNxbZxC+q2xr4P5abbNzrSR9zvI9WYJ+K/Wljmp8RDW6bFKezduGRIM4HNaf
Xwr4EVCk8wcTuDePqjEWE1qQp6owUkAF/y8ZRRMlmaj5I1U63z5nVrs7i6z50tUq81tZ5HJqjc6L
Y4GZGk/wV7oc1mgYgaxKE20dQUxlCdHgLrRdsfFiSKckleyvmHKdI+1ZWwqfp5l1nqXAzJcNh8ik
fcN3WHcB1cAflm3JEg8WKk5QNFlWeaoqXcsi+yFWA2H9SXPztqvcinYqYaO4395Al0gODvJLLMcD
MbZRvZRgsX5ZzFXj0m14EwdFomRZt1Sv8jJ2hXMfoaFbKa6r1sapVvF9fu7BRMGSZMMPT9tu7riz
BoMUAbzNqiMbE76BlKP23lfQ0c//LoRREGuensvrDgtAyzrdgjDxUXAqHRwJpH3NLDe24UMctOpu
l4q1oq9i1A5LY5vxaUqGBgua1N54c98Cblprg2OfMTtfPEpkhSFNtkiB7X3tphUDtxvgiHDh9uXA
pdLJ40xt4PAD3zGhbabfqoTFLCLxcxxCTQ9uz5cMN/ONmh4JBOsbyJf1LMvq7GeMM7vlnD6gi4vW
zvKRWyHrA87xA+FP/qs2ksi1lap5MiSwEYUsPOqKwRcLB0fU1HVpUrlZdxY7PCecmGFRZ879PE8B
I4Bh7VMbKFP4klIMRK01VY2AZfVdpWuO0gxs8nlLSGTdeBDb2ab4vqxoiIX44/XHJAcVu7ZetWGu
n384M6/5ggQ1RYgUoYMkJAaSLWK6gFYPfTl2goAaqRhIUWHnvBDlCgs96POpmaSYYPesijuNpl6P
x6BSnfu7AxcJaa8u4egpxmUi+ARROygrs6WDXwoWzIKbtigSRCOu3aTG4vPMFYUQfukbG8AeNEFh
S5algNm3ReHrD/EOuUqsiA/bSaEEwxzDfJjhJiqplFotG5iWdSP6V69wRaEdDppPk5f90Hg9jI6z
AYqcP0aJ4cjhSgyAfa9qe3BF6OBOtXin1f4rzpgyOYcZS7BDUzpqGw6txD2oEu3lLpBJ8Kr2sN4e
mUpfia7TzRSzfsex/oa3x8esBdHNniHj4+c64UNWPoFVkUh3DsDRrLoJkDLlF06ypQrbX46aO0Or
+T52WO+xLj5Wg40ikMZ14RCY+0KsSPv67pEV2u1uf2v0dtytOGrNo1gnSxl0WxDTxuHoi+8fBISS
JT4uf0x/3O6cxoFy1Z0hDkdymNCxBIKZxRgc9agPpGipka+Wxg/kULpObVPcJThs9684Dj3We4Ud
DVY6v6vYyFsZtlN6dblcWW5QPObCr2onKZnlpbqsArb6wGip/MyUP1tspSrM8WeAIK4MPRqGrj8F
J5cgfx4Th9vaNHnphl6P3qmu56cd8Z+/gsOIfxHuRgCW34ReTkntnq0HapkzjEN6JoQfBsjoty5v
KbFvMj0ku+XukSnWdf/4mWTb5W/koAYtdyvPhkujrJWJRmfsAseXzMqA+hMApwB6QfoSm43PcrxL
3+vAbik4rOkJdfaDgdYlVsllkDCEyOe4nz4slPkhPFqaXOJqen2EG0XcMyXvknBjiq1ulBW4DePB
MtdkpLKDU15V5MMxFy+68chcWb/xhoBzf91/qv3vYBvLf0qeLJYx5+iRTcaf9MtzECQoD6dXK5Wk
/Y0U/ervnXw8tth3sdaaIhOIvKBg4Y3WMYghJW0tK9Y7SF9Iv7WUts61Xxf1gLOHfjs5chxB92Kn
7E1Fq/rCwVh7Mf5PZeVQOIivjD7IHB37eGiSKqEwypehG0w3GAN7Fx1iMaHvyCgxt5NyW5GetVbU
qAuVNv7oQmaGWAF8BBp/tnRyvAEfF5K8njoUK2c3gXPhd2PMsWUbnuXXFR7T4Ofo4tkSQ0crBkLn
ePLqgWnD55Vs9+Wi+kOQm5yPnU2kw41WiyvwHCgcA7KrRrkqfKyZ8S1eKBl6wyVFcYtBaUQQuuD7
Br1c02iXUlQkwEsBEhLP5VsuU6JVmYsMLnafBrGTF+pMCfrkOAbPpfgtu6+YOkEaKG73WKRURyYT
8+E+KqsQXo/P1FDF3xB6N+AI4p0kiZhELQj2iwTZ3Sv/81ZCYF0zbESpQZXfhwgyyC2VuNvjWDl+
KBhPPwisWCemqas2IyJxyzQX2gXwktvlTRwIkHdICdiGjrcShS9fiXVCWUpcKY8T6OawGz4YI1Ci
1BNi+KkZDgZg59BzgOrDfWTjswqwJnyYhNYZ/536tSP9a8D4QG8S5QoGGViR1ltBLf9RsjQJHeMu
YLSVX6ieSZOx0misqZkOQs26Zu8ZbYUTsawb/evVLj2xvvOtAbZg8cH/wl+T9A8yiU88S+Mz6ovb
aofqHW3k+h6C2jAX5s3Yz+L0/TW9c64pN0FYwBvIzOL1qlktwkgjWhe98072HCrrE8lv4gipuINh
XAx58zrLpGRN94jnzS7p8iYlIhoOBi5SUhwC5+VOGH5AG0w3hadJuwNYNzDxKxpdvqM+FNitPW2z
lgPRPSkUH7sHlnaDvd1fY6WO/zbucXJEjFFgSaP8KJPnoN+f3OiuHDLxQD3V4bRum4XAyxouXEQY
C3LPx4HKpIdFv5AUT2OZj0PKIzJmKjEMbXgBDfkUV9cou/l6v9GpsMS37qIJie2Kx9w2U/opj8Df
mghqNC9m4f1IuaC8M5oLgDO05BgNXKpBN3LHkEiscZvL/6ySQyB+2aGsDe6B6Axo/LA5MPgBHPcW
l/d93ZawogHFP5oxHQzQme4Gei+JbIGO4CzaH96e7j9f4gLLc0jw5RuD8/oGUMHvYG2pNrEW7BC5
+PSperdlueGJtHfPmT0uwkuNAZkPXHOlSg6J9dwpV2wrQePRv7h0ZmOgydoqsB0w7aI32xLBN0YL
QJSvwysexd7HW24CFd6M2wFkGPP96NY/h7UfVqRIKJjtzey1LRBK35uyTSUSfpn/TLghrzsdWtvE
UnN2QN33m3IO9pq0us2486nH5o8y7RIqBO9t88z+RGuD2bnxwzEP4KmHIz4d2lAVufdneBcQq7wK
aqbBi4llIprxASdZqFypeZqEE66chWOPiD2qg5fwtUqvwvSa07v6/fLGPF+EN153vgtFdRFWY6Ra
NfV+FmNc9tyfzr/He2g6qad8Aw9UL6RSWpvgjL4lsNY+NT94Gv/KHzvhrd2IygDxzUj7Sbk6Kaub
PkPBmfCOng1KB/nxlb1ey9I+v4m6Ja6NX/Vb5XV1kJy8N4/lEOS8kav+z6pSCbLTJ1jXCcU5uwuJ
fBP4f7GotCx3T1Z7tKDu26eHPn32G32KLJAiGs1WCY0vr9AYuk+vclWmAxyBJd7KMbeGSk0IDino
G31iRF1TpFQ9J9FdHg/vpWQW2A6lfDzeBr8QkWXSAz1G7AbrXCy33Q7mHMse86Ej4Ha+OldGhIiO
BDbZwqbI4smE045x/sR/5wKRH5LU6EVTZB8PLS98XICR6uu2reQgwmu/9t701qGX88hTPJCcJrdt
X1S1+SAuSBuZ6VlKzU+swqI6KW25RX2VwhUkq6vjyUwz92HtrVhvi6kayQg8hg5nO7hty+QvjZYu
YQlC42sFhiPC8cDxH9HHdVxSor9M4R4YHFN0DYclafOJaPJYQMD+AD1ewl2v1mn/BGHDAkKlZFZ9
AoEDSdKm9W5Z6hb+ywrUhCYQV9uuUKUP1jc8mnH8O0jsZtSnqp3XC78DtYNbVijAtoC0S9N5gu/b
VAtPzdzWjjGcc2vH4FGYbI4uCwTn7AzpG+4NshW6RYtVG/+2DtA6eYXdW8jD+nmG2UgsRu5g7doN
xbxb5Tm/hzqB+wvATQlWEFUAkTTGuXjq2vimpTz0hphPvA7Vxv6agC7VV0DzvBS4ufmkWNEuSRP7
ZT1IAVk9MkqpBxIQ7xL4TiNAvs7DMAi7XKKy6ivZXWbVBthxTS01KW5M0GxAS3x1m7461tqdV0xe
qrDARC4RuAB42NYNJPjZqj8qU3eqmg0kPr/GRfs6ZFvG+1KYt6/guqT2PVYX+RyrOdE0xaZsYBBG
SaCJROD1ynlPJ7xCLKioEUx9cdeVLvKd7lUt2Yn/5TPnJOcr42uqBMxi/ZKSs8w6rmms9RvUOdBY
Un9WFYl/VfgObk40nzxe/k6sQHkiFl1VvEyNt2Pcc8dtglHbt7ZDDoZkm3nezZShqWkNrXHcGVjl
j3wi6TWc6kRsg5+KYl38/jZbCzqfLx5E18ksVlIhp9zemuQtxe0bLNvoqjiWCtpFpo6p+GaDBoIw
FqIVXa6zX51XGcr5sHxvgJAb7M21CZFNzz+wgPzXktdXTQ8tpCU10RBICEPxSANEqrXPw++2I+l1
lZcQTQIZY6z16oNYpAZDpXSw24P9KuD29VsaQxXBjYy9D3caYAfvxQdaCr6UfMm/EDzA+tUN4juM
L+uzVMR0bQQLjpDnE1gbBm/dbcZ0WgpoB05noUg4krFo2V4UlASc+g0yJFcSnTw4RHVt0O0v6bpJ
94XQ1cok2bXXtmI/AWMerkl0o97bMNSjBIOepYQfmOq3khf/wo6HSL05CgvQlPEjoHbF8iGUp2A5
8eO/52Y/ni3zCUVEBIzZEWCtG6O5c+MSBVzUBquwizM33dPnIjm0noLoJeuF8lY7h7z4McUBJ6p9
396Cc3XLPyZGtOZ1wMAL+I/PPpc//iziIQd6uNFOZ3baheK0dzb9y1zbzq0fkNw4NCZVevlBu+XN
IIuil5ApFf2JKrb9UjhDPUWCOAzO0JbrIMpsb0yBfJaKKMq6WJliG2HgHzkUP4854/yazT6qDs9k
u32ogSgguI09qeoMD0JtYf5qyvdADoYHVsnRKaOGNn2oTMr1hz7JZpE7VodluoC5OD54uCqI2qHD
9JwnY32S/WsHLtf+EIFQefZrvQtmJihdm2OxjKWxNlKDRxT6/HRAUCh9nspTqJY/CFUF260CCxPL
F3XD86G308KvLEs7BKqxMACNTctO491nQVZ/iuGi3OMzsLC4AM53GPXHxW9LTX3wxfmsudXN+Eab
5JpDnLWU8lgkW//voe7VqE8v1dhl6AJkcBjInAqsurgzU3thF15NvTWEGE3KsbvQ1vRQyOMPfVWt
Fh/3Ug9s2BCTeQVZWdSj33Kz/zgDFA3Gn6d1NA1lcDmM6AK8t2IakbQ8wlwojavP/2ZQuijvRNyi
D5ZdFZDC7COMti+Vdc6LTSdP7mq3aC1DjuhejXIVaoJyhvewJ8octndqTr5VA7xctsJmhjxa4EwK
7mQcVaBEGO8PpZNzNoPLoGIFY9duix+rhMqJhg2FajMvCWKJm3DXOKeapfQ5QTMwqVRGu1+UGnes
AEeKEdaZsqQu0gvItN3BzVp1EO33QVawbbQqpreAjbPgQaYiBnC6H/mQtF1f+RzrbFabMbgJujUp
F1FEzwXcevvD4A0M7RPPE+Oe9IEG71ghhQs3DNUzu8mO8krex8h1aS8kbSG1GIt8ufDXt90UIySy
w4gnDWrUkOVdYEMR3tDPS/SRCzM64YIYLkyI0dxJiV2Tq4A10TpXAaZ+lCZteNPy6D1yHCf5dkqu
JW0Zmfems9NC+f2adw3GnX1fF7hfizoKUP7a5vvlT5gLJR70lMn5UxrObkDBfKdPQdpE5OlrKBgD
Dj7GABPveddzTprPsWUCeZxN62sC7nUDkSjXrsEbSEwvwmDskJJgbMLKtvaZ77dFtoyHO55zblr7
Fcq+sM631RJbRke+GMCfMrM1JyJ9N5CusGledJpf9gA3PJbZb77umnxmBw/cu43vNq64r3qyzI7X
PS91srxl7IxrOXb3Hiv7l4kRdnQwKqf/+uvvHd7q64AO+Ev1PsP2HptQgDHjdM/pECBTZVm5HpX+
aMd4PTT8S1XB49YFGN11lunAo17druNRCqY2t5D7ThsJM+GNdS4wmMRCO8dca5/bMlqP1Ae0HEa3
ANAyvY4enaNGtS5tTKeXC1ruZIdXy8HY0tZH4seTWpmJFVD+iVDwYZeSrodzxkqgVlV8yV5MlIti
oibhtp2F07O1xb2Wt+c1PQP844MHIiSLAAzyLeSCip60xSka3/Mexf/SpXTrFK4jd+LnCInq0RoL
UyRd/NGvXKkzktgigC6lUm73YFPG/ZtWDkL2/Zo+z5dNxziwhKzNsZD//ds+DjP0CXTwKqX5MqPb
Ln3/YHqbPD9VgPOhCsPt0wDUQNUBpu4Qxm5ZBANZwsIHVLY6Fxnx7oTpOMtWY8oP0f4V+UVYYPey
0F9Qwlv8wR8A6lY+tc2wpCdxt6XHi+V0vtf9vJ/puJdq+wz8F/Fauhzapch+QF/rNfbZP0YYSjl2
3NFvsVzIqiqndE9Sphs2tIu5Xwt1JVMhWTcwQ5onKD1pchUsVyPCw2bok3zi0PjOEhNEoj/G5O4h
ylSFOBj8I9x7rT+mveAplxo1Q7L/umm6KgDE1RNk09v3XxJnfENvA5PInZOK1X0Kyb8ePO0y4aH/
O79g7R6T3ov6OTQC/aN4R2KuNy+7yA13phR61Otewx/+ofHCjPYj5hyZ95qL+b2rRSuFHaXv6cSK
2oc0NOHuhotB0Vsr1+BbSA5PcoLMFWGZgeAn6dbuWyqzUGpUp3pMvqrtDDoMXYyoQjrWx+1POpNM
AJEqdEX9zKKDDjyQGvI7z7/w4FCPjlgUg2vr716EdEQ7QSwS7NG/n2zLrZfVHAtnbxgMsqY1oxZK
n9f2mge3yE2Mw3F1NSLFemS5hgP8erGqEDu1sOlxde9Fa7q8yYMy62CZV6+dnr5+rB9k0bN3J6iD
gAPTg/K0glO8/PTjn73FTVgQf8pQ/GFJDdQmzlbdWcwcMpMaR+S4/pIEOSgakc63K2/xUxBfP3Qz
CRBYHG+j5kUbGs7ZtXENhzKd5FKVIezFzz4AcQrr3+cI/6bzBqI6hpZiCO9NKMqAQAQoAYSH6qsO
truWdCv7AM4Zxj7w2/gVQgYkgkJ1Reif1Xp2zKJH/+0hAnxXOcKEif5CmYAQE0hOcdI27gCm3eU1
l3YfgrtYWszXv41xwJurUbhiUbq9jGShrtDN7gYhJI+y1Lw2WGiFfCgm/E5DNPOBTV3AkY8KmVwO
QsZ/H+qJgOq5tvg97YDLYiCmhXhl/9cEd4M4niZVSrGBEmqwjBPNdKtSJWrsdO7xaPoz9nviDe0k
9Xcwdh/7uhohgqoHwSO5LAEqmuY2nk2SjlkuxxZ3ru9SrjIYnujY3NgW6Mvqp3ZWmpuxWthPxOmK
gil1gnUlhDiX+U3p1GSZaHADv01eHMskYzHJsQqeVc50ScW4khRmQkQZz8jvI39gKpyRY6Nnv/+b
Z63mvw6nqHck45WlTNFuebOnbRkzjnceS0fGG0i7ZFfmcaogZCM5sSwlzAatKWsMCiZ4jNrzAUL1
lweZSqx1Cn35UNaj4Xo8OY8giu5pbgULS+pADnlcNTHlT9OAcQBGzBTQoy4wpMBha6bT6e/xIDHQ
ibTzCpiKb2irY2f3cMZQ+Yc0Los+Rt5nebfQeXWeGiIbOC7RsiYlJR4W2ZGcMa4pRphZycExQsYA
oV3CUnoJWsUlNDcAWhRaWO5g8DeFjYL2pbiLRbpWuOdVi7TIl3ue9T38NSx1tgHx+CepNtTqxx52
5FZuDmVLUZvhdMUl2KJ0pdtcvYh8KZTfLve8iR4ouQSLgCcLWWskPN86LXNZ/mYVVEz6DI4bK6Ni
Em4cTPAmcTbJMbwQhpNGw5ljPNxu1EvgkZIl/kuLA5rlscV9sBeBDcflF5BmEs2Hpu5LmoaE3n8w
U6HPpGuyRKOEC8VmNpU9BU3zaPzD79H3ZOxHRHZ/UznsOGRTSdcffKK3AfxroNUt7pMEIiVcEyYE
IAa3ce4Q0OGb7T1aXUc6oLSKpedStO0/twiBSqXMpYH+hj5S52DFgw5vG7N+cMiCvKsOTOv39Tgt
dLS8JE4DqKQAx1mKhJUsq5u1OGN8BYFlw+rf23KmF8fjKDuHbcxnVtnECPgeUdaYM4ZECLUPcyCm
s6ueh+obGTjoG8ef/BaLiEc+VRzm418UrV6WvHO+cx6LK+ls1Ltk12QtWIamhI/6t2OEAA89Rzti
tAwRhlGgNcIrV8g4MCDKv8pvCkFL5NSIqQ3L//ZTNGv54FPFP7+iyptdDoqamDk/pB9Bn2uOBzdq
ByWVGftqGbh27K2YNR2GRLhEANKGtVRkgj0AiqnPptcYAhGMXd3ZOdXQniMBUcjtN6moURtFTZPg
sbXNsoTbKgoA5OhkpXm0g14kroe3U0H8D1lRp8Bg3QMM3WuPhGizT6mCX1Bk9xkfOnoGmr0tE+M3
Scce+BSLDb0LAaNkXrbHXhf0ajuIbbC5aJP3m/HdjBhsWJLEWFrwmZDvln5MXJ/lhShgCZB0klG7
UCKgZM8EZQW0IOIzAomMhZ7p7a511d3EZ5IyzUf1XFNivosS4vjMgEC7ZnAP1e7u0A7OygfkRl8s
z1+tb0+t2GM3xgJNdJOi8Vcs1udRZpOp9K0f6/F4tYeYeZBm2yQFitmBNTPiHLsLsTcBySFhtnLT
oNsY0M9igcXBoTeH5zw8QkYgr+RaTz04mSS72ga9I+XvDqUMTCoZ2tjJNwCBNsJxHzbHUcVgnjQP
5l/EJ91ufwVb1LHalIYAvnJ52DuUm0wn42S+JdIFP8bGR9SyJeg/l9hqfcuvUvoQlOMzxZu2e9k0
YPSJV0t37q5biufJMtDR9Cn8p3+IWm/CoGMva0dP0+Pf9QTvajlZJZXocXBH/BEKb1XUrLysUdab
Aj3Py7N+ybcoG0iK94fj0wbjc9NN8tm7evT0UxG6i9F6+YvTe7hJXgKvOvRtXtIzBjYjdgDtCYiW
VodDUXq2xEI/pBCILHqTPgUTrFs803LLKugJeRImzBeMPfKmdNQmqrhCHG2PbawEsp24mO3gaCRL
6jfu0JJrDwbJZxEbabG/uoEQOp61A1kB9SWzpeoz8neoMZzUjSj+Gh8+vrfESJKGdqIPp0ZuMvaI
SE00oZo5L+QdxbsO7eISC+xNstGVT8INTJjAqZQkXbxZFf4DSKXaiyj3iT0X6+z4fbTF6AF0NCLJ
i/P27N6zuTX14Y4hGJM/YozMWl9KX+HLZulR5KO3Ln2LT12asMqsRa/VqS2aUszK3XfXnMxdcTRF
0/DJTMzm68ykd+hHWL+61h4BgLlET+VoD45Bmqs7b45197rJnbetpZnx6XivJBFKhCB+WCDSEmMC
1AWYxae/RR2C1NbE55DfdFYHMJ08VcDI/ny0hkWM0PKDXxI41E2JrXvk49SDo/jfKCrCZfgNooL4
HOU7zLB6sa5foTNNv8DyfBBPPkWB0hrZpG3fzH/ErtZ8a8NrSvGYBBdpOrpW8FUy1c3zINXB+q2f
X32PlDUKesm03cJ3/BKb2jWyzwkddQGS629Sg73xouLWAX12NpEfXaj1HN8Po+xtpdrFC0CDKfJa
0ou403St8i8VElQdMDu0arl0SJleV01SFzP93kC0Sc50mJ28sF7rpTDChQP5POWz4iEAqSInvN8Y
EO1osO+90hjcAtZwYvPjLLfgCkARYoTM8aGLsEpy70Mt+A3iviV8MBIG3ke+P88Kok0kPNngCRwt
HD5jbQx/CyWCQt5oxUccKXNeq2ejXV408wBsOlF4Je7eq1jIVWzHVU9NZIo53LgGO87O/Dj3KkvP
vChPJVjoDGLk+ATbqlZDE0oIRyTMYp+ClQCeFqLbHub/3Sb7xWCJQTZUC1uWEZ0vfcwJwA8fc7jz
mpfIeuRwwuGODNrfz09H1ovRgQC44s10w1Et08igBVxai9DH1ztGggdSdc45z3VzcL+BessNSULs
ZIrck+sGOSDJTkbk7djKyZ2xEStC3nJ7Gq1E0m3svUjHJt36ZsHk/QIL1fXyVErxG5FBvIi3GG/Q
2tck0OV7JkSNoXA0cT0GjGiJWfezwADrDHijoaXWT0eUD80q4vcjdYROKKNdax5pjTcAPIBe1O1i
X0rcmsufyEWJzl2KemyQSOaCEGGk4ZM125VuCdAiUFEMuhjBHDPDcy6a+E/VEekNzGOUWEsl34yA
b1U8Pzfsh5+aCGbrP8U0zuu783Rdl49XY1AUyK6R90I+cMyWPL8BAD9F1x3pbTpTyuH6VaxncrNC
pd6HboSq/msYQGFWMAN+3Dmcfn0KU/4JyB9GWKL5VAlJGwUQ9nCjpJk/6Jtpyhe17sFnGdfOnygT
rBAms5y+dhfSxmntLos6ccg+2FpzbwdRcyauKznBbk6hHy6vI6kZbpcORxfggcYMaNydKZJ+472P
Zu3bePlBOmMyj+ssdGriJtAflp9BDF8UrpdBjtiw6Yany2ZRTEQoCDot9UCPj+FP3YvR7aSeiM1P
0VGtaNqd2FnhY/1gmmag2rVd2TkJHRbiLpV9ju5TLZDcSlvfo3ArNZD+ANXE7BCVTaoefBZtQtCV
OUNSQgUPxoqLo7PO5R/3ooFs5ax09bVBPSYRpLZD4tTojxRYV8tLnKo6YY0efbexm7nlQ0q6hDSG
XcdLn0NlYkSsTTMxsrjKZuKKLJsMoLw1lEL4L0Okwebu/gujEw3Hh0u0a2lCga+uuOtiAtXV2Tr3
/p5PqwRPVxLtJuROgi6lf5HjzhYE5V6w4jWi074oCZhUDk7Pa3EyLKJzyLiHVqKtN1vZtKA1ICyV
PdJJbeaWSJqNGEXdYmFZJjnQcuNkcMfSj7BNCL7Qbu+d7r99TZlXgwg5AQQJsOykTgPpildRFdqv
UByhq+xqYvyFlVAtNeFjkByo1RD9HsB0J3mvjDm4rElchSabvGC20H0aOyZ2GUvi883PDHmQGrUh
fkrZii8ET5/I7Vr6kFgM2fhZAFaN1VuNW75kDtb+2jg0R6lCg9+egEOh9WdN+rHQ7pifSYJ4vGTd
3trNX5p+BR5D0VO54nelPRQ3Ea7kFPLrgxMIZ66H1leSHPFzGfX1InJwZnG2UoYaD5zjrXBxO14h
KhGshKQdOWuZlT2bHTdjCbbnh/H3kdEdJdnxbmAWjfBfO0jPFV4RyyYYIsjZNXZ9JwswX3mBftm1
4eNwXVB33NJGVjAJJravJZ3a94oYyh7cN4zlOWB7CPeiuhei4CF0ZInQC4J1CFpydN0onitu7PP0
gltAvyjPlqwKE6p503KUHshfiNvw/TXsKJ2taXE6/l4JdvXXyyWW3bnWm2d1bS1OFc6U1bknAi0v
3kQjRjgXjpZoZ17pR0fKx39y3CuOZV/SHoOHhTzty0pBanIT3LSE7CpWd2YpYGtsevMjnVMeySmA
e7I4nQ33BBR3775TvHXNm2xO5BoiGR1h1T7C12LXKnGu2JVvC1dv0X5tPxI17HI1rLsDRfqRrWue
arhomfEu7GHlJz8fBktQUnFApOZphz4XkSOmajCET7liotdVNfKCdxfDRobBzCviOanvWvFnutP/
56TMIAoXcY59Apqc568ae7/mTC8SB2yq0XtECeLBXN6DIgzkWtFtboVQsUSdLvPSjm65xPb74wc5
IsySVi7V6Z/9Eq9LZT8XTVc9b1XMvHITtkVUiPg2APfwkf5tMMJYY+WuoeUNcBNK9/P79ah2Wv6C
CSFYpqGe3xx+sWDP6dK2iH89RXM0gTyUyF5rUsebCvV6yhsKDPJCVYJEvWONg7HxgC4UPa7lXU8b
kEHWupeI8wvPQA6fwCsu+TB5/UCoWyHWlLUpddN73lu8gyGud84C4aYKWi1eDY16j/Whk5pLpe9R
XQj/dzVC91N05cyGIF5V82rT7o/uB/j+QbKKxPl0Si4zpCbXPtCtUDVG7V6SAdToqBsJ3UnGbUqF
X9AM/4yZ/AE/eG8+oiCNhPzsKV295GHbJd8qsQc122Jrof1MomZTZFJYsJuJqE07xMP+XqscgP9u
nSQD3IzTFU878W+K2jqu3PbjZ3yHFpRNPn1gttPxpJ3hax31Kzan7mglUypBEWlc1NoXxxHGXlTO
VNGoj/V5YVIY+zTSjlAfL37x7dsVmbrdkxHs9SxGD76CoCmCTMThTqbAV6FYzsupPe5diucAwYRr
8eJF9IFXA4hMyB7pCyFPphTNlyrUq8scYSpkFyJGVS5QdQgBWkHIoqEJn4jiAUwDmPZ93kFFnIK5
DkGDkWVagA8uM+fQatzgiiW+Zc8kGa4CuxrYA7VYLXtnGNE4ilL70w9h93gV1MxZTGLn2xE/P+U8
JDIN1x5qoLx9SVxQ3v9+oIaFXl6r6tl/0YJWcAbzilc69PibTGrkFBaLv2ivTtZn8Tfxh6nnUxRt
DtLyOYC2NJCeCNRpBurEYBrUY1dpcEkDpzNP4neSc43xv+MsvI7L5quEngbNeqmteq51oOGn42Ff
8jBOKkKBmmlJj+62gsLtvdZXP2xVAWJTfbSVAL5rL9KYLPB/voDRSQeE79WwjQYM4QCsM+U4+3+i
UPSkgKm9PulDoZ7QObolJhQpTBIPwTZjGkhYVeH5V18RMOor1E3Ye/YOdFG0dzxfklWSGfsGNeIY
I5qD/L9ixW0x06Cs8btobwf67/G+p1BiSg6rLZYwFMKycDDj40AUvlBjSAjwPSDwQZ1QIxk/dRzE
gEDVRewJf1tWuuzoNOI4xC0XoVCcAk3P6yps/DsQv5Jr6C3VD3V42lgQNHddX2vgs46eNqElYe10
VN/1jbZCMMvQvP6dFzsB+rgEL3G8VZZpxJtWn7v+0V2KoBTzsOiqA8tJj1vb+FnY3DlK6NxOSDay
64uNgQiLaxEiG/80WeM4ogxpfAE4ZDLKKSxdIxlffigEJghXQz/U9UHlCqVdk1SK3D2+HWvJcwk4
/HN5aUXP/K7uHxBHAISbIrlZbmdwct293WPn05LDtsu44GDmO+7J2oszgSX04GpCBaM30TuI6eKB
zVJDMQ9KUppQ/ASg3GEhu+2fp6Hc9h+uM5Jvlk5gJhViim9Di9v3jb5P7iAffoZ+cR8C2QNKvZeg
N0Kp6YlBOEYNyOWpb1fhaiPBRGutz7GYWAEUyy3E1iKmVXsmMmISnUBOVILsJv3Pcer8BertvF/H
dNEWKk8RHhcaugpMcYnmGMq3nMin5q6AZxqpEA86hpQu6ht82mCO4ZJhJ4cKiVFRhise6PhFoFZj
fChKJO8L4Ur1mhWHI6QfO0xlpqRkoNN7aeWgm68Yq1D7PlqFi26n4KrhxJJwgkis73piGcQlmdyX
HS4M+ExQ/9gUdT+T2AGAkTVvfikFhu3VO4d2oEewxW4P0wbgAT+FukLpoZHSF2Fx7a0QQrm3hvLj
4MOL3OH7VWmIbA3NG/6LswwAn7OGX4wawGxkq5+6CERdFYw0uDhIyjt6QdrthMlBEwcNAsWLf35A
qTaHizla2qXRnfwG9Z/Sm6AYXgUQGoJi9BsSkwPQroDNYhkVOp21OWgK1zvK3IrfMrJcOmlm1bj0
8M1K5aHPmihbK3tRoI3EuUrFqeKGxBT6KgTgGNgOiYPxfG1++Q///wrRGgzLueH1/WK1c6plUnM+
BqqfE++QOe6o1ZTQhdFd1GYXC2eZeAI5B0zPY45dOJkGe4x3fxsgD6FdbstVXyYQm/BkAC8puOiP
7z38PJO4GcpJAYI+axC2AkvGM3ceXyLng/gGn6Cgwark++hjf/UfK80ZztNa8p5lYeG8asfwEQzZ
aXrPB9+fAbdRqt6ScYUwXpALVoRcbkaER5bmbaVHJQxiTppX/+KToSkAYnhiuH6U963wS6YqU+dD
nQjlMc7PCrSADd9ZBBoQ2dplt0Rj6ku41gJB0ttKMiVCQHrbUK5pK+43ZR+FRX6MMzJXSyGD/mLF
X8UAkOXxy8lvQ2vxubnSkeLpXjoBrmEHYerkcGoUz3CfeukfI8J0r3mQ0ugNLOFyoTbdq9c7CAfT
TWwAXZzdhu696zvUiRAR+UrNlFtG+2wSFmgjCR1d+OVW2mhizp71Pt7oAatXZBirSvbdxmcUAcsV
mB4pELfvLNPmshiIk1UPQDtHslEC6nOzNirilFJ13szDrL+9IeApQumWWz5CilpdYWUh+fgBaDGJ
M+sS0t0r9cFTe5xCTQkcbtqXJ+qI32WuhzRk7OQ5C6d/xg9rwElRq4La2zQZ13rIEmdGWWE1I4CS
Joof0ALzdQGR+kwJPNYuI7Uqzw48RKWJcM3HIYfHa1VsD3n8xxiiqrHj6ED4iLSv4Oh0jdMuAptq
wJGRt2eUzT4TzPQEeDcwfUdwtQCA5Ob8wL0I13TBPa00aXh6wvDDVrJvfH9BLqL1u0moMwGNcST0
uX/3xXpQn28a/GThofIpoq9in6Pd9+sMSjd1J6vjiuV49koGxag/I1mDAPnN7qDjRqgm0XbVA/6b
1AHtBP9xgU0Am42msgFjbxH3IFpsF9RLMzboP58a8cuuiMArIOVbM2QQpPYJLpo2E6lvsrgYeh+i
eADzqmt3k8WM5+Rq1NJZ6GMcIzycGnjew5KOIC3YI28IAS7f4Xv4DyLlbAckLYxRP9I/saurYvvx
Pu+qsgriVzJrMpv+H7fBWxGd7MX++fF0ohYfhEsL5lGY9JIp9uB/8ltosL8KgXrJT0UrmqAMmQND
iBU4FcHQH7FG6BmzUSLD1MGLksxzqiikIIndMcI03NU84kn7tazaNcJCq7sd82qr+Fm5UcUGLA7T
SkSN6S9PW5nd4y8YZtVCamn8FbMsJI8nnV5UxQmxuQO3Hh6+ixdrFanytznqgYrbGBGpZSP+Hl+0
KYqJNTsFvDnOM1Nf81cb27QLm1xcoBAGNymwt0ZpPUSWx5U6nCr2/OZ/bfFEL9F2ygijs3h0xC/Q
1ycK3fGYAyJVmBvxMNbPIuXoNwJqeYYwTVAY4395XpmSMh2aJqta/xhvDxA5hv1X9W1+nDjdHFYS
sTOMbGx5Q772fTIbhLw/1rmoThRSAxLfdrdwTySwwmqEnF8NWI+sEKKdWMCFQQink2NHI0WuWv3J
AAs4NctP1di7qEUMcwiZModsZd6R7o6ALsLVPnAM3hjqJozK2fYRKZ+0wVo4xO+IKr8Jt2oO6YDY
OOJ7uKjwRPAQlAPlq8WQYxZt+bCx0oVu4iUS7Qeia3mtFFKXVw/xWsz59+FikMgbtm6rRajOaM/6
jScex8ezFUPoFTMP61WgrClzBTCzQU6MSdJH6WlFJzpcVt7EQtw+Zyu8SYBgSMszS2eJ9QUhUX6/
wn3Wy3eY89AX2VvzRcZ0yCEinEWWTNV/EpCKyAauCvtXr7UZHu7pbWd2kNGa663jlvlwMyNd1E1p
V4oKnCCQw47Khvhiej6yeZBxMdDl2Jqt9RH7TwxzGVHiK/GUwQKkdO85CfI0uzkZam5DXenNNyyL
uVWkW3xPAW1nHv7agZLL/FIzfHr7yLyfS57V244pAaGVdP+5zJJYoOSkcUNS5RvkP5Li3UbYvSeW
EDJgZIaHpcF5zk4PaW2Z4PHtSokD3pfWOJO8w32JnYLMb6pm6vTmmhQ5ZhFswGReCsJmhEN6Xe+1
+roe4Q1hTp+uTRihlQIJx8OpntclNz+/4Z0rn396qlA8kgYocNT6r6vpB0be3xhDJF3UUyQl4+R6
oACNWg9bAGzj5CUST0fWcnuj4vBjXfl7USJFicpHfPcBRKlqtn23kNAp10St0Oo9ephrKrhiz5/T
/xAHZndIY/C75Q7o0N7YAiXsHXB9mXYsgOoV35+wyhVFPFy5PJXjP+xtCcz+Z93JP3CMkXEm0vmB
mS5/UdOzTisbBxMFjpWvBkqhkbWAEgtD4Z36VS0YSao6SmxUHcF6zhI1Qap63O1z2kUqL7u+Bkl6
u8ZxYJOF6c+woDc0HsYLirO1dBpHfmlHaMptAz62gfoNWCnTnho1o1OEIJeEFPUggyINo3Yt8pct
Hc9HxS/EDlvTHlFQ1Hr4n3VOFar0ccTy9fD+WHuyEvUh08JFs6sdK5an/H8nTUgA1Gr08/EXPxDo
3K6B6Iy+dWFHI8SIuKDJWMa4OjcSAnKi8L56EuloRZcjGA3VSNlXqNZ+5rO1E5v3dQ1pzQHsjP2m
AX632XT4mghkVxSiMZZ49Z7YyQHfIolYPDL8pkSGA5+8eNtXtSpnwUYSsIEmZ0tbEAteZodWBHXu
xAjqBHkNO5Yf+9SvviQWnIsNFgcIAULcPCBITh5oyGq46+50DY9/JFcge2FYIupUYwD1HDANeU6Q
r6Qc+/NJwnoJKHmHnNP7++TraOdwzUgSqDK0ybuH5bjGSHxGqSaGEbFFrlKHQrVjCQULWB3stI1j
HtqgII2uVCdnba3hZ9VZDBI2td/eJRI9mGyefySlrc+D3kq8tdn6Q/8d9o8zKJ0MBYVbp0aYoFgx
ICqVpSkCuG9McHP497AxLh61PUqu6sYBUaF/jFBGIBDjZQq2JScQulNzzstFZRf0delAYaGcqW6c
CAwLGCAuagVjBBvrleb1AGI0n8+o8qPP4XIFKrc3P0yFwEh/nfcl1nwzbjZ3vLoZz972EF2jcWpp
QMzQ7IocASLn6K7S/NYVZIIXBeDs2hefNaJjqadAs1iQasjEJHBeqKe/WXs12/Np1sn5rVIHdbji
/tyy/N0Vxgc8LxMxU92fMXkCxtmMdea/1SUOijrgm5wjNuwdHawcKJ40B4GN77FtzCsChyN1tbCI
oVC57gPY/041Gp6IcgeIJjxWpSZLwqWoJLBrdGSGpNL67hirDvZ4QCVZpwa6D518U6ZAWRyhMkwi
ySjFmQMgNZbrzH7IxTWHpNAg0P0EPQjJY56sLC9Gv66bAP8Z7v45AMk3QrpX7KGnwYJ/tM5vGcXF
vcra7QnyVc32sDu95AeQl7afU4kDYTnjcw7Fx4lAVKiogdxcxOgGWty15Qe6n8AIMS2pdcx+ZQmQ
oRlS3hLZREL9w3QCGZIw+AVQNu/TaZmx9V2dBdDuciDtvfZehcobNWRRFTO2Mm7G2bSS2Xaf8+K7
2FwhlRjTY5PYLcWrjSvrmNe7y8vv9TXHruL47V9ublLIDVok0hgK7yApS1FwzCtwlUICn54L16Bn
s+RWwGqSNgr+sh2e2TI+5RVL8S7vdVJqxbjQVDHsWIQUg9T3vhmUNUVrc4XPoxBnz9Fmua6/dxX0
7bwhuWDdAlqUWkaMvcuwUC2FzNTQSkjzwvvTG0AzCETUfPfDFk9jncbj3Dlb4YfTIh9vRIF07eaw
2zQYpodjVOg7V6BXdJZ7oBx2N79RSjNRpFytVYiyuiUiXG+XW1spU/pOIY2o3V1f4HLM352s+/Je
8WSbkPk6Xj0h1Hwkmgyn5DlF1Xw3yO3WQ8MSjLj+U16YZfpW8VhXMLp6x1C8NwMyBM4B35s0ggIw
5ClITl+jt4NYsFl1+iy/+qzQpSRZJRv7+NIzDWM7RspEQcR5PaS3tdPbBNUUZZstUXUD4o0CpSzt
wtoCE9f16HpJo61/G6PKLEXHVVMFQKDeHIxxhQY7wm2J8ufMvMa95PywVCX1QBeJI1sdAOzs9T+A
MxRerCq7DpNxyWkbO68Id5nCW7wqQOp3W6t3xTrNhFb02IRsIP+wLKUl3e9uoQxBU7ypLc1mUYSZ
jLeQYrFfv/744Q9ftuAkJ1pIeBm8QlPRapQSnYhps3jnrfzzpdDRN39rOOIKApWj3pNPiAvXiJIT
42RbeSyLgJuQxbUl2PZUl0SDhkbaBfwkFLONyWNGk+KLU/1PxA+8v4gtr91ZxbNV7078p4/MoATr
JAnRrdafRxFp5oKNIPxYcJVdY42zdTsIjeOKdHe7s5jXRFejR9+kRgcd+8Tz9JlAJYLX7zVtxRH4
L9wVfWn/0MWP1tbiL8/3brka140mdjlXNJ7p8q9XEg9xpq5vNg6GtFGahSv08WgPbzmiYnNdsteE
gqJQkdiRJomc6V29btdBAfC1WiH0fDobnwxXC50jx6Wx/WzFPgOA1siUopaMLjs44h+F3aVI1PpB
Zqd/faNADmdVPdu8USVq3LYNHhpVTwu/GmPx8IckZGmSwNhz+ytLu8TJtWY4f5utlTKHXo3frQw9
lKoa+AQM6M6d6KSAg8x8JnR0s6H9k7sI2MDmrxX5mqrB55DMWhyYjgAM0XC+e0rTVaxGskJfhj16
OZokdiveTYwQ/cd6ciPRRVxfDHzk+OsGcZmEBZ7tMaCm8aeYtF2YX/9mOhVHrU6B2F9gZb7GNvtE
OlfULapwv7m2IGJIGcWAxB10LJHwVS/qfU1TTjqkEbhlp2JAuTo9QDwiemxT0jE7e3BoSEokG/tV
Lkf5FNuXkBDJEOLND14A4NRaiVGQns+nnPdCdMUaBjVvtDp5fKDjtlhHbm1CWoHNiJ8HqzRPAg8j
c46bLSte628IeQJE8rBnwbqdhDV9EwBeYpUuAeqvzLJUCHOEf3ME5UICLWh+54reXKZs4IR5UqDc
JsVsorynVShOU6QXA3ac3nzAtSEx1N+1HvAcG+JHbQf5zz2TtqHQ5xerbJqCDzdlxtg6IMbFEI+k
PcGAp3E0eo8fl4dk5ZpfvS7TNPa9EilBj7k0zVGwyMMnD5qI0981+oq3sZl3tRX4Z6fsDRy0Lt3v
arKws1nuWSf74vNO8VZaPImq9W8Yj3GlTExKBljUnvjSyfQqESsyBa92tt0zStePoEw6KFWkr6uR
qnrthzOmpGD0DgpE8+gHAZBksQiMMF9C8RagwlBTvGYYQtaCLlvtOwn2vfPkp0NrEliwLjph5XH/
MU/AK0QauZ+kp0F+J2A/STiY8unJ0UJsuJbWylAP+KppjUYyHlzQ1wodSxcNT/b2GMwFolJU4zpy
HIDGol6hGr0eWWRi4uvhGb3430Obzifsw2PfQfrLvyyKf5o+8nZ8U3DgGguSSpR1j00I3hWRxpzg
S2fEJjzSJvbBkjmCJOe5abM8RgWOlyf+p/qWv9uYsPs2ABv3SacsF980wtjnG3bwt6ySIJA5TfsO
W3xx/8JGkNf1xdUsPTWkbdAZT6aOc7J/ppdcg5kYw55QdRAcWB67ZlCJL+2YaFP3i8gcodtt2d1f
XUgpUREBSwsSb4UB2Gcru4D2fKo9KlO1H29B+FTWNguBkCvaJzeQadvbmVC7xsYggnVA8ijFLmh6
DGajN1X4jIx0p0tcJmiPopW0Smk++2MWq3fmC/KnHpoxgBT0JvpmxFT8feeHkCJcCqXKWTh8uoSg
ffUEIqdWcLXDJJ5UNmrwyed2R+/7HMqsWLMCbsgcTWQtquOWahFLklWFp5nlRO/MjePcSzFokQaD
JVSM/QOp+9NmZOgx/jTTrCuvr2ky7PATiTP2FPhO7zd7O0TkQPkzmJIOSJf26DOOpheEyw+cBxqT
Ap0cQBunu2QpFimupbo4c+GfyZnIedULxbO7WgipTAzsjDuK8IdQsB+k3k5IEyw1WzffZ4DnNaCr
B1U8z/yaxq/gduShRPEgGG/mynWdzDn30eoVoxqLY+Qo0NqqnD218DjKLBadKsMJW9+iyDmg6Hvz
JDrUVArNWRlAjHI8NfmLrMOYKciIkpljdEe5u6Cfdant5ASUAtcFJhtOPvBvPqtZkx3y5gk4vY3r
PwXVdxSVolOADRQzAx/yCExO77RZ2I3s2gKC3FTRRAvPhmKHS3xzaEQICH3IKsmC+WN1wUfDhW06
/0kKzSRgbVNIW+u4T4H43FXyF4cQLh9mW1wjmTguvWA9ws0fN+Av5+4QHEX0t6Xfs1LdsaH6Df3v
RJZRtFlIaEAu644qFKTJIYsNJHjhHLt3tgoN9JgqbVXa96yXDn5wOfrjSDCG8YXJPz8IqhSnEt5E
gCgakxB7LqlrTBYUPqe4+kT1OJAAnKiFDKuTi+T+TMaHkVkWGbAIrQ4byxBPNC9S4nvfJAgUdHj0
wv/ZlKYWylIwzWLqwn50A0WFJ1+EhsrrPEBcpCuf2ascgRmPSKe/RWUsAlJwO+QrbpPZwn3ohILv
doK5lxdFxnF8nWK8JfPg6E/ZrDALOE0anRjTuike1wVbOMNeZZLv5AcozuQoOzBiy8/lzCMvI2eQ
T8lHMBV2YkRpv7yUTjP+YtXN7iv/dd6i8j6/6T1XN9y600OTX0EVkoDz0t/96P/xRC6x8pCVwf7c
xvDEGTTOgzvRwbEMROUnDsP4AjsunBfUjYfBXFnI/oDqsgLADq3H5m3NSb81UUyKYaxG9FGXvPKC
X02gtiDIHYsIJyslyXnKUfz3vDCz4RNucCFSq+7gJtiOfoGHzPukZB7nmoVPLp7cHoI/plVQ0V7F
65LfaezGx1MXgPre7Km7+mPgE4SBDPlcPhI74bjZhLCQrn4TTERsGvRT1npa6j9vIcqwuPjhgXam
odW0rP9rk/CP+rlSvToG/wVv5Al53gJmoDZJPoo4CbQXY3nklkflK46ZQaZUnNjc1/WVnzfwnDOT
q0P5ZhZmFo+4Cy/pWJPgAiLFyN2ClH6IKL8RvRrvtCIybGhEkqrUqx/aeT+wgBAfT1ZNXepjVotu
bH1hEoHdPIAUUf1tgsvZEd+hSFEVPTOGrmUh8gk21JVaGDE/QNj0HrwNSWGzEOzd/lzqZszIiFWh
IvjW96Mb3AmOVcQx0lGkysf0ggEQX/eQSKHYnaXhzcI9g2xMg0LkRdfoulQHRipHYz+97mtum4Zq
02+iugW6fxusje6nG2VuggyW+l/RdVDcUGM4bd2jxHUPJukuT8hStO00Y2dovpbjZQH1NdXkrisY
pSR00IeIhjBy1EwyD1HjrFh5S4brMDJXq0JBYNfSqEQrCOPph1BJNgQq8vSHM+f1o/ZP9joD4NaK
dWF6C2lXu7oPBoY0vDd2UVpw8r1ym2e6VIO1iAAsK+pxv/ipopT64C0rh8l4acYeAckDAuQ06LIh
OWeJKntlkiCdXhwNpIile03vLAST1V5u5RkUKsw8vfdQi7W1qRrLKOOfEZMHAY164S8QQVnHWSF9
kHTv12kEJhj+OGvWuRpvxABRaocGU8Kl2Yq7TfcZ3CCHKm12Rm+Rt6nDbrrUxOf25Kk0kdr/Kl+E
UkUdw0sxdQN9Me6idKhVkQOuVSfktgVZ0PzihOIwFWOFE3d2Qi+/m/BG8CRQ/g41/T35WkZt0MPU
FW4wHMVawarKxjMIhXRtyNhqYNufQocCt9KY3h6XnNsoi/JBKsK4de1Okw0OfNr4ypvZC1/YSKnk
sMFXS8YXyVzYki06dmTVDk/0qLW+rQm9ZQJD/LoxcfahrAmxXzW1OqQrsi5aqv9qpTz98DsTRAcG
ndY2A95YaOOT2Ot6OXvfU71TPzJJ3TBMzHXbNJxzVJLHu9675BJcsYieiXYYEbTdobHqSh0QCHIm
vMDbtbg7HLY9PudOSHdu2TPQpQ5nINotrcNJVpCMYlxZJYOoJayjciTrBdMN3jNHnO0vaByTBs9D
dyHcPNKuS3vhkdJuEHukh/178tx8Frx5UF5s5sh3bUaQfi/1ko3lwnAgUAcOrSPNYjv/v2LVuqFp
G/YpVaulW8p0FUeR8GHGtkG4JMk7iAZI0By3SQbTBkivAPIgpa71KvyfH/MAT3Un/s4KDFvbgYAG
vPvAATx5pyULkpDcwfZ79Vgv1tdihY8+Fn2QHg7+klKmfqjG25BO//PN9vQsmCX5+YFyGKuK/7yT
oUzFrz7DgN9lY/VujMfULRKn+aybYY0I6zth11HZISpjROVXHpLUPyH1nRysuvwl7apzKBZ+FRGh
IFC7SQOe2k7DnFrz+etMx+fiFcCd1Vzyslz9xHUsxGidUluxPbVVfLX+ElDtBDrE7Gf/hTzSYE+B
n5PUrlAnKDpBSCUGQGnpUxloQqqeFqtBTZsTRgt/2ohsloe9TIGf19qu+u88B/GlmM88c16sCZnP
a7ru0ypapPv5j5pro8qJxC93QBTSdRQcbMGDzM5jBTgnKjdwI2O/2be1JaM2CIiLKTFI0dZ8WNwb
Bq9V9w+RWTK8Qbx8NVCXgb33WY3JXmQVZ7E8J7+S6CHRIVXKBi4eFRP0dJnOy4frRXGwn3kVIuZL
Y/R/IOUqt0bsSbnU0zbMbZ8cLiyQ781aRRnVaMgfSHxDJPKJdirgkyfps/BMcKL4A3EHPR+IGoES
qgnczDBkt/aEIWkTwbMAWXjvgwhpsDOZDBbxja9L81M87iorcbpp/nis7rL7ASocOVOpThftEvw7
RVnNW++UA36v5/mvQkuVGQwClMGTfR13Ykznrb0ru1aYAXpMW3xuhUOGBdCdoVBMBaVQIw9UPNBH
q2J9PlMPj0qWuQxhCSQYHYyVS44spiVUBisg4BJzsO286WPZVFBAv/6COhgqb3M4RbRTmQrG6gax
4C2Bb1qXB64JAYZWhLeTUQgvsyVz/oaz+qhUc//zpdljjqrJawRe89tUKgbfLBMjtyjW88EImTKW
8SyORgd526CYR1e2HAyJS3CLIJ8PNO76rd+mycLP2FvvQ14gk619U6mmjeIBiCfRR8TDwarsM80b
vu1t785nHvdnZjLCGR6wR3ALPP5d0sPstZ41QzMvoNKuE844jeTU4fJGpksBJht5IQMzarleq/6g
9yKiYKYrfwenpM0uSYFZlMVqd/rQGdlkrsQ002eUzFs8l875AqVG1+QwKtusnExAX9KBfIW6S9On
F7+0qxe9xQ/38VlSIeW2ewtgAYYHZLxeJslKXTwWog7bvXL3U0Y/LDHdEInLQjPAexwAheQlRDZB
6BYsIlBe8cbEXB8Llx077YnlpggpKPvBskj597+H1ONCyKc7co2M8zCrzYbI6XLPU9BVdLlOjoJU
LlYJkAn/VIUrWoZQbwL4fOAkubo9rAN/Cfwi7jvsB31dAgO3FoHFYzz/ISUNQzZYX46EPiEcOy59
v6UDR5Oj29os1p0oOQfKXRGLj1nbkCnZZySD+ya5Lu6ZGA1lR5Uqhgjh1TQmV1tOwym2rgTbtFCN
t1O695nbjAAm9Mfl8oUitOUzrt7axz/1olzV7/ymrLi+TCbNx8LQTrVCxUw78iHnfFUizMm+CKdx
rbgOKJ4a0tkTAOpXT38IRQrIhwuViTfIra6ItJ8VkSFRdgQ3sKvojFiUItuXoBfAxLsdcDeQ+yx1
IDxqze9AGlPogE4cPAvuxzPoH3oekyozIPcBlbBUcrwCrT6+kV+FuBuVidUrmuRBePZmAyhsOQGo
uFklOVP3eX9VUdJvL98AipMKQXYBaSSq3dV5D7biSXMy5h7v+YAnp2CobdBXaQwYNNXm8fDvKeMf
b0V6Kt/O6gi6esfvoRlXneApUE3QLeg8Tb62E21C+XO5PvJNPNKGUwK4GY1D+PD71WmGF79rqbSU
jX2jkfMOwTazpsufa4Ugk5UROiy1/1BC/oo4sLJ7sBcyolGPxn03FdOXRDf8sWbTPvvUaeNgol/N
v2s4BptZ22CdaUazaRrdTbk+XIl9VYRPc6zV5zTQtgDDVp0jIJQUlULfR2untPU/SorO7fJR65Ih
fLoTm632PRAP8fwFBrMZhyKDUp1UM9eyYmBUz1e5U8JF0WQ+Z73xF3c8NwvTbRakCPlpf7giB3xZ
bLhLN3vu7kwEt4xUIK+dj1Q0zZn0w5n0yoB3A3wl5qfcS7OCY8PlDNvSCvK1j8DSGICg0udXsONq
ZHTGLunZqXP3EJmsaEqox+/svv5UMdV0JO658CiS7e+XiQRyJpuq5ebPwA3XmZmLY3Eeo7YjN64R
r14jvly6XNwchwJGTd6i2rsRk4sNbHJQxhRHzkdzZevusYN9CNomOzzFqn3YZsi1Xr2WLo+r51Lf
z6R1ZJSxscEL3iJqVy+ysfkiy797GfQmRxcSot0eWSX25yQSgZNtL9UPmyeSPArc46qYakKVUNhg
oYmDPYpsmOSnuqy1NExNZe1to9/3GF6Tcsg5toP5w5kwSnDFHJURRIAxHyjaWmSI//YPbON8bBv5
svPWvGzBxLZhySXueeYUux5YrRm8vz9Wc/F2aA39O5E/CKpyjbMVq+MR8wUrGMH3F22SvLUJWN75
gq3mXozehibfb0lAqsItNavxk0V0cEX8ID8BUbCbjMAlgLHQbFz1bmYHs4B5Ca7nstKlxdf/rA8g
E4cNqFd0EP3XAu2IMu3XrtRKhz5+j04rjym3opv0xnRgT+L25dSzTRS+gg8MNoswGlHNC0sf/YCE
GilZiLDXUFc3cVGbjjCt1EiPyOGiBoAXVSMgEUAQtkrovZnNsDwB0R02itnrodGwjQYrBWNvizYO
IkmFYFz59rhBpQbB0gpJwpFe82eufPnLeJ5TYIFVaipdD9urJE26JJQCk/XXT6GeBdDRiL66YJos
bAIxexopzkXaZTeCoP/L5GgmW+2lL+VZQ/ghF7e8KsH56xdzDbsJOncvm2xpK0u+tHh4sGSQ1USi
3Wrbdb0wPJblkk34cezOQ7glalSoMi4N9hUTlEKetexDA2oLfWe0ksuqgBJj8mRY0IP/cBZ8JJE5
gCbCEZ54Qo4WpE+gdCMe1nqyvW1JA+N0GO3xY4VLP0ncXPBwsUBA2A4iTMasYQ7liAfzeUdimzNW
RYjxC9169cUJbdl6tBTm11stg7Var3KQLRGtkROdj8nfSa9CrG7Spsk8tu/Bbs1cIutpplfuKNmB
enUa1nZb3jNeML/E2qTYHIGNfAczFOg728d9K4jVZj2TCBULBM8Y8nxLzEOf21ur8cEx72jno7xG
zsTmDOmrjOY83w//WsRURc6uLHbHUzvmBjwitJqmPv8kpEWOxTs70wDZPWwrLG35Em8hJlPnA+1d
Nhd4lsMXSN1GNkt/M6XZgzgpiUU5Dv9ZNo2w5QjoyFA2v2MbtiWncTHQLVcthkqJ2geF7Sjg86eN
HxMH5rfC2ZpOblwdiVu2TN8dr+HXZ8ILzKCB7BdLqXJMeAQ7bbfqvl5YoRE5ZtVRd3bF4qFmuXcV
DbJ723ImZM7XfrizfkX0S6ps6TtmIEaFVzWIdWtbEfeoxPthNV0HCfRl0lj83MEsP3krYI3CHwT2
Ba8vWc0KzLLNL+rYiaeQe0gZ3igDUnyBe0qEc6Aoc8mh9U8//0t5AUHwrmk+mg6Mn/ArzGKBg6mW
Ppqv8TmerRp/mW3gJx5yu/+KB62V7rQHRp/h8y+H+ERtmVWDxkFUQkCSaLjKTS6MRjXcKVNH9l7u
JsCEqnoHedCCtPrq+tWnSnnwmweFyKiQv5kxlF90wg9vaOma4xwptkhngvoo9NoJ/eRyXQ9oc9vP
9ogrxb6UqQ/F2MQqETW0pjFcWOz5bH6pkmLzfiiHXz2rRWDJgDxulYJzZZthh51P48JZMQzxJgMC
tocwJldq/noa9qDBUTCYARrCQCn1fhev5TUnEmHlcQ7zkONyHuLJtxoGmWZZ6La0mNl8GfvvPc7G
XbP5UZNyIVIHWi98nlhYtrpZNGJjXhcMhdebUw4AYj7BrkhJ5lUJgvW659IqmSQqaHycPDRVgacm
ber8oFg+ppNlr/vqbJRtZObqIe0I8t0LPWz98m66xJyCekZ1tDS5TKhYTzwBeKc+MsrvsNDRWVuP
ktjH9hXHw4vNAGKhwj/viFEXDAdXAXXtAtJ2IGMGESXXwDo4LA+gWTXWCr5w1WQJN+SAAW5AccZS
BAu3ZO8QSIKcKRDaEnUZXGAm9bwqg/14i69zUY8XRG82GVv6forXOWMHdpk664McUdXRfUehjPeM
zL+ZmCGbt4yAp8AIcAK1jwrg8WzdikohJ1lG2Tw/jUrk6AhKMguYQYjNvYON3XgtQVD8L9QBqYMq
XjmFp+yT4EBzz1q06gb/w1cn6SK7uTpNXSLyvxttTt1XNLVuq1vkwuxNFCIz/z6ghEl02DSN/vvM
BC1m09I7Y6gjn2sCcUhMfSiFh4bqBQlKVEV1C13SR7NP3ywEEA3MitgNxDRG7tRBXhz6+EsCR/cq
jkuMFw+EwHVhm/8tuiGB0xoljvgGuwoZ0FDA/k7Bs1e8ssYH7t0ZM8p+DxIz+QlLOCvJDo8CeR9Q
LYZK+7dE6bzEW22hSoRfrUDIw5k67/x6N4/gKChM3HHJvvSNcveTEMH0eLEPmw85P8sDvC2chaLT
d2cl9elW6g/c/In2sWoTJRLDKjfqTXz2OLDeSjUYDDUPu3P+WVxNO9x49fb+zMFX0rVOdD63dWwd
HYSzMsPOg5m7yGFV1MRj5f3QaVzpzEiKW0Zi+v+gC6/fT3Akh1OGIntLMqN/LU1usPZCQ2pVN4cv
FLgTyaPM5XDB8xnRM1f0uUJaNWWLkEPbXUnTmqWYvsM0oW25mbFtZGqrmqUpn+zkYfQcr0K2M50K
UTYg1KxOdVcJBcAnRjSjnH6rZ3Vn0jaqRuEsuA+8qpYX8dyIZNSydu69raH8GJcFl9VEPVIUr551
eoJFIaluBOZWFdJeC1Ztwp7hNwUgVQUW+CgX6iEZ0/tslAAjfA0UE/u0OFs38z086kcL/OTP3uBM
aLQJnvkAaUGE2b1qp+6zOSownFlO8Gi0OYcPdQROj3XCkzdiKFcOv2qsShKq/rzoVKmsWe1ZSptU
Bm+DpML6isnJClqtXxx9QBM7tAOOIxQmMpuBQR3N+UMidCIt/GA2es6JE1H8So0pMLr78D5OEZQV
SG0dQzeC1DooBRjVY243DEjRJfceqP1EP6di4yLagIfynFEjJ8rLZNRUFiIjPKZDfUe1UDNiEzp6
T6f+klFkmc2oy7G3YEVJVqSPXDUZWNvLLuuImPtoNTYeKUbyf0N6rj23DpU4zZfIdPCI88O0/eFO
n9snWuDi8lTq5ZajWSOX8TkhvJxCpP1oPyZqTOFW+VWiXzmf5flCEvOSUvHaZcLwMQ1N/wD94sCX
NWQ2HhiCmoKXAuac2bReBqaqt5t6xvrstWLNMapDjiEW2TLIDxnAVlDNO98LN8DUPnHbAhr87BHS
nLcyBvpg/1AO2iNbzdQmjHw+rSLZlzOx5HDscdPEXGxN3EximwPK2ZHFa2zPUqAcnVJfuyyri6NE
Xt7fwoYcJvYsVctk5BSojX/NOHqmxNVgPykWDN5qb+bBFY79hOCRtlbNcpXOf7X1Iyeear0kTFeu
3uVcgK8AKrO3YEfXD9mPBCPjfVccOlIXxLgn3JSyKEsglwY/ZRAc4ywAanVjXTM/oAo51XMFAYrW
p5yjhJuWbgruVv12e6TtzkKBb0XIz8hlKhVbRwMnVpRAHqDJ7P3z8i6RizhzHLfNhUiJSolDs1ba
jxYOiswQrGtkyU2gVGYyom971L0Um+tZBcB58QB0woqqeX0Fx1nheQiqwNHvnqY6hU/eVVb4BGfe
mlzA8q+5fF4yASS63k0vepdDcLPhE14fQeqIwByx9SFO70/OhQLSpTpARtSrq11w+7OpsNuAcwrw
1ICCLeycqbsaZ/eOTxWEt4xPClrsJPZgtmcGupmW/HcCyYQ2KGPn/NA/B3sV07lv6UdyuaFaaIjT
sb/eKCXGLhJ05WeEM18ErN1m9RKpYmb6ORQWR9zPAHo7cnI5cS5+vRGbOFiRMypId5mhpTdoN0Jr
SLn932lhlcHZZJ2FRtvLoVit8Dusl4Gf8HdbQHQbyoDUZqPAlXl4FKbdndw32ZPCVgcENzJ8s8MC
lzauPiU+TPw8F1Rhq486FitFXwortAVkqHzkEC5dr8piYaNTVR1gtxodGZORtqkSPOyPnLAn2bUR
XfSvYNJcdYFfkAXRGdw2DyNaoWOj9Hbl68pA1fWS+LAsAjFBrXLKoxct7Y6vVfZxLBcXJdyOLM3a
tjJrngUVIARKPpkiL2Y5EioqEwoQ9rBC2wEsJnWcjT/Iul1QHbxM+CfIGQ2objqN6DU+PxV0zrwV
UVtzK42LiRs2rWYV/3WGx9tym9CeW+Cpr7yMwgpKK9sJz/9O9JELcxjOb/9Wy7pyavz135lTyfvB
XzLT59/FqVg7ot53Msnsio2ry+9TTDIbDdOh2KPDnNhqlMRDVvbigcwFhu6H58qP76y8fNzZbupp
x/xkWA2OWPEoTTZwGsVy71/nUe3lcdadiVKDmSCctyyB3wtJt5E1bc+WGcB4U1q8VjFGIu7YNuKG
1GQG74gsMofrMeLrpOpvge3YXqRWUgeaUt1aZ8Krv4bM+7eGS+qrpqsyqOvA3hAQHaTXbujy2Bq1
1/JJfOYHRLe/u8tKGI6YL8DnsljHfAqiPdCQisvMDSvbij9VvbdqWiGgHArESzT+Ef5CcbBkG/g9
LIxiJUaJMJiOrf0/pscBRtF5ohFuT7XqVca5Q00x99A70lAp3pBCmmBB9tsIIaDyyps8nzbBlN9S
ifzs0wkWAdkMXf33eRqiVYL6t+jS56PX6hnZ22uCUb4SjTB/UfzTmUdago+6xU3k6tT/kg7j+eJb
ofdj+WK9frF5Iw5cq7jOkV5CMHeE+UxqiSR8aQfeblTQ6uDpTPfzHl+48ocIbmCS795sNzuFcx33
JtykT8vzQDLnWT2T8qmygaqaFP3jbL3TaRinSimZWJPsLt5O0TnWOLrNBwga+DWkH2d+eFv+9dfz
yXsq+Pamlo8zCZteqhcE1IIUCe+RGSIsEl2TGRXwa66L+idMcFY8aTokXiIgRrhsaT0Nk8lGYNr/
5ZduZl3hDsXCvX4RMtArb84KNit3dOkgmLFmQXfHkeiq1sSf2fBIU1U6hgb1+G0kWhpu6i7BTsNX
LcuTPXL2zmaqSIN4m6ErgqTI0n7/iTfGttrBz2tMLJreg4BJ2rvKsQOtnyVcqPjR7fTsdQgGZQL+
m9HWTssLmrlKW9zb43o/HQjaWGfGQZwZbhM9yvfDuD2HXzhB0mDCsgDES4unc8XIZQcmwnKRmwr/
nC24gg+uJn3RrBP5fPVPouGN7ulrAH+c6Ju+EArDN+JmxoqMnRXmcAbdzNjlsfdgtvQVpJ42ONql
1v/x3bf12WPhfuDYtNgTz8Gt45sXRQUNcvW/kmvYJkbekhdPevPByxmc3sYBjUN9D0qQvSIJVQNG
zEAPVax+v9y7tAYJEnf06oB7ucDXLX1mO58b+AgAzj0JO3qRdA5bxSkqspYVGZFDvhblO7KaGUpO
HdnkWhmLdZ/173L5G6pnIS0zzPPFRHfDIhRwttUmVY85+OmCiyLLgWskylkRtfLgxbI8hvkodjBi
cpDgvWa2W/PxfUVhX0KyRDt5JhZ7hrjpkTLMNM8O9rjyZSWuKw/XqcjvyoVcKaphqGOVYfKUyTWM
yOZfcV2SDNB91tir+hBwxFwqrKSmHXBj0TeOFoNVuwGb0a2JdHDj4JSePOs9fYjKBdhfVFoKsqIT
GzCd0H0IUv/GFC182Shu1aWiYsDR8YJA0yhyqo6ei7t4wUsij3cZFNi7GyHjy4tSuqCkRhknqYAr
CtExPiV3WZ3QziKtu2A4CAfYTGkZHfQ/yJczypPXHNEcPgA18Gfpi5vNrHVLaBryLosuWPLohiUK
COAMsHOGs9hW4ASTDajcH1D7pa2GHANPSZkXDh54kWoZ85wYk2laeBl8D5T7AA3I60uxXtNT/U0l
bJna/AOO7ibP5LTcY2daRibnMRdknvv0NDMC/gc843ZAx1KZZWjwDYsD1gA7Cp1xss8kQ86ZRc3x
8gHLsWhDHH/WrLU0IOAkwdRAdoxn/GpllXK9Ry/w7b9qxcpPFM9ZvcMefz8usZiD7/1mX2cD9+QN
TYnhEJmqoqrXGcxDynhvx3cWZ1O565IOWBzDIrFe0Lgx04I7wlQf6xRfkEfJB/pWyIm9BJXvANUD
tHSqKNikT5sHjSp6IVhCNHHeK/2pbbCYFsziwd0PMfJLpg9uH6wcpZH1yEQYcT0+xsz6KK5jlp2d
MgUk/Pz2Yn/N9UB+OQ0mOn7U0UbTdLIHmHpPB9ljyUUemrQwk8b77i+9vU/PLGzh5ErHEg6lfMEo
lmCpwJ+LOTeddTdiHN8zvsqxzaPMOQwpjmz/tBLRCcRsKgvu7GFoF+WP8U8+5nWKjxPXioxL1JyJ
pFKLeXmv2PE3ruJsuw75WIqUy22OiMRtNZYo9vnMpjClEvlPKPVIfDQrpfMz03kxWD1bT+XZfFP4
97xzRY3PuPqO/vMlWO/bVBno331KW83OFYKsvWDQz0ZW3XC+9qne5chr2qhPRDH5rnvHKB7be+Ar
RbBCWlgiI7x2bFAmHrXNBEJ92GZDMRvCAg+33VMZvwt4i7q7KwzXdBlq2hZsZhZMoLqk1rt3Bzf0
9MeKkd+02262okqV9Fs5Zx7UCiKA+VA6npbm8xymD5os2jbiDyqwONTAUe1CvVYRStjQtFaCkaFw
tIkof4x6q4JGh3buUjMDq5Z6xqDegUkL5c4MSdNlc81WNU+5P7rEf7IDFY/KMqaFw7hRUQ6+VmWU
puTcdhCYZdwNu8tVdBWT5pWJ1ecsCIMEE0napNzi/tyWTGCSvbQWx3LDfpVj6jRi/4jg4PlSWskn
WiSqrLCAeFtcmXPjIsQoNpTs62j4RWVTXFGrsZBL5FgwUZaHSERCYhQJbEiKY0MOIIX9TSbC1+b0
RNjc6SirgOb7/EROwPE9wi2EVJGuR1Iv+YsMVjClRdeeiJZwyv4OQ53IvFyO2HO37cvS7/AimFqo
NBTjW/uuW1Tnq0iD+zIdb7ogF7qAm/RIA9B9djLX+p+FL7Ybna9MBRgAtCMUpTUSlaRFHavJkCAw
Pu1nqkT5oWcquZplAKUL9rqyRUtDEqxE2RpWgsLJKR7fZUezvBPIWCCvrZggaIpoTKA+zZS11k4l
QqTDnR9ZZUClx89Qxli1E3z6BwOM3RNbG7Wv4v73mC+5yqC16LlQxA6zCJDzWcEKaob8HgwMgO/b
5RtcAnmrKOhR8Yj4hcQI8xT0SdeSmOdiQMXxRA7h2UbTIHOfe1J8JS/ODGqbGWJ3RWp1Cje7Xu2f
iXdR6AOZrikyeA1LcRJrkKWMtId2Fd1Qc/EiO5xeQ4Yy2JoK8nbJ0u6rrMMzdrnU1PCDbMFmlar5
eR3hDqfO6Ge9ehsJZVivmXrsA/1sihCgnY1FIMrmyTYnZespDO0hkXICqNHIaKl/GJk0AcK6h5vU
yxb/m2igGwixdi6k6WikcIDl+zesbTCkEzBFla7ticvX1DF66bag3czYhE/HDbsJqRa/gjMd7dMw
q4jhO0tTDHSAeJYwWMSBAyOoDBwBirgpNW2TNjsaK3dkuq3pXs/wNtvqPzOTOzrYogW9hjuwzPy9
gKFMuOYWg9gAx3aFTzStIYBIMGyyOaRuZ27pRw4GaYcQztQLsCduJ/HswV/zhGQdAQ8uTtJzLwK4
QD0nMZNrIGRuiQRKOvAlobL/0jtzJvikRlrl3jl4PoCYxDCSXWrWhYtNKVeqzT4InFA7w1e23I9t
F0Kbp7aFTxubVl6x/TE3H68u9bT9v8SrS5YIo/6QCoZe1OWRiswWVkHEEO1PhMaCvokuIWlR90KE
b34DHwBsphuASuT38PEIT37sFlbgFXO4LiK6gFPQgT4mzYnpvdwbQelud3q/YG3BZ5KM4hNrRETg
q8P4A7VE2pmcGsx3YFXw0FoXlPOf/8etYMJnbn+sTznOAoltX2Y0h76CYT8eCaAmfzxXa8rCthGg
QdjQCfb6U0+YdBsztUXAO02BYQA6bli2UHSML0ngXupbiLQpkQsjmBWqiBQTowabMvcnVTpybzi9
AQaLO/rIUzangH6tZ6Bnx+n4I8HKg3wyq3C0QqPVnLpT79UXrsqfRHKf8Pj51/b81pjSum5vRues
JUwLLfmxdGd1+Mn8yFMhdegoQDXM+5pJT1PuWCFWzh/OlFnr6rMG3F4nYT5s7Oh6SOr3iHmob8t4
OUSHQSNTS2AGUIflXOODh1qe1tTY6xqLPmQF+wWuorsG6ALJoTTkbnv+rDFjcfkHBb8mRY0zhKFz
b/cXNezzL1Y7TTLAibH7NlxpZMR3Ir2AwI77HSFGKUGYKHTxdFxv+nzGCrERi6GM4OJhGkMlP5G9
+/ALedB39/0z4IdtMNdZWaAcpl6JY/OWpvvb1SxjnKNafhFbtAdE+jfto1wQxX4w2PH/86ODYdfj
GD98x/hTgzE/gM4w9WulPyMhI/ekslxAKYN46MGaxI/YpqYHEPwNKG1rq4h78aSW8kgo7zf5JuKX
kGSAgobLnHhdkSY8NsRGavxNphG9+MBL6kCMnOdDYFqjN4zlO9e2rpOnd4Ldvp5MI56Yq7J/iZ/q
16SkqZipRsxlvrxG4zJFPVr++aEtdHdLmGlEeuxsTVhMYORlomhkYQ2PytIM1SGxZi4zHNu9rHbD
1eFah0L97WckEQaZB8BAx5LWaEgJPkFxq1Zeck8CLX+vcEn2DsBNFRInUelrZ5VCkgeiCPqCN/iv
emeSlmIhrNQhwdFT6Inn5FOqJzYmFQLfjUXGT2pv4a10Y/R8f5CLPKzVdqd+oRFH7S3dmTmDyXc+
7bLeb3p0ao8kO4VHZEkR4qJoUiUS0gGtPfO9d2eVDYr306EC3nfyzSwtiIYi3YZsCHd5SHB5YI/S
MNTanopRdtEBbjIAuprABfM4I+mHaLeuv3STLvS4kYIcEC5PIicSiegeHOY+oV5fhmyWtmgXOzON
z6yBYMfFjB2OP0nPKAETFQ3eR39DySuvffDA4A9JmFvpxNkl3Nz0mXWBvQZsGl1nHB8hi+5deZf8
PH47cOp7ScwZneF25b7TpJrquNaprBfZHo5VkLvwIq2ikV9dGDcyzM4sRwifeAw9c0DIFpDq15pB
Fkk5N9+yOFuCkU0GxTrZUjnPfgD6D7pggjyq3nQ1TG00cdjsDUZ5Wb4Pdm2xRC9Hkc3mhATvVuHo
xYucKDyLnMAXvl2QN4cOyNO76/SNKeK1UtO6rzomzPYSs/SOFbvz/sCQgzde3iPFlWbEfasc/Wct
6QQpeX20IOmJ5s0Vyqjvhl5YUk/sG+JJm74V4dkFg/Q3bUNvvnOrA0v5lYVjOmNFisOfkhdr1xyn
JrjwJV0PNXAw63PE0v9r5n68vTJ7pouma64haFYNI5EqC8cSylsFyPqFNa7S9e3hx6IDDfKrE/zI
ObvUnUhjtiqtJWI4hvgIC8Q1r0uQLPq1fHKzg5PpYJTN2r2CizPoJPwhX7ZNK5TO0v5MiL1EU34Q
IWmJT3qkLyBWDImRwhmlv77cqzORcP2VDid524nZxMDrbV8m5yQc6Seb5MKhBRYfpwSlxdztjxRJ
XDfQpZ3CFlkoMR8sDBtABdcoIcr0YKXNEZJ1QexRqZ+CimmGQyVe1DUD0pa66f16sW+lsyLQ2B+/
VcUKhVeLj9M6Fp6Kg+6b5cFhnJTqpR9iQfGKyLLoBSK58iGoE89oEgYM6qKbNv5wRm6byP5bFNEz
K2BK98YdQThRiAP+PactB2+2w7mqIBvN61v5NTEExXQ1AlO9RzGyMJOnioXQjLjXUnamgKfbjlMS
KrHN6krPt0X5G42j3Vte5TrmHBJwWCLIMr1odKVoVf+o1SbvQpCr0w1Jg7n1pXALXcVfU1SBvWyz
Jp2GyfP2ydED96E84ws3I1AyI8Rq2s7mTNPqLOf9e9tdukSYv0yNcUdIA2Xtw6aKFMgFg+Hhf8g/
ivxqdEFieXlhTZTTSEQNwBe31xFYlOLmBL923I4oF0A99mb4s3hdgGJC955cHmmjRVljLnAoU+/j
y/gGMODPQ2oacJ0GG1juzOhZjs964ueT1YFLyKDonGJcYWU52jchQk8MYIu5NfDAwZOFMLtti2oQ
/X+3KGiimqY8MBY6/7CwNA5j9sP+to1fJVeRkBliZc+xN5pChxmlwtt23Gg/PMoMFKj5AdjHshdf
/k7w5WPZ/qSMhyotUpBx1ATw9VcoVJRNSsepqKcneCnvi99y6PDtu1HNZhxWmt9EwsyzyxksOeVG
/MCfZyd7IaXQyQYN1unt2q/ZkPk4JM1oJsQiMKk/DId7WM1QY+H3KCbsykC9mFHoPhw0S+3Cx8DP
ggKYYn3vemdKJSSSO3b6rp1zrZvNU1wscAcwyEDN3HdcqFNrG1DSNqnj0Nlw5wjqqW/38QYBcRzu
CRxmtLj5sgf8oARiIyxM9NoMAkVd+bfVonexBu1fAIFCbJFG3WrvueLA/SXCyJtoEQcF1LDW+VjE
SFqnsIC/0oSdgZxWzMqcR/Eju7Ndo95W3tRhJpRqqUboWRfN3lvY+SxbTfW4qrF1glrB/wD0RiWI
iXeNwnWkKJsG7eeeTzMUsBC25pZ3Xd7s+sN+BssUY9+d6RfjQlCykSP+CNEDS1xlE397QsjQrBtT
pNcZgl3K1kKXdKG6Nd7Ec2Zs9m+77x5Q5U5Sicr8XN5CrVpkyr6Rc5iEzVNih925dB27giBf/KQ0
v/PVHRigl5wzGOTr6yC1hbkFYHyAFKrbfH9J28YHI/hN/QCFPSquEH4NwUrEx+HcKYxu4j/ZDAA3
RkGEsYT4tDS1el9LUlQFyEBVZcFPLupEWPiul69cdNFgQxfhaK51lymDYkDn65AKIG44wIdRj3P+
yQsRNNUEJUIXzGpcP1GGyG75q1CoH5GWMuJIYY9wCWKvKh233SaD36qt0BWOMI4saNwxfadCGnZj
tZ6EoNqbo2QjzdxQrskC7zBmKOj/mrBN0L0Bce7l9eTlg3mQ8H/bSELNEc839atnMe24imu5Cl31
0Q0qSntad04NhRD2KN8juESZN7/IL2Bbx6a3ubnWaN8SLpb+cvOLJbeAnHWPftrFFb6saGHIZuYA
TV/2m09FIHq6r+0XVh/8Kk8sqZ/5iH8AnLqIfK+nXHJO9qqOOPBV2Lf4k9oK0nP30aJ5DJvvCLWt
4sEXTKa9921Hl73/OGBmHbEiVXwEJxIhwDyvgcVBkMrFbz7hbAvlotKl9FPqeoI2i5Q39J67uA4u
FfU5yWAbSdQLU6G34XvSoRaThYIJJ9UPnM8gUMlQvJ/n/Ak1GKkIMMqA91OWJcNXkapvQFA/7/pd
9JE5GkX465h5ljqAPZ7cWVZtwdw6CDagZo+iYywpoMwnGX5YCisPHrxns/zhQ0KdzjImYqv1J5Vy
8FX4LqhGHuPCpQeZueH3Dyg2r2dAETnYRDUlQFrEYJ5GQtnZHnOV1igtXKhdjcbPlkpZzhQFmehu
PA3E1DDxtybm7mVVYGR585cDPbEsALuUOoqKoAiZntxjdJOZrhPn4MWnssEB2+n0XHRRz0M0Nr97
UkVOlCNwvWUP8+dHgsufWyqwvkxX2lX2b6WGOuAh2eE/cxhuZN7R4/7m0eHxMrIpH5lwLUI8t1QW
ov2xC20p4xZQa/EOEOvpTshI088kHJF/uUrIgeZ1BQSKrym/26vepiiUQHbduWFzkj0CKCR+7N0X
Wi3c/YMkTdMJiZndnozU1UMQ6K34wfR47LIOeojbvC+NCNgim62dZxpKO4AZyVh7NdKJhGltQytQ
8MOe07M3iT6w8oE+8195CoMPEdE9OALENUxUp+PMxu6WNpvMbln3p/NiD09zK1JGd16pGTwY0TJv
3s1+y4pKOOjghLWs7HTVed0oz1DSy8ioZeBcpEuLcsfVo5S6LL6XsqswEoFNiiB0+8a7XBse4WsN
kitRcP8Q5kCKmGqC0ZBUt2hvV+l8UVxNHXrDUTe5025dY/jK3AODKLGi1rb9wffPu8/u+GKZkvjc
mk7rG61PHaX7ZoHIXLvj8n6FKO1KOSWJTIfvWFO9IMqEO037wkRYDhupZKEbhVFKZDVka/+eHf8c
0RjlOXttsneSN0t71EW87vY/mEZ6VBIvTho1wecgveLTdcW+n8UsFYqZ8UMToSdIQAYeyl9b6vKz
Oy/CRxcOVMlZJObOq5u85QHzUgr0MfvnYMGRb23VXsgcm4nMjHhPmgd9COd8FwDFUcW9nCHPmOWd
fRTNLbW4BhO0dk6tMJypBIltNie9UmJUlhZ2gA86l3xJMTpW6qfkvuJZC7tVAHFWIOd3DHmQ4K/U
MFY+Na+vyHbGfZVzEqNIqL0LAYKwTbUa89baCfxfqZBIVsoT9HJOULM99odpTkOOujoLznTmHpv9
G/N1zR/EmVHyOQcLq7LfZfjHU7zrorljJNb/XOp+c0plhPDh/LGY0q42ZxNRtKs5ibqqJP047EhP
MncQui/4Bca4sNPZppRLi2EuKWGGD5aNzRe4aFxcauYmUGQbiTIs3JjWMgJQfxM3+7tACShxRTrT
OBneuksz7KVnGJkYMFVjewPHWluuNDNgj5GdpGPDXVKa9HIxk+w3yoMZLdfAN9YH4fDrygaINOj7
t1u+Y8Sz3vnFvW5yquZW+Nw6aiZjYjq4x/5vLumrY+wkB9MmglcadN282wYOtySZmJvuRkBzFHdd
tLkSZvhCCQp0NwwReaB4uaTdYlsDtwIEfp4JFUcGY7csXbQqzfjPtlAekr+SYfZpPpWmoN2zm9fM
XQbVSSOsS5Y/SE5F82Pz1W6d5is+Vg/pISkjsO+nvNVz2KC7UP7B+cOqp2CeVt4VAtxqOnYReY7Q
75xrPJW3smgZKvkf+B21sCLIuxwMqc0VzjfySuZAauMjdT4exkmNTOmt0JhEOVPvLD9hABmF0Wy3
88hcg4VnIUoAeCC1XDd5k1G67pdQ7H1h2fIV5sYLrMdR2/NPkm0cRfLJQrtxihfFWvmgzbQU1Nkt
xHON3o86Bc9DpVUvN/gx3LRfQMTqwj0DL5bf7hVw3fO9FJg390PCE+2UN1gAqlCzXa74RZMWbY/e
LNbE/AEkKK1XRUYsOWZCovM1Y+1mRloLBKvEttC96ss8vpOkUTi9zahwTfNosMAaspifmaXCiPtn
+g3Yooy570QzlK3kwOyPRbWowbyQxuUK2yfIfGa5wS21hsScCtXkrGuIzA5a0qkpAdw5mwQOhH3b
27gjnva6lAtT1FqsdsJ7d4cRmvcAIbcjsb93K3YUSdOjN49EU5H9Fisz3N0Z43M6U0x5+HsZPVgD
ECniVzlT138oCita0aah9hrP7NpqJW6BL/3q+Z8AWwdBmml2LNX0K2xj9E40emxCt4Hmn3DElKhI
A/9EWWlLnNB8esyGvNYNMxkyLTn/HvAKbB7KyEJylQPZOARGK8ktZUE0TWkDGEqa0PSxFNejNMXN
gB/8/QIwiJJOZFL3Oe/5Jxc/e3V9m7eYEdk6Zy4wMBFN/H72UgZOtzTRtpbpkkQvFAWbtRKw74bR
k3J5BCoyxv2k3N75RPrDPDszgEJ1UXewO9LScXLws/RlVOTlX5bzg3r8TRGE3RgzQxypPdgXcyHd
9jG1VdGWlqMIZBgHAgfIeA6Bst3CBieh3MKyUTuklT9YVmfbkRFn3vZyIdUYJCCdd9LXts+ofdhS
BvWxFOaQ5Qs7yHJueTqLbTbMWZ3QQPT7+89wNFrKa8O1W1mXgnwApQ/Hxb0fllVzH2EFSKnXFrpV
J3cz29AjQaNuRziNHfb0bn6ZpmLWS9dFspEy9nxAIQxOwCGbM4BPeeWWaKKEdY1qGki4iZRy7FNX
Hqm0BRjdt6v/532111ABAiL5/r8mh3CR6sD4fexGaoI9ZK7n0iqjUCrNwlyfvW0hjS7bVlz14jKx
8lZB852oeaevnfehRCGP6d9/olUAwJjqBX2lUVVEVb8arS6645vI43+xmhjsg+yUl3f6tTtLGXhi
PGms3MRJjq9GEXcASV4alnb6t5+SFYIFaKyeE028z8CbJ+xLwmB3rien45lBAvWU9k71o6veo6p1
mT5QaVqIUvaHLEUmH8EBzVUJuOr0Wl1szCR/NZMoHLUiEnKYSZ99YrMedmqamTaULgq2Q9fKY0Sn
GtT4b7fsuzop0m1kpyQuN6ofbHQzRMmrvLhGa2KDIjx5+DOjXmmKQaADyFwxfmIg1zgmtFHcT9eZ
xgaKfo04OP6uKFVIV5ejjAp9ZOSVdO+xMOKpXaFCmRlM0BQS6Y9S8IHUULCmxyLWuEFA9LDqAKOx
u1sh36eMbP2mNPK7U4ZNHzXZ8M2zwp0X7mKAXsPFlzUJu/Jnsy6cmamWz8rnaS8HNfOovvDetTqT
MDmcjiG1lQDy1MUlRlYgkf+wDIthJtCYh8vXbC0xsQgliHVTXZ64QByJiYJD7tJmsmIrbH30L3vs
nzk46pF8c9SUjOKaqoeF5oY3yUZpMpO6CqfocyytY9PHqS/EpgQOk6vYjh4uG5gFu/v7bHRIBej5
tHzvCzQnHWIagMlLU0CCXyyAEagzwZiVy07NCh8mppR5dD43/LyozngLp9JwwFQF+MJqm4AI1DyN
doKQ1QLzaC+xDB4jCuUiX/v82ClrGRetgl+zK73Ojc/oXB9cuhNgd3vJsE0sypFO44oTCso6lQav
3zTPe/kUunLeuoqubCpotiVhN7tj5AdS7i7t4Rlb++Vq7t3+lW2iOYzp/b2aF9G+/Ki3awCs8krX
KyB7gZFUKX76/l2My8/iJhKlrLFAaRxlHL9cF7gx8Ji/vAvW7rXDiJ7VVQPlwpkTcCUWb4eMztaX
ho9agj2GVxGu629rV80Oo23C+qlh+mr5PqJmVXw5ibE5V1TLhBUASEa3lRPl1zSVbpK9m8rNdA4e
GWwyBaIzsKJC1rlrxIJhC6Gh6BqluFWgbp77RfmoaMcGs6ReWOLA6ztyN5V5bbyAILfLfmksWCz9
NpUOdPn7n/7vapiQ7pRox57cV656TH31HilQUZaBApiFqznyqA5IHGSNTcMBHnBBzYgvwdJQE/wS
DujKncuke+UbUvaA/n32dhfxrVMMspAgltGbe1iW31JKGe1JmpKcLZvaegIC8acIEf+gSFpazO0x
RRVIUfXTKnE5AaS9SR9nRmleMaco6HoUcciI/wzU8G7/Wot3TWVnkJvGEWyuHkhEH5+4M8UYq+8Z
4Qcp59MkeIpcG/HE0IR6rRHkWy5PAnXq4Fy6hZdd9dY9o5Hh+Qd7HVMR6hkmgEAcMyQm+1cyovaO
qn8WuOG+TV7UjB+XaeA6ZKtFi98DLFsATxYfHw1/YikBg0ve9xrA0cWTFVfgoYM/uTsbEqd2OWfX
fznSqxhJEj+bvAkDZxBT/OnHmjSJOhgeA1F+jHl+PANWMa8vyv9FoCQvlfJhjGNt0PK4BWMgUuBq
K3LlKEhhP4MCaq52LOv1DIycTB2o1YYyWsRZKMaGG2SwyADuBc/jLEtEfOZftKl+cKdN0Bo7ptyH
Osi1qGEZDiqpYioR9zZP4TehpgN5gXN63Pa4WUWlcVe/SBH7sTVrLYg/UYScRlZSY90L8jhwdA+M
395L7cx8o3YuXWJNkLX4JtQrbyDO6qqBP3WoKcCHod6C2j6PQ8LWXghWXNIf8jkGakW1NqxtfR0X
HjNz1fHmZQqj+XFpzM6RB7f12UcCl8RRzqYPBcmdpXEzWHtuS5bJ3gb0t86VAWx/cRm7vYxunqXT
y7j939VVXvcjPlS1powQQQcb3Bd+lGGrudF18pIWd3bsamozZJEwJ14hAKhTKI2eLzeIOlWgu3SY
VB0BA+RSBqW+p5sxjv+AKbJFh8jIY6kfC82NMOA7GMmCrFKQMrsF6w7n0iyuqfdjG1egwzmKdkm+
eE0lf3vBztwEMFyPhxuFnduh/AQ0xq0HVD6jsagDAyxIQfot6c3pKtm7LC+RIFtzLlEQiek2wJ9M
UeCnyBGKV9cDKIwYVwYcFCQPCQBN1yDwb87lc82pBwJrkiptIj9UruktQbpvoPka5UOCAxEUBVtm
I1c5g7IrSXPAHhCXmaSfkMiQSrzGyr7XXkigZCxn8fFaWzL1kU8lPpr8ulRiHlA/O8NBk9vEBX+7
lHnPR1FnYdYXwahvo/1VQvnVXMkb/QbdCo5F/r0deAZlCRz5jibdhbCHlIIo342kPw+McGr7KFDU
t/oPnTSQh+hPZ6AAVKjvqRNiasMTwzl+GBvpXCe6ZZ1u0LrBjn0dwvtBQLMQW7RjKl4D2rwrqnZP
LBGBgt8YOUSKaWhsU85lH+x7OZy3goiT8EeNagcpw8BDfr41voCf17wHc/PjSrd2lmTQPRadLmGN
RXGIIWUQeiAvBFoKwt1RkICMz2CQc5x9IDWt99c3Vi+HwC/9icUGhEi6IdjTqlFPYUo7ovw/lpGu
sN6vMtHPcpDMj4DxJDAWHzNfv+cZdk5K+athIROSjLlvM0BRbQjKRh1VwdBg3VdUyk/qhyw4JNH7
wCqk9BE8QEpB3QCMiP3HWVSdUtYu23j/DGsjSowgZ/6ZeCH9ipzAhP6WbgzKbJ+7yoArr1fsCyzE
H4sglFXwMvEKGddpVNetl2WcT6aRwiV+zgTEH9oX9dTqh+Ove5FzUxJIWcqcQPxJb2++bzpP0LpN
8/JJ+vYofVCVVONxpsX9G07QNaYSp5ZOwvJq+geyU43254Ut/pUJHtuF2WWDGw+I0nKUg67UVE+f
gW3JC7VqZfTtUOum+8yF3uT5fpkKnEBi0+b0RXZWUW1U2IOFWDy6a932bxKh6+wukdcYEW0Ek1xX
/UtRP2rz0zj3MkVqyaCiRmwHbq0fCGGS02uub8qCZmHEGFcMwOtaWv7sm13vs2fF+vZ7xptPII12
lGCKdw1JHBqMjoqbPj2DXokXebBQ/buX74ix/YVT1Wgq2jw8j/4DAzL5zoVEBo97wAtY5rlCvRB9
X2L3ZdSaAd6oCWi/RW6YkwiebGb7+78IEi/WcyS4xAGMwi7v+HqkjmN3pI3RhB4asWXUq4CTfE50
CDFQ81CAG5wK56XsF7TiauZ3RQdrz5VqaJi6pyRSmQOie2ZU8KTD0fsoycQnuWEHCAt7faI/jAi1
1Swl+ErJ9queI0pTam35rhPts8JEO/QmvGduzwKc9gQlViKU+fGEW/WHJYLGCHBuK20mo2eZai/Z
5tiJCwQm42sDcjubwkjK+G0tELbI5HjRSfHyiGZoXWl/VYgtzM5q8pBQiaje2KkiGNSHIcgo8qSl
Vi3eiWWstJbg/ad1UmJY4WXDMNFGCA9VGoNzeQNJdiHeEAqscaTD88ACkS3Ame87zYoyN+G2jqOp
FqY4tym92PbMhOkzy2QRRLXPj5S0kgzz7dv5+h5kuw+LqsxMNKFf52Ro/b2gmAL18K4F+HtazNXT
jGchbNP5WRwTm1jFo0biMiYFbNvaG9Oeydqq0esnzr83816N5xqbt7iNgw1cBliZCvF0pPnPIHki
TNs8xatFnjFPq42rjpYInecE6Lgpw1ulfGbsyF28cOgblO54IB9AbOxwwldJ06vbZno8pI275fA0
ChJd/8/augxl4ozmWl4KNa/M/KvBukl/dqtdBhCVfpBXsE6PEaUIZEE8ov6XwIDgRVV6yIsA1xZn
RUxIl+vcxrmvOpvI2CKZ6emV9m//wF6Cp7FVkGZNu6EAL/bMtJ0TT3BuSHfWRrgOu9l8r8+ysWrs
5UJqz5jOaN1E+49O70K+kOSz21BYgj45rzT6dQimSrVGZ2IgFcWNyAyzNs6W5QCmtyV6jbEBK+jV
0iH3KsivyLS4zs0ZaPpb2dpitzmAMD0TrTFwQdv9DFT9D9fFJ4fvdWMpTUmsscqiOCxTpCz7OhQZ
78e4XdAkauV/3wwmYZy0xhqqyZeVxra70UCtKMHyz3CvJbTG9rZFgmoaEOYSJMywmOgHhyQCmJ1O
AWaNmVRcFiv4khJzHmAe53y2azLqKeWYPBxygyHa0teUZhpIJZt1E8Ovz3VyIYNhzlJKt1a9w+OM
fQZ+VwWlynS9NNs4hP0sDaTuhWrCp1JaU+aevAxeoFWwH4Yz24dL24dHUhcsYGw7ChauPCrfF9x3
tLAegUsM5VIqD/pDetBFW+GSEedu6U5uVJi5etjsgX1jDHxxoRnJ/h6lfvCk/58QZSUb1Foy7dvl
ll8S5L5Zed3fIwYVvPt9HVboh17iDcxeR+EFYs774QwxJ60S9RAoeA0z5Z9kdE91Z/OE8AnP/Xf6
ahLuuI3jk+5RBzmGfFYHztyy2EyFFiI6oDNpt/2tLCD6W1o7QXmb6KxcbLWmvUTLIjJVir2ZEJxM
CJCbD2SJ6K3dP5wb8RIVCSoaDjiPWIxz/KbBT1mlzH8FUOKQVhSkuMpT0katQCGZVONvrOKQtd/i
fGhIiC2MBKsOnfMB7YCqVYEeHOpp2Yr32wUZ/0xik8P71qCfTsciK2kTvPTJjUZAnp5Rk88JebAp
LR3RS6tb98C4M8t8w7n0iWUuCm4ztlzTS8qH9FAAEV3Vmxq1ikWVIPTn9XnHHTIfrr1fzqAnvhrC
DSpavDKtosOFWVvh6Snix1mLPtVFDB9zA/HLK+Aeg2YQ1/LrJpi4YwadZ9aFxz0tzMxhwUjmPkOf
37WSAVqnrmrw02qWyB1mOnMzrIScztrDlRyOBLhxhWhVVODRD2oc6JFauS49mkNcB/2khDMWOClE
vLABiZDoid6Migs1XM3oSGjAoIyBcyTBD1ie+reVx7NXMjRnRIaYd3C7alCEYggkNkUGcZ+G9p03
XbPbl/LHiodERVBlIq3nSwox+vqLLgzt+WC1Mjw0rdsklCfkmBcJtO+UPOrKOZqDvlKOfFjpsdAC
bFRH0JuHbJ0sHi7ZzJIAKDr+UsGDNigk2GgI2zpSxL+quUVopCXydZv69jXodx/ARB56kiUbbg1g
DYPHgKBrpPKtvMOMOsyKQ6XfcbhCnMyoHxRiV61+/AT7b6P56jYx6O5B0jzWcPbdrkzmjZaoEqP7
skuf44bmP3X+ODOMktSs8luHDHqwMHI52fNliG0aVR0kmaCDtYwU69nezqT/v4xm1zauGbFGYNyM
5QitX56S5uj1cC9FTrrpxic3DgwIJ0Unb5PN20HXnW/mVwd4axINRkMK2E2DU9z7V9odL+UhClPe
0PNulc8qcSpYQ+BNrwqXiAfDU3ePvWLyIS9IA65WImWyQ7aSXAkFf1ztodhUOW1AC9uGivc2XZNE
R8gKKwVvFLES0j0rHoCUYCE2QUUIsmlPpzaF96KTYctMPYL7Hnpx7u6nTsYR7do82dry9mlyhWeq
p5OnMlQpZY93ei5uMu1EFvXFXtkf5ZKAL3hzU7zzLCviQxFKgyX99HJwROsHQLwKsciEoYP6uObJ
zldiqqNoJAdfJwpT8zaOErDahrx552p6I0xZf1swP73mXHwMB8CXAVPOkWJvE+tD/H2355WXKijd
YQhkFqd/OvBH7AUJTTjmiwEyRtP/SS8TXUiegm4qPoM7Z+zvzHrtLQ5ZhiLQSL5qCNFGoG/8hIKn
kIzzw9hEX/umhr2kB0UFwRd+IFwVAPIwDiz6x9+FGBFkqbVvtME0+DhZ15nTX5PYTsCyDafA8jkB
wkuU83vXs15/yndu9dHwVCcCZoKDRJ8Pqg+G9aLHT3/qUzK70/xMLptfMtCbEmSoysqgEz764kZq
8f/o357lYAPQuAuHYZOQrMeyjuELHzJAwEF0uylfojLCeR4JKYf6NyWeb4WqCgo/Eryw54rLS6GM
0e67H6A4hqTOCSecPcB6c0TLOTZDqCkSGzP+rPBHJVTzufyQ6MZeA9vIJ6YxVzzkggzo7JdcH4pd
F12FWhGxHkwk7iMHimYc2VJl0HhfVqKEoilxScTN1oSZ76ZvD/80uipNbtibNcJApTQvQ1QIZhXM
/g8lH5+V7pDcynQHvKVB9H4q7I2olVeHrVt/7FVi4vXfm2coJ4PYtbZ7HrecoToOXEd42Qqes0dV
IofQmocf49xStJ4NC+/Y6YdfvQNiekb5sVEePhVFPE4vMaUZpGo8OezVTkhP2nS49BOT3oNAJNLn
2sdW2TExtJuldBMsopRF1zgS1D0RPyRZlVWJ3nbG/+add92sLxwHoRD9U9SDQEIBTmkMiqzKwNWF
UTSb0nEhIh5Fcu6/GR3QY/p7UDdKzhSi0gwiub36TT9E7edJ6uev3xiUUmzyuI+mKlwq+8Y1zLAp
bfDH0YE2maSlVWDJQLoDRVmoMVaZ3S1u+rxIlZw1YX887QNw7TBbqaIgxpg9gVJWZSKJ4Pk9c13G
mJ3QRTtPc0wh/mk5t3xSsHwQiUnOP2JOHQrYnx2nRbgcaEQBD7mb7Ei8hl+SVi3OnbbiocGHyeNt
9VGQ/ohVRvPuyj5bi3XgOA9DC/yv48KSoPgEI/Yx0MXowmVpei5FtrQNWww+BU3H6yNt/1JIBq6n
aU2eMBYqUTni2zqFrSnvd4TwVhP/8FD6Pdk0wN6cbsY/oeD1hL7Vo+1Eb18WNI+C8Z77emEx4GpT
IiEYMQfDSvmS2bgzrnYBZO2EZs+k1XoQMgDfRMACRXLvOKaWh0duUVkjWR8Wl+X1wu4OhPlYJH5u
cUcjJMJzvOmXqi+PcDHnZHMz0HWV+gsA9rm6aeMhIrh1JwSSNsN9UvdqfvzB+2vy5kYRr7e9dhAI
L0ljiQR2fqgrMRdyQZeiQ5nRf9Q0HyL3q4zW8Vf6gLhFlxVX1rnTtM7qkV+VJ2dFQzoTD0o+Rmch
g7koPZZwmohPR1rfs/c0E5nCkeDdAaiqV+mp088JXlbMP8xkCQzklFctcm1qBVNDEn2hbkSlA7CL
sJ4KWOExHjLWzX7gwVRgNWU97KfBnfSn5vxxiymOlULab/3ZPVjTv+xmnKsRPg/9RjvWCSi6NFjQ
26AekOFxZhK/8lCda1tBDu7NMUXJPvVcW3/AbUf/Vw4Lq9UM7YJhVQKHTsEOyESs7j9iQi6OvKHh
LK3bauXDZd3mP/bfU/ZKwbyoxfbZfsZ29pH77hFyH6IY3jPv1++ujR4rUWRQLZVxTX8eMyfq+yiM
54qtPr9rnly9Jp/hRdZ+Hy4SizD1DnJd+TJSvzBmo1D7AojZlEtO1QhME/sxh0O+MUZ1HPO8gbOS
1d6bHDny7vjCvKxqqgaN0iLE8auAc3zbF5yvy3ZzTv2MDDN6CUUEg5K4sZkronCm9uE0V7pnoR5E
4fwJZmcSknQryy6Fj3F5e4RE1XWrSCEwG+YalKGyL0A6mm1I3lGUdgwqGj1aPAWN1cyezvzLgGbb
ZkPkxByV32tS1n2kVp/2fJf7TcRlJNODEiWsN+zuav664woAGUeIGGNuZkR4Sdjq3I1Pv9xNkUc5
9odwxt0gUK9LoAfvDE7w1Jeq4f6BSSqzMK+5CghT/MvsX1qf9lhqZH340iMoN/gm0JKxHwdqIsWz
7dRiW8QoQ2dQ7vra5GxO8YMa0UIkDaX1KTcg/Du36/OHca2XyojzutO221wVgU39EZrQYCJpkNVI
oQDDTpZXtHOHWhq9nPIl3xs9Hh0GU6VinUllsDtGtxGHDomvySCkpv96mAfu7CRFX1gRDhX83EDB
Q8T0QVGFcGSYY0Z6WhrfbbotJyhAy2lUhWiahX79yOuYZuJShuEJuYw+hEATCwyMoWyagPpQj/NQ
fShW1zhUg+qfgBcKNZwJU+t9I6OFUdPGmyx2G+vJxcEB6jZ56bv1cD6MT2w3oMu66PKketAZuV+A
dusFoyKgpX/drddhHPD/oamO+/FSOz/HFuifm6i0GBtBmxv8IgVwMa9B5/xXyqNPCb81pUFLy1oU
NAxv4Gr8pkTrz0g/xGUQQekr712R2OtjZFXvxX0VzcQYchVy0DaQ8W8BPqOXCQq4vGSQm1smarXq
8ZR0cdZ5IaBsxNYXrayJYIflcxrdzEonFSq2t//lVAlR3l4nC4GRcKl6giAHYbonmf6gGKzVPRRx
9KszFNhSAOs496vFZi6p3K6jGZ/yM5bOm3dx5+lH/Th0NTYYKaSYaIRkiLEf4ceJ7BV2KBXKgyiE
wPPjsINwHGIWxx/T1iPQRfNSILD7CeM9mBunRJuDFHXjvHfFsa8EJiRKJr2EKSyfRmsVCycv0mON
Lehs37kn+eHcIGWYb5Cvt49xQyLSOMJfoY1bk/K61JE8KoY4ImmbfTtA7yqEr1yEgnTmKvzpgf7D
DxFbptj4/V9r4t6XT3NC2ONaBmgS3GYVk6eKfZpTZRRwj526J6IxgTgEYxN1P3U5sGv7M4zX9zzq
I/Fh7vjHmVxRrLHGo0ehe8wpsf1rsukb6110qWuqF4BkT0q8wSuHUFSZTp86dWXe2Vi6F8GvCA7V
PCcpyixFPH6NoI2eJ5oPCQVuU5q4Z4jd1dnqkxjdp0RNO/W+cBT3zkfMTAAla4OCmLeOjBvQdTHg
09I63oKjy0Y+LjpfKEM8sRprZAhNtC+1v8pktgmB2a3fQsZsAuxVEIjc95TKU97ut9LdhcwpXvuv
w5pDpFbacDp/cQAr91huxkQFn7ILCJx+pi7pths9W3CCKomGWMqddXbPuWPO31ZR+WS3Q1J0Rbi1
WsyADjdF/dagV0DXoXWD+CDaPLoNzwXy2KetqyeZMPmTt1e65jQVDp/zsLgK6CV7So1Om8p6/L5D
ORsxFAqgeZ3o/wfd4dQhPAPTWaqWAxoSHoDRt/P0aZGHsixxZ4t+OasMmwLr2Hy63bNBU3bhcD60
Qj8u3eZsr0N8Alm2hIqbh8kXSorwTXTPjGUl2hTcRQ5nkMV2SauL4dz5nOKRbk6xrTsvU87K7WvE
Rw5tz+X6Diuok3R6PQKlmI61tt5OKGQ6/pP0Q8Ot+yRDM+ZAZhj0fO/w1Yj9hTil6QIXbc2QxUaY
LQg9iKUKv2wY5rz68ehe9pB/UleY5NztbPDHGHjsx8lzQNeOlxKHcP18dxnSFw/mb1Iw2tDkOW/7
CjYPmWN1X0xxP3/AaaHzcEJsofgtqUuTy5/MLSW+ldkaenuf9+fZ0cKwvR4+qF7NQdl8h9gP2M6I
TI1Berml2Hzn27t3ImjIOguRFodVhLMD3iVsm6FKGAXp+nO0t+n3z7FLYFaiAryDcvrw6exqQPiy
VhLVaBjzkcYR2eU1t6fo+bei652wyfelZnyzR+8TUesm6xv8M9DhfANmdf9imXRbSf5pZP3BvzYR
3SZ8smVqbVrU94sSv5Bx8oDOmSPLc100zzFveJgr2+fExiNDbNisrowbiYAiUwEs/3fBBrAzo+yH
PEITPpejLU0TbgwBwsiaIBFs1vAkw2pOi/gTCB21u/0BYDJLyqRbspdaHJ8chRXd6SuslF1lR+xQ
FPndJ+AthXMpb9MazT4IXWOkE5PtuoCCVP9NylQo75mpsM7V6ZqMbyRhCxQxYvhUVmcDtfAoxHnJ
Bj6BzhxatTGLs6fuITrCcoIHMgA5CJhDnHMNl4oJNEJMghLjk86xOd67aBFU6emclgcHiW6ceJ8/
WmkhIjyPUAl1FaVW6an1VO3mPHxoXJwohuP3wZHxIw84fRtsPl6TGJM+0bolDCVv5PZwMQi8+Zm5
CZ2m+G6MHu1e3h0U40zGxfosSRcizfY/VV+yU1RKB2w1pNslRTSve4/QhOx5/th9RfjBw4kC23wB
ZfX3ZsGNCvNVRb7ufhiAT92eU1prgKOrCV4c4Hq64bAE8yrjUFxNazipA+IRxvchmifXczu83dAq
IUrvyYM1cSqyT9+SOqFHxDLKvRGkmJUwVwgxoleo1eqQcDaouz0eoSOsD8yIL4sEYxdI854oWPDz
zpCws6iTwXL77y0PBsO/6AP4aFFjhBX+1NA2tYTGZ32qKg10hAVxcImxruo2AN8H9VnJk1ZGJDdT
fIZq0gxNnx5GHbuMH3kd2fMaiVB+BqLKmGTvj31abf/nRs9w94AAkm+l3iMyqNpZIBMan2attX+g
58SuB1oQrHVVDhTmpDxx1tPFHqXYPJcHUNmmPJV1yd0zMqZQJgTV8ZWjGSZuOiDxQQiLuTunbokh
YWm3ozvVOK4TQYCqrFhtATlxGgUtFRwu0eqSfbShhFJ4dg2SNwBAKgwOBwGDiQLWEnCTG5cbCFrQ
PRpCl0m2gGRWMM3HU49Bq724pP/eSnWqPOM3XcWVJAtJqtHpbyexRrwteZlP5DsrTbwj5E+5laAV
Pi19agnwMUxg3/4zzXZOJdsYRn2txQP1CV4JdXda57vBLX7KRa3Jh0FIcyv9WpGTm1OHxdI4aj/D
khj4fNVIDaJNsez6LJT2PZVN9rpX1AZvL1mOh7LebUWeywho1QxabrM27uSdO7bUK2VQlc4pPCgq
7heiYDudKznCE4bp5ORlC89AoTrzhPfbzCgx7YyT+il1bnVXACZvGfCB3+3nm+CvedDh/GQ28bID
BYma1ySxI4w5dlRO2kosJxHHaCy8EHZdu/wNOO18Jv0wJdVAOMPjJEewz+zVkBw5Mnabn3d/SMSP
NT/doaUk44gqIMe9vuMHhAwWVN9xuU7OtIMjNWSv9hC5GL5S4YjsHcKHcvb8VpKKXOQ/DhA7f//d
qi4Q2APocW10WXZK636M6ImoYxK+aa6xyzlkv2PBMeON9rcGilDYDF0KygVtyyhPaFK+xGKF1Ggs
N7aN5LcDaDriYk/wnFByZIWlcKaU7gTdJuXpwSPLeOs+EGgwY5fBPBcKieeoF/h/9pqKC7ANsEdc
i8CrftHJMO1CHmbpBCKbMacQneil/j4D3nwBFn5wMhY5ap3dIfhb6S5Mh4RJT1TWYS4ECdXxRuCt
FprP4Spmg0TvQydhiIevUPAK5h2jZMmca7eSa69FmsCBA4F1wC4pxoIzW3otokRTSbdh9oTZCJbZ
a+bdJyaFNY86eeflrDYagHHjC/hWdgXvb7QdHOGQ/oIhpaMPzj+yAhu+c/ALR0L+SUdbShfWQfb4
naerq/m9/hmVN0w78ubE/hZvWeK3oI4d3zXMflmgXKssQ/kP6++5Al0Q+S8RgLq/lhj/oO6OtXVY
j/5lcqxqEE3u4oHJaq5AWgMikJYaTYhVJ55DMCtsQr7+SyT3oZO7O5QA3IyUnlzV+V4oUGNgWWLl
u6Pcbu8vwd9H8PwbH2EVs0+Ptdf6nocN+zDRHvNmGHdZJ2XaBfX26/eJ8Jb0ysr0f9p69qy9XLe2
LmuHmTtt2UMPyXXP4+IXsCp+HBspMH5fmLSoS+e5RgzXDzXhkrz3Befc4qvL0b+zJdFwES0Rjaay
+slVN+V51cMbu1WVf1v/mV/k0JnzE5lBMNPLWmODhda4Rmj0hq1XPer2BLmd3sTegMEXacKDVR1Z
OxlKrSdB8Ra9/ITua383PLj/2HbznzRUh+ssngyFGWQ5rmvjJuP160PkE0KO8O4AqjDUoh3QF6yc
qq1cobXtLlnOukIzkq+9U6HwPayL+Qm4xMDQk1dhltTzb12YIth0uOLqrrLhP4R3YN6so4W+ATfd
aEDJvcNk/pZ+QzoJKeDskp45XfZXknC5B0dhgjPRozRCo9S7Xizl/Rp/tMYX8Y4gzr84soyypsXA
G+NCYw4LdHUDtaaA6G6IoVBhIOsDrG6NizSerGc0A3uJmDuZ7CbAUHtoLWNyN5JlFaJ2ixWCG5sH
v6OiFisX2BumV6yRoL1qzo7TCml3/ILLcQqxU7YF9jI4Q9CA3fgODvdISBFXO1dZDiYF9Qb1FgRA
Iolo88ah06oMeSUM95A5a7iVGnzX8j52hmay0MUt94pYuKps4vn4WwErz+WQN0hfvHcaPz8SmibR
9jZQNNel5WPnNbHFEMQIlrlU807xLnS7EAWemq+uwwfUntEGv8GMwrfjewB5Kjz3rNUH52Jxso0p
Lw0Io6z2Zf7Zv+8R5XJmeKYL31JTDZ3myN0kXYo9zucxqLyqA5XGXdf5MaodGqIUSkYVqRYtEoTu
3aiOoUFF95P2mV9GRpcjOgPeBF9Rzwa6Dn+O02rK+8WSWkvxQtmQmMxs0L4beS9Q0VJPl01RuanQ
RX6jgqXMG/DNUQmsZs8fSSQ2cm+kQAyQCzLo4IHtBwjidb5EdvWFAkqMl88hpUfyrjM+cBdSNca4
pmu7jrPiopkldR5gqLFqpBoJQy0ofv76CTyv2XCrQ3wrYRX9m/gJDPs/RUQvJ9c8fzjYEt1zZkhI
SHmFRx+/lWbno2DOq7wXPqfXD13/+wY3Tp5xykFxIr+yEFf0GSuybdNmY2msjrZQ4M+emqCjhs/E
kavKq7aALuqQSRbb95h20aink8OhXtBvGvzJQafUdjqUbw8sote4HHQuiQNIudIN9Tc3dkiZLu8w
CfFPmOiPbLTGFM6z3Eo4N5JhkDKRTAcxWY8ar+lgupJhYguzwBHIjtrl8BHlfV+JMg51givHEExY
s2ppOnB9CIPQNeSABUquH2mOOyrhVDNRO5v+ckm7JGWjn+uxj/SMjYOjonOYWx8By2m6GL/OO6BG
a3Bzs2vPHHHhi3Q1CvDLDt5ieG5XprnBlROj5bhHEPSXi3SGomGhwaTT5SX+BuvTr8wA6nSn9pnP
2iI73yKHQ0vdX76GYjgds2Z6is6YeGxJr8r3ZisSU2Y/jQZCJs+lBusGZ7Fg7WTuZVkSopU+KTIg
ufDLzwoyGYgaGxXUTUtejVwVJn3kwe6CD78iPgiSJ2uXeVcGDUjJlF0uwp33Ye74yldN+PTbt0MO
1I5QJOCa/8URDd6g8qqa7nGMXze+FXtg/hOiKFUroktcALTe3KziKqELpCQaTVACZq/n6f3fyy/w
obqDUrBCaO5Hv9sfmPbgKgbGeFoDtHwGq2qgWkBIXMsC0ToRhp1nUdHEfaNHbZJvILN0512vyDy2
g16ujev106vN+TCh0xIOqEy5Thc9dxxZ63JzHINgquCgEoBYjPVGo02pQVR6BkrHC1BFMbbjR2zQ
nv5UK0mEwdbirB6flaa+MPaUWD8S3/c6lxjHw3/Xr9bRBEHavVFIu/b6KZkVkU3bKBc0mt56nL6X
I9SJjVbCTt2qdd3d7Ltf0ySQyhjXb3wNxUV9kJFauIUX5m3QCyZxRkhq1HvrIxVxiqdGDC/bckig
yHps/pWeP7StJHC7L8tM8phR3lOhdc/W1ON2DVRO57DGxXV65SrAcfqfYp9RYan+2OQPVNb+NIYr
0trILCtTWM8iBqUcVv5umN+oWKU4Xrnw6hxnOC8fHWDA2fuwGxcSf+Nn5Z1ezEpVEhx9f3QSY+Lm
vbItyYHpF59Z7be9TUSTqc/g+XYBKdTdpptshJhZq4uNecKyl+o7SP7ucvc8yal5AmjEzO86xQWh
IvLnxYxAfMlse48/NCZwpwyX+Yzrr2fiJiBh/75+uNqFqncygBdbko1qVcUHJplRjqpnHJUY5QEJ
hWWE5RBdYidH0T0Q8DvEBTSAcH69NzolzWPrzFIyYq+lvvF9r/3GVzfaGouOf1buh6+ku7hZP5IT
4JzGd24tVVHJscavVt6ax1OM2upBSAehjVCQBYWUWHibrTDEKtLlzkdShW2Na+QXwJVS8HMUil9A
GMHNrzMPEjqpy4MFCKL6YDdoRj50q0wO+YCwtcbXBPHyKSEx/S/mNXQuFjtuIQ++KZcafdpSTKJL
FhxM/KKOSzf1GnsPIsPx45PmULTWmRiZMDkBEKOBO1t2h1+UAJnuU4GU4bN5uFaPR+uYWiQcdFgd
JZNyrY0iFvIKDs/w8j0Mo6jG9RvNGUirCQsXHfsPWJ66Xs5cQkHs0W2DzIMi6JKYZg22hVv3Lo5d
J5gqDsJL3AS7b+i3GdbYUjPwpONuu7pNHe5/GsZMwGDkTuRo7pbPs2Oh1zYpP2LN0pSseIZZnmP+
yfzCMTLB6RLkVzFN86xvRk/3YdV4VvklZGja3bZgWJlk88NxJith2x3EEzNWxxNWvDi1pxPvE/18
+fDuKjvC97c/1owJn7C4ZP4+UUzIxh5/25pcdKR9DoF1oUbOdhpScCuMZydsDEq7zL4GR/54qnf+
7ab4BHyUto0nua/NCo/FMzNSPv0oep716pWd7AKJxVjvXmJpXk8xJxEzz365I8sfx/OuV583my+T
/ufmojtIwPWdnqhh4xoWFvyrqB31Wh3ejWjn5hKhh6kmGuMQdcmKtEFqCLJXKcj+3AtTRDRpCux9
1kk5F9kuLkHUUxcbjyZVZmXxBz95mHmut3Na3+pjfzzT+aI/5h/ivQBPL2m5AitzC4CvNx/od7JS
DjI1hYgKiOHsyR8kywVU2RKIHCE5oIIOwCVF5DQBDZKeg0SsE56d1ZEo3nYNP7mDVSVYkAlbsHA+
Kx9HrH3vgW4jrNrbUX5z0gFQs7oK99sscB9AtFo7c5VQpq+jjF0i/OSTEF0q6WUvGBI40QaG8vxp
ca99FudKMSyEXYaw8p5Q2SvdDuwVjnk4IOh8K2bOUBE/NCikL3916ruFAUqDkBXD7xawEOR7B84F
g3qbfSUj3hvqFMpOUeg3Qy/Gjf8aaipCIb6knAWpWV1Jlha/DDP9YoSImtRyfa2YP6xfEFz/XaBt
UPO2xiFZQ7W+HMKEh8wGnbUZMq9xx6oj8Nkxp8T1WxTzBWZX19Q+URW1n3PtZjSP/5OOpghvedBm
DhsAvZ6S65tpejD7BDys+5k7aSCCGvq+BlaODDEXRRBUo7WEYeNFVn4Ql0OlHCUStiFigP2Hmw8y
AFU0r/675IWqKnrrejoTyb8saS8ROxMETQGPIgp1ni7I23wg+cmfDkUTwFSIGN60EKGBlPJD9rYZ
byYiXbzRWgswXN6mRLJzks6CQtZOfNMoTjFzBBtcMi5d7nQFkGZhiitN9Vp3eeonu2ovJi+7V9d4
+2kqumdvqWrm0CSN9jBWHwmmkm2V0RoGoiMrEn+c1rXZmUE/5vsgQHdezXOGgFgEzkgWazM9YsS4
nHQ5S6WegzNFkGh1Qb09bASCtLA8S/x1/1ntGK7pIOx6nRPUUAyJKf1fgx1XYtqjHKUxj6/ahYTf
IPF6gAR9dojvAnRnJX6xHyWH3yQx0n2gkmdBmmjWtJk0pP/rt1HWxY0trf6evN4xVONr1LuKzJ57
w8NjWsM0XU7RQLX7nPihsWqgis23TxvWJkBc6n2jHL9C6c+pS+hSdgoqKbic7dT0B7hSsZSVlJHQ
ethYir6X6iiV7FgYoX8MOZnBpAuO9XanToMcQJBgOL8XULo2sNrjyCw+DgfZ2fe66PQyBQ142Rms
zAX1htRV8YZx0KrW5PO6xaBBMgdfMTVbBRofLily8lYWjeA0APkk5A9wdayiLWSY3Wy9yVWSQlux
kggB0xmMtc34yffirIW1y1fqQoazkGlguIkoxXp0vpALDKrF6AFys6Xd7MaxbIk0Xms7KXgfq6C6
fijFf7t1do0DGIsm/4w6pgkTsg0QEsb5vTLkOFjkU5xztpJTMacfD0k6bLJFPX8/T/wc9AhKyV21
8fsxy7jcV/COPSZ02aLoqsOHQmQwtYqGXpjCYY5LPIkYSrjV0k4bItp05VvBFdioT63UBprcFbzB
NUYkSQqM2UzDudAWM/BJq7rPoQejzDET6BZnOIu9Rur0AGbNfxc/LZCjEL38gujUMnHY7v5uXwzQ
+4pvogHhVN5dssFj5HRxql89Dsq/e5oO2SjFdEKGQMEpcWJPOsTT8q+PABVyO5I9ShqB4dW5bAhu
YM+0Ol57eroEuk2ngGZX8SAvbJZhEJX/z2Of0jTYgBR8ItNN+QjNGuARuo1RvGNFZyyDNrwbeJXl
woQ9yOAvARfPqNfcan7ndJHTW8bA93pudQcRUUb5Ls1RGiPMfestrpnFEgUgyU9AmsuAOIZXLZtV
IYAaFMbydUv6O6l691FITiWi2qpQLPKl5d5XbzyooqLOZ+0xamsGKdUU3n41duSo6eZqu5rukWTG
0uupvZak3NWZ4zud0MyrNn0nVRWTixZ9odzUOz8V7MmCpx4BDIo8U7+hLnidAdQcCfyGBIPiL2iX
pljrT/07MBFvX9ywKyapiszJ2uc8NnQ3G0KTXQQc+pE0OUAcGPk8jGTuf/wKLD+A/SdQ8TistRI5
sWlZYq/tQbfWCfJiZ+D5vTC9G7vYrUDVDeLYTOLQ63FHKjGxVG3Ug8WVNki8VvyRa1XdqyH9p8k/
564I0s1ohjK0dgEFi76hj7Rw0AteKrvqOQpAERoe4xXX9/HylzNPUAVXFqpvhUjBaIM1+saOkmPz
opR5ljO41mUroVWuik5c8SrydkXjvkuZlRLEU8ShLWmiuOVlEUghaOA/TLn7dTfAFQ/Ivh4pp5+b
Q5VI7Z+b/3SBiWPnYAUHiYtQhv8a0zjSkyhCag53wVXedr6S1QCHtF+DZmTkiNBgXQWE9Bk2PqSa
muza8x8kgIbFq7TD+ntFlzJrthPJFg2zWHPqB6F6Fobf3KHD/kFgL5dz7AhIugRAgDetZvC7ZzQm
ipigMET/tmPvEWBlE0dFX+QAtPTQ/O6RODXC+9EW60LgJKzN6POy9fuqarWNQXKKS/vUTugvsb1O
9b8CaLG2QgheJWurUGYc4l7HKbmfFzkYuoxgx1CNNRGOkEZAAo0hjMmpw4W4T/+117XUsoYZxF0j
kozHeTUqk8E8f0Hu5E1Ge4eQBx1R7QJ8GpRgQkqPaZ9+qcPYP47U9DJHFSZk2F8XAQC9kLc4Wy5N
GuJ1WaI3DkxKzcDJCTWEtuMkwE96aUxuyrwJSCGPKnCWXpdUf3KxJ1ERaGiaxuFg/MxlSvLc9csl
Hx5YvzE/L7Npn5szQMHS6rCHNUi1sYhxCyGkTlR+RUopeAz0rGTDQIBnTCHh4J2zZJ84QfdYrHjn
8329Ay1CBWI7h7wWa0Cqbb4+5tKd/uCJj4b+2TEjbv+RwRV0bQIeQwdicyjO+wVxEaL1GTkrmyAg
xmpOA6ZChLG8GAhdUhOV9iJYGO1PlzEJt2XINJEtqxgsnqvqkQyhBWiiv2h9n9vTqhPnN7eGt5kJ
iKiyDWlfmGtn74PkydImNsvFQ2ckooNEZ38UjL11319BOLsCi+txtWhs9+TiZCdmV2+SwV16CGdg
C6Ikp2TjCGyJhNVxfJ/tSc+2gTXgV4N3o41XaNqx6sCz/K+A5en+chfJYb1nJ2R03vk3pAipUlIi
j/nC+dLTi1FnN2tUv8v7gyrf6ku15IQ86i1kOUGoq6vHbFjzrmFbbBqhcJBs3DrrpgWOKYprtJAG
zVaY7f2QsvjYifjl9Ba/haviDQqASizqizIQxH7qHRWuOlSnOsS3HSq3R+bRvSPEoj9B1UF9KeZG
fpapBEcpSzr6//j5Hq/ZAA03bmzMqfJSYHefY0bElA8J6Ev6pbw20nxHshFl4FbvJfGnETtgt+wg
JRxRv/yRMTnQfyjiymlsgxXxOj4LEQz3vZJ9GW7cV1j7KTlyOdIJZoPySQjrcJoXV0CzgUKz09mu
ZejT6QzD3V9S7As/TVWx0WDlV6yIYy7sl3fxnJa4tz3H7HiqftMxp03iqtnPdJw/MRQBNtzyDi4S
DJFRT9yyMVyYLiV5eSyGTETNcPRWbOLvn/o/tYMi2mbZuugGRX55lZ1g+UuZKJVn0baHwKQVh/nN
VdKo+tpUxbFZSPs/bjl89u2o2OH1U3dmES8iizye4gw3Qyxl7Gh84BUEYRmeHoQC6Ryqpj6EoQYv
i9DjIBWiDkg5E2fxbJnzbddmpkvzaU0SC4kbcPR3Pqxzifl8BUpazTAbaU3LGsbSvVYR3lHwytnq
ZWDBHWpk8XI3Hk6EX78XkoxHWOlfzQJa6/zO6etr1RjLwj9HPpE3YQ1m2jBqkYqeABKPyq32Jzr2
f2vxItffLC5QdnZp8VcqSuU19Zoj//D9XzEVy3RkC3jtlEqB2+l8aEbbo8eg9gm/fX8Mz69/QQsm
Wix0phzWZXY0Lf5+NuFLG6ssaMDCsst8pTYkghRh09vOLb+mydqq85HQ+kcWwyiv4/RevP96WRsW
9/9P6FRdmD+1JGJhktoIJlSGqMJjYewsKjNgjwr/5ZX+xpZ/0+Ir2+EP0L34nRFWzfU8jVkkxrCL
R+zwl+mSRIdxjagl53VtbtiqAmVGUgvOKRT1In8hLxu9ST1RFiKKMrqXAhJLwavkejCg4S1E919P
tvL2qyU+zeYd+mENH0W9TADmZxhxxBtNp2s54dEQvi8HSa40RlrCa1YEjmDVUQx1hUokFs17r3BC
MKS1lMtvP9tZO/ESGbiWbTdd8Nc1XfyceHPFomGcZg0Z9Kd9eL7Z61fw3ckFep2b7s/dyaxWgB/0
onMeu7xp7W4bsZcFkKhvAxbKG3AoIkFDrBuAIQyftNZkR4zevVRuY4IKi/ENbqcBL9NvW8eDKRrh
ivmmhO1L6khn0UloZRKbeb//S0Hn1RB57HiZDDLKaX0VirF72OZwjlO6ebxX35ISD2J5nbzKCrD9
SdAw3X3nDJLNUsOb49DniMCeyNGsxlKeRV6lcxX9cxI5pcgFAC9+67+T+PS/TqhDVgFFZcoZ7FgY
jDnrnbJuinrGTF3qHeqfaxSQzE4QkAD37jRVrf41KZ9ulLhjAbrZUnvUWu/mQ4neujwQSZiNOtPG
Pp+jomHlMXFSjU4MOYF7XziGKM50cA1Lbd6DRjJEyLGIjycN4qDIXDUyN9hYVWL1X2NrLXdNVasL
OjhUqSPTxh+t5rVoLXGCiQ/trKdu3RH/hq0W76AJjdxatrxv7fCWXu8v0YqsxrilhkgvJ/QlIjjj
A9T+0w0SMJebpbPA9AnHKnMCg94Ga7O7i6vzO2PQxOrq3BVVk/rG1WA2hxZXcMY8uE9w5XnA56GO
4uDpk6P9bAb7yI/1tO9wwoOLjRgO/F7eKd8wlKNA6XAzW6zo2mV62ivG5we76V8Gqc81j+SPDVV1
R2cxnmrBP28MZPhfgmil5lhKZ8NlbshHjJC/r5T0V7j9Yvkzdvnrrld2OUWWTXap0Et3y9G5ngUY
1ACp8cvJ7KIDtn2tr49aX8DtU32EblvyjawforCamM4BCLIAFa5t/7gNhbEp9Nla2bWY9rY7ddbE
aXsiipuIPU7/w5h8HYjWbo2cDCzHoM8FkD5uD+VG3JvHfeiQLswCKxfV8bXtRl+I0hJ7YyKANtrA
uay9dpt1OW62QAN4b4x0KyrrE8h3j5Zpy1lIAL2jGCUgwY+C7tckPW6S3GmMfyb6PAJLd4XTPZx9
uekDZsJH55crz2K0xIKPjdwRnDmULRgaCPttWKZxSnKzS8G/xfg2O6lstaSGITa21R6Ex2He6Psu
FAqyFz4pGlHUfBOq+usoRprKkzAOUCtbi2dVi8wHYJ55dAaGk5ntm9f7GEBSJTxqPrdJ0WvpJ5TE
3KdGX9GAPPDNOIViUDJutZXzjYa2CS6EqGfzT99aZqm7I7q8gEtXhrr3d7wmU/pgniwF1T6HfOn8
+PDDWM1sIMidsLLawWL1z4WIh/fH6rrY/4BSDhEpcBmVZEyMslSnJlLXZbnclkiHEapZe/kDtJoo
xGStQZQJmrPJRxAzbnUOIsn9id7b7ZXtO5dYvoheuuDxZ+OqgwDtVjdpDd7qcRYEu8lLeRiDkKYs
2jXG78GfrMXW9p0k2FV5R2e9I1CGdFPeJMDY0kFOf1ziz21U9a8QnGDBGBhXRln1FaFWz7kSIiMn
bzyhanNnGUUvus4p8lYgXFuzmm6glrkQ5Wyk7mz5b6Qc0vIwwg+kf5J7mRVLULSa4uO0Amwf6FjV
uLVIG4FdTPMof78QqPU60nrXYf0Ubvka/8dMkKLbR49+xx9xIGh/UYjKnL1LYdIneV6Hab0rov3v
IEHGc2VmKt+tOO9ozFcU6QrrDts+uFmzCUtX+1NIKyUDALa706u+cpcLEw/BXx3rEX6RfZO/D7oQ
TBbNaBmMg3IUrIyLaRsn1i71GZnHqosKnqjS2kW2sOmLhZ5URi0MPyAiI0nVoehoFKaS7x8lRRzG
adPKU1uWhGls/JLx4jJWeSpeqJxwaxoZ1XwtS7Hn3OQqqG+DDpoKN3Q7wYJcB7zI+FcfCaac6GFa
+Be1laIICkyOuZQyW0NtENGT5DJOcy3dKnplwCoiDzZxTuq7DRfXDsYloG1IdNAOmtYNUNJBo5Fx
FpFt7eG+O0dRNdKo0HdkMWt2Z/ozj/ltc+7SNnLBF7uYAc9N9jZPY4IFLA8WoK8XImwUebSHhbo/
tPiOWXR+ojpVNXWsIDNdeMoq0knyuyW4ekGT5lqvensxU+7a7RmDPGpFROeQ/65qxEBr02mwINTc
REsg6Se0BM40xkxthjNE4BeKc1k+GCjsIM/vq3AEj1cgqKF9BNxcERgqRlLPfcNn2fqMfeIpfqBb
EUKQ+CVYBaDMWiwWzU5/rfKJekekOVXeKPgGoIwStYUNdR9lHHJpS48rVDGUB1sQ4BrPNy9+S8cF
ppNITRJSXCf1vYYgn+ZQ/vC1/mkcDMb/HF5DONsrItmApvJQuSNsqk82Za7w7t2rkYfLHb60tptK
5S+zPtvHjy/44FchbP5Tk9JNjcPboCW5j+6uKb7uLN3hXoiEeUepGjHRVMsZHhQQQ8tmh1GPk9HV
7RTcn7LpfOjjW2eYJpINboWTVv23epJcbbynP/wePOxKN6dX7PhUBnx92la6I+miQTsXju6onq1V
5WK+3fnlFKKMop3dyFI08v3ZeMEenVw39sAvTr1RcNJYZCLxFkTd1kFQzYPwncbGrE+X90jBJ3Gd
D1JCWmqj3GPMadiPhQQ39V+6QXMd3m3B1hoDLEPLUJOssCeIsa5gjMFhrHg7yzij/nGm6n9lszYp
G9OuvoEQmcmgOxUzLxRcAO5t1ff+67OepHeNczg3HHXcbaPVq6AV02iiYJTu5wNdiBAJVOZAnoXA
aiK9l390cxumNl6qxIyvcGDWwgtQyGd1eAUOpW185CpizWosyDN3m7lnFJ6alKWfKnMTwqkGh0N+
8PTzMJUOLBHLgaG3DpiQOlQRxhc7+BP6nBNuDPzntQsC8sUsFspiK4Og1kHi+RylbpW4J1JnhSfx
cSvdJm4vqSVvgaaD9XNBZ3vl7h80yt7sZ3UkgYMBZYOdA1YqJpNU29JgGXse7yZlRTvBfq43t4rj
vS+RNJ7+lW4jwz/R04xKBo1kJlaVqqdZ4/4/VQWU676KMkC7+pc2aRd1IvjeVdoB4llZg21lxBuy
PrS11EHDE2sPGdoGAz3Ov93Rm6cvjAGW1OMtYSu3poyYZSD7I1pj7brD6aj0fKtTMkuUHKUQhX8e
JkU3aXtLZPSSm9ABNIrb23IYsk5ifBAfBcirWd3O37flVtdbOIXZ1LeGC9iDZlZpPRfKjxxjR3IW
SensffGHLBgfAomnG7oBOWuh5FwqT/1weOydz7mszi8c4js5ZTpSITJlS6PMuuELDb/BD8bwsxAf
fC6uYmxeYhFWCuW/W7A1X3ZAF3VMv5dNw3n1gVtbR2zkVTIrq1t0CLwgdNFvBzHl8EQ8KHqVpjcZ
iKFIWXzCLdg3n47hHu6aLKkCunU9l94cujdsGiVrv08j4M/tzRiji5BLQsyAueyqQRnE2cGcI0Qj
U1yXi8Syr4iTy9La5svx4uX/mH/oetiRRpSNY8jL3z1JVgxapkiyrXy/Ux1IWQYfGbLudX5OHsce
4HoFG5mO9vZce3Dew6RxozbwamLyrQiAjA8Y8iJfXbkh8KXnuzyZypQ2F0yBQgtND6mizpJmsw0q
6DWqVQDsxnOYiwC2R7b6ew9wfxhgztmRhYpzZamVjtRZ747VP6eUWeBiXQiXXc1fQeL6Ub6Ej6we
KVKFEbgBELQatkmnkpRBWHHTOXGpcpB6nO4oSRiaFfwpdK6L/KaygbePTW6IJflStx7+AyZM0/xA
uI+bvG2R3Ee7MFV3dBPC1vdvOQurVT3d6LPfZhgl7HcDF8nBptCONZdR/scKV8LISTOZc5bsBSyA
CQIb2WqlJ02Jeyi76zuFh/qomEG6qp94w7HghU/R1owcF9CVwHf/gI9pX39oBa8700TDcFiqInGD
GAh4ni9CDBK4AiUF9UvSy0SvVtygvGtefW/Pg2W+kjQTAH3Q92NUhgEkok10FcDqhzRuTfSJEZmx
vppdYNFuXOvWjjmic20DZ3wrrS4t444Uclk6s9CyZF8HYhrt8Z57GpAimBiUnj3NackFkDjTg+mJ
mnT4aQZqxRoGTzjK6ZFnur3guacxbb2ch99ob2aHPP2mSvelFfS2DaUKJd6gVKbM9FVasBBlUc5r
RKSEHri+SaS2WmlDJivtN2rcfbMXl4jyubu4k6pXeSrAq0ARGoZPkjDsnTE02u3VPM8tmeeQgrhZ
dSY8dUTN4OWhrTXVth2lo4Ej8dMQcs5KTwvBYgKseRQao9AsIpMIxhyGlcjennzXOacaIaAj9Qe+
i18qqWmezjf4ul0Dio0OVtFjdrRc7OGubV3EGMBjXnhiu1XVIXOfu4Nw2P4Q8mvQIlWryM9J02lQ
FKEUU6oEG+cBvvNq07K9x7Esl7XV6uNsiRk2kDIbYvfMUbYhGyo/cvaaL6LfLGzrMn79lF6Ty7yc
PWY8PKBZKwQ3nGXIVz/UhRyp4h+5sSNJarbarFFMyPXnuyfVMXqrkN6zLO7NACF+Txxykc92W5iE
QoYM2QaFil4fgc5BHqZbkO0ZGDnIybgsJiA31QGcamTUkH746HyrN8qby65Ru0okeiWVK3fMKXWV
qSapH0dkcklrwXcvXwGj2mg4MA5Q0f79qGyVCMclBTq9/Cf6Wqr5dGbgX9M9/cwmBORaLbe2Cr/a
bCqmnkL6ybh0HibiG6yKBgT1lltJsf2OrWnS4tDJuKJMJ5uy1X0KluQnf0lLVkIW42YH9Qx1qY5c
158EGLcSTM6PIpmBLQmMSyi4oTfJ00x67o50dqCBaJ4C8N4WR9prERj9n1t6E4C2hmnvNNu5+mEN
K30CHDZmEWuk8PBLQ4zxYNxrjn7qzSSC3cehjtF6PDGB10eZzK9owDNoLHoYtdzer9p18HYmzO1g
6AUU0Fu1naaaII+7TncwzrdFhCZ2Q3UQlZTHmi4cFjz7k1rV3C8xizQ24a2OdAxnEpZGLoBQ9LLl
5F7GkqpjlvUq6C89QpO30oD4BISEtL4Wubebh4Pj7JTVAyadaScB5quwiF8tzyOAspMDCrAnF6j2
KotPEsSC4Llm7Bo2lWUAxz2cQ+T9VyYd33CrCK/h4VUA3ycEOh+LLdiTtGbKGRmyA+Qqh5+G3zDE
4bsp91K6jdsZWhdZQAdGc29uwINdCbopoMV54Yo+4BtJfiuyKe165j/UNRS8mW++ZU+ZUUnHkFPh
XLysEKKsgIy/SCMQO29Xdggpv2ing2K3VSySG8IBSud2h9kYcc4sFzHa4EnqZ1w/ZtMs3FWecZwi
CWABKcUnzfVpWw1kYFhjwKr9uUHksBnCp4ChgTu9Aj96NZgevxqpqeGZl0S34QGQdmJOp9CcR3Ni
0ffYU1ZDbNmAqk6S0A1Jv3ukbkGvzAUd1m3jkuOuuxFAvv5o6JA5bozV+euES+IwePWgokqS2hK/
nCQQ1vuFsBpVSehlx23Ipn/retL6OFJhCNY7kJlvWxRwGMfmBXBjA74DDgyzuO4SFMCHzTG4txEY
0FVquIVHB4v1KYS8RJgi92uzzD33AotRD25EJwo06mSVTdS3vNPbQrxJxX+joqgS85ZZW3V9HsDq
y7/1UVu9kQrKNnhdlDVw5ZERY5aQOMxjC0Xed0zfWeVk28r7anki9UTsrJgemc+w7bhc9Xwd1qVK
z8fZ8xzYN465jP4QSxJ8S8ZJ8fPYuEQqjxFJcidlzUO2sfjo+M2evYTCAwBqju7bxumtMvYGWJuV
j3d+/tHC838z105AS46jkERp0l8fJkFxbWVcPikx/Td/zyFYnq40v9qatm6KGxXpGuOUZVcwIvF6
SgKW4FJjE5q6p+WJpZ7gSooEF1aoujuAgdxnuShJ9AUrpB0jGZnLZLHis3IcgZ/X7hGBOR4rBmY4
VdpHr4C/vptAG3lsDYEDoKK4WBJxylWB7DRxBa9I9VV+EASyYXhBexKD6AiydUqdztrge4geOJIS
fkDwvRwtVuJyeKf9Q2KWW/EMVuaiW5zxfpN+Iyer1V2xQ+GkXiN8u/w40jijqnOgeFP2na/unLV0
YSv+6Y+/seXanJD3SGzpbxiVW1IcTuZBVgedrMECRixcqiHtekokT9UDD4ECUN/Uq+uWRd4YaCHQ
JugaJp78aJwhMSduDCbtxgQyRZzj2vhVHoZhjy5NhrS7I2fWMR+VZqG3grKiXY89RZKPw3PDBUj8
b4Z2BWsf/8LR7ptrQtpDKglqm9fSLeqQwqJDFkMQfgYNnReFWik3fN2U4CgFxJDumXF8gvZ9GHSL
8xr9neP5fNnRMGItJc07g47DXx9Fhc8DmGMOfIrqhW4770xv+fssxyRvg3T7+fGgyPOqk5/xS5La
BNgPZHl5OShYQdG+YWHGx5yMro20h1qgRm9oW3n6GPofEDW4LNuxDtMz6kxZ7zmG1hBfENctIl6C
WrJfhsK9TQ3WqfLF7F5rorwXfMzMnlS7fapt3ByzEyIv22SvNQDWcLgoUQWn2xt4fg84fUypiyDh
9jroTN1SN1W0VMKEHn7Iy5fG6he9FX9itKRR/B/gHT7pbf/4BG7Gp0vsy08ebEcu5NUSNrXxl6Ye
rDSRRAMVCJlJS4ZOwR6e/kFLwAxyh2T+wp98SU3hbJQPPDqaQmP1bwfE6buhHSCvF4XVtOZXuG+L
Kjzd92jtPFedgZ6spz6ieISJxSEHkCOYYyiWbEv8hF3PGQ6h4qnbaS8jpVKi1EcN/YdDjm6Ph4tG
fAg0LxXfvB61Oeq4lTrLzcRMJC4l01nupl7nodo6DybuCgVQmzuwFY7DE5HyaR0iui4tXjLnpl7s
4XEmDrKijYIAqaCdUHGRbpsnmguUg/PoW8tt4Xdye6KuVoo5JhtOh3UjKOVnAphY9wAcUap4jHWx
Iv9MjVsrfAJTPU0mDNAze+LBuYHalEJrQRtSKhK3+dCoCejqdMZnhw4M7hkNos5JJBiMUrAnIngG
ET0ODDtf0HyfHD7NTh2RuhfepiM/4jFgDmyUmt6Ounq4ceXVrZovuEFVnrglkJo3/xkNNnGlNqtw
Z6vsHAZH8UPcST8grQ7Wg6HnZkmnEXzs4YozlnwjZyfW1usR7cWWF6YD9qdulbF+a4P3cebEfdZB
4o/lEPfmN1H4EL+kPlcahY47aum2spsVw1nXQ9OVKLtq4zJ7CJJRQghosc6pJR6miRBn3oI9INeO
GilbSCTLNJs92upAmogQZc5dlt+4k7/+mwncJ1EHY8Wbn392s+oEZJnjdsXLRX/Z5iT8o4j5I/jj
A9W5PMrzaHz6VLBuLkaUF5Qi5F4kBYukMeAIK45aAzMtsmH5JE5jJjTXlBmyZONWzhVxfi69YHKm
PKYfOvAEBiOX3XphSUnC6EqWgNVrgvJoTkUn5Ub0kzTOWr8jS3UFY8pL1/kuUgvLnHMiHBmQ8xLF
27fBX0pMLvqlZNyiOyHvN9Ey/vEGG1JLHpWFtdfhC4jSHUy4FiK8Henl/c6ZS6rU6M0lfzi2ysil
z+9N2MlBpbEf4iRZv24gii6yedMldlFluz/Y6SgbXnTxJ19+S/+FY/Bfg7rd6ybUosPwivucrzXt
jdMrImg6Xbpgt6sZUnKB8qXof0U21BgR1yjEs+rP/13V8g1AEpqGyTN+1gaS4KemC24ncHUH81EU
98pzsXPqpJDpPc8hH34ZPHw/eFN1dWGD7bPVCQ6W7I9T/gYBeMGQ8Pw+0TJjxnuekaQjqCzpa3RN
1eVShNIq27et8GaEt8b45n7/vElPyIrR5hq410XqDJNDyzQejpoF//TUuWPvSu72EcRDZmAx1DtY
XL2ZPcbqxhBPsdfZC2n3676CrvcYKN8TkiB4tH+tIZlyTpaZd+odgBSmTivA0kridsvwplz0LNAp
SMP8RnNgGsNWLTWnJZ34gQUEK3jsB7ZDIWthZY5xPG/VybHzYhnVSR5HbUlKwxWFcFCL4xtPO2/f
X+6HduIbnsvkj3DM6LCfQJZwZUYf9rU2AO2DvQBvEFd3I5xVGt3J3CHnVr2I9VwfyTkD73u9DkaZ
w+nC/tNMwIfVhc+60MbDos0EjDIcd+mhQ9Km+4TXdVIRS0q+Y3MAYX3NIMJKZdRKTxgny7DaAh6P
pDBWRkZppxnAaqrGsgklsO22NiM1mij2rP5P2K8W72dHE40eEiLOGqHzjJTXSU6PBhoq6JgxPrBz
NjhU2TAgcA0+I6Ji6K5/LETTy9qqw63kXZ5zW+ZgkFCVR0N65Nx14XUHi2jIfKOizjayz0oY5h5J
G83JwJ8UcJL9FbF9+1ZeldQi2xcy7RYX/M1cEfx6Sq7phcuXMtUOqLk9XA/Fyw+xZaY1NVx+5oM8
5ne4J1Vi78hosNKpoZlMgYwcQ2Jz7pY4teAmK3Of23iwbGec1TpSUKBYOPSNbf7Ff4ehDE3YjdQf
Oa3LCxC/3+bhhugLfUSV/7q4OM2jF33m64Cot+CUo6HKlgfAAOjisLKVB6BWP1rgALZjJFyQM2M1
5XG9oVJ1CSzUFaLaeesO5XNY5BahZFK4ruR0K9mHWdiJrAx6F0RQBpLsINLyL6Hv6bwgzkNcUHHU
83+U3/7Q41aZfHsVN7BIYimMPbTIYBVyakRxghL5tzC879kGQR4zHn8rhlxNw+Im6rLfoTvURNwr
Zov03BeTDrJ+sXof4xt+kh36sFgvzo3EucGhbbQmb41jLFLg5JaFJfZvDaLg7GGbIqo8wjpv5iti
8SPC8bmuTqvlYXO/kJxuRpsyDLIOc23pAQ4i8mkIZesk7S7Gkbfo3FS9Rx6RFfrjHPOIN4WtMsN4
0akYke+h8U5w5BpsooiUYBcuUsWCsKncPdfef5KzMi/9lCIjUCTcbJctl+vqb1OYn/YLF9M+Ah+l
TxB6FmqBRbNZECwn7Jc0Gu/qd7FkCcNkobxz28R+zDr72wqBe96B9E6SYtQhVJ0OsFjfUA2F924C
Gpx93XnKmckpeW1cGeQ/YlOolA5GyJjBXyXhs0eVhOA19o3wGc30hUOaUiXmivvAmBu+VkEQN0Vq
mjDCDHr2/fb7d0eaQ8yr/NuAgr9PI/tKoBTeFR7pmeSkcduW1LSiz8t5qxMXG2Qx+Z860jbZKEWi
UZwOtJO1Suu8m4bPfw+PGxu4sEOVazNnCBge1i229xVpam1h/oJBkZlWHbutZd7/5EPqhMMq24yv
Yuj/ucyRHXWzCcFfctFSjefuQ0xwE2Xr1bFrLl5qWshAMKSLbamum2c15mywfA3ZsN8L9EJF0Jdy
OE40nqqs8cOd3HL+pHu5GRQLr4PQDsKtljERdkyi0IKkSURSnz2ETZXbajP3SKF/UDdCHcnvyIRy
Nf1JXbbbVoc69vbSVVoRTGM0iEpKyWJsDulhZpQ/mJ4qMYUT75JZeBuikyNobtk3d4vdzO3ihpCH
TWtbhrrLcLtfB5qnd3/o2J9PGqL3QOY639E/55VZXM+laN8euy5WwXtfEPUS6bHAtEsXf55kyvZc
aqFz3sqYjZwLe8cUQcLnV5gvZ5NM9ZZItq39jRsiBZKZlAunQkLjwhsSzTqqO6Olpd7X98plWwON
Bx6EhLJds2DsWwRTpQA7DP7qxAZO7UmIw+WupFGc8EolUfrCPlbfCgUMPcUMkMgHUgKgv7J2gyqu
lMh1a+FIEoUjq6qRZHV4PcEqq+bITPVPA+h8A8vwWaZEy8HDgkFkq6hbkl2Tu88sPFBk7hgdxkBs
7Gy5uT1rTWtFlcRguO7ox6hvN/sb2tZE0GVd8YKDlBwL5QSuS8tIy9x6jHR/x62xXVrJW6egIisz
4xfKz08AAslE8IjAbmKf9cXNQIR5YA0FhATsSZqV42ULPPlxb7EiToOHrZ0S09yLqNvH/HEj2EfI
V+z5OVdNVDVeBk9cxODbqcRmBPwmthAdvzEOyAhqyz7/IrfxNKR69X+5jba0JWvXpCdo5DKTvC5I
B8w6bAoHVg8J+xLrsBZz4B9FpO8fmuOmg/B984qBIfhbhDm0kjWmC3K7CwoND1yeBVzY0o+8o133
eVNtyvbm/FVdyUW/EZRykaErhMs5ymt6HgElRwdWNcanMDW71rZqmvOSkCAW39Z6cTTPLOz+bEU0
4FMUmc6uIJVJyLExervWRdDGOkHC80ucPPfwGJMTaO94Z6er9CcPwTxpbY+SC0X5SodoiYYn2jdZ
DzaxQY+c/zwUmALgjLtBPKRwrU72X93dPEtehjPcrSpyBKzlm5C/r61RJw/XuJ9mGHoBhFyeii4w
Yxrl1d5eaHQwmKQ9vJ2i3/KrXTSI1QfASIxyiV1+TFEhED3dIFQRFa+5bMz3cdXjlxnx2zjyTgWb
q+xgL3Jecmr0xqC461kDFgNyMLJcXe4wEU8MUvrCi0mdRXI/GmxjbkSHv2uFb+XcxNO9UmTlX0zr
kW53fRUnIqRgP3cqvP4vMd9bQus56DeQiDkKo6DmIW9B4l4rODb4KNCYkjiUqK3sxQ8cZfybc9Wl
19D1DSwOJZLezZw1vPXxbCydJ6fsGLhiMhHQwR0WUwKL6NWqBZwlm51iay7Hmt7xSLjvk3QY9yvk
nGpK9QlOiSecSYdw+KFxKll+ZeLThWMVa64xmMrcyLiDbKIvQ/ZOUjWiBT/mhHaGZXQQSs0ztitP
1DAOB6EdIAlpB7E/5e10XwaXT4TjGtcewfiM9hsB3d3ZXszjOh/9nz+p35Ij3NYOMUcIcyzbmRbN
QyZeGKIjVYTUdVWVyC+UD4jn9b64/tyNfzxSw7lMxG+A0NTwvqBm5AqI2/6Wy4QpYff36LsSMkF6
L0vngSheshSAOYsJ8HRyqqq88QWN+pwlfWQl5R5U84DkaQ4a2/nJElmZha0+j9Pvjlsz5z5f0EBX
ZFfIhJZh6fXmda/juxfMPc8UfOg5oVS16/rbNejw+0XQj2ImxG+oEx3SUJw+e2qBDpLZE9tnd9Ve
a/pz+0RqKzFIJI/As7dRfLyYHNbTjSImCtaa3NwaXaDcovt8xD2LjjXl/HWMn9sYu7gsDp7So8wS
Ii6ntYmMW1vSwFLIbZ+V5wd6/cV5QfTMjNFDNyqsK+1ANgHdCDF3Aok8w4oChSWROgTkP5XVmJGk
3qeuRU4reeisSSA5vFLUN/V5tg1zw9w+AxViGtrWaHe1zVTfmCuTT8H4/C1pnWUH1rqnMvZCughh
4kG3TZrj7QtO/sISoJF08s4G690GitJcXCYcjCCGyb6RHlPJWu/GK3D5GkG7UTZePTW06xcKQaQB
0w1uD8sevMyMaJ13P+l6SBd2kv4bL9CDaR6MHtLMpMg51VUEuA7eZz2o9gyOGPGBVF2lRYHuLI6P
xNDiiKxwPWH/VTydAAOrx3SJTUaT/iAv9N7X79qCPcNB34uTq1K+hAnLz6A7dYynHWMN/dFZLEqH
03ODiDYue1rP4cbmY4hIhWj5hIorfu85AOJZKKjWUsf8rxYvkL80+UCft43jfzBNeIn0/2xjvHgy
oblw8Zh+TVTla8IH4uBuyJSr05suNoUv7hbJ6VD6FtJ1ry4nsS11ndJAe7vNK10ZnypV4kE7rFSW
SoHjclW/yUuwRO8lB2RjG3xAEWmUPoFrPh2WfJZSIsFrDvO/mVTXI8a07M4wxfILdACqz1+pJZJ7
x9/DpCWAhAEP2kByD4/VmkMjMl3+ET4AtmWSEVjnt/XXdkpAS0AfwjCLRmIhu3ALJ1JlyT0CPWl7
AP5Udg4giKAYnlyOkgQ5vaFTGDULsA2QdZ49gcgFEkjgPC+ZVOMqXTAvAJZXfD3W3z7Efs71phWi
0n+ByOvk1KpR31adqA/tuJmh9LIw/r/OuCjNMYA2+qnMUqUwDn+v4a5yNckm0nw+TqkzoGx292F0
780w7sV8Ng1DgmC78H/UmLQ+P9RBczaqfsvQa8aN7Eh1qh9bTjTVJ8Hf/Ml3JrM5SKva4N3RN3fY
uWo1N/8oP8vKxdIN/43LTcVf6/a8yNpWGXPGE8VX/isKsFaikUOpYuv4UpgYsPe9icIf97R/TLS2
ioJv9tHVm31e9vfrTDxf1KLiL+fDTsdiI9e0+xv6UEaZB474Mjxz6TxWgeuJqDeGLk9MBeLrPXlE
m+YUiL4/dxve6dY57pqdm7AJfGU1SKg8rQL3sCxzAAGUIYXzm31AOFnrGprQQ7JkMIxcRIqo7qkz
cCBuFGt+9U7NY3xXZ7+z9vX9KWGyeFwwo8vur8YuivLo86yRIs4Po/yqiNExEZI0hPt7xNJyT8YE
wgciCgQ5+ntCLMiOVx4Khhabpa2kVulthn954i44GLe6xD+pTVcswyn5RYmYW2b1+W0XPR8XPsRz
7j2d5+4fJLEI1aDV6ZluKFB9PSzmgAZ4vnP/U14pAwetxHtNLuoHmphpySRs6kttkrqnBEe8wUaW
xgi8lSRscxMW2lL+Xv/CxGG1Mlx9cosB8EHx8c+yJwBEkBFY8T3y9ErlVM8K9B5kpt1lu6Qr0GMq
Hn824mv0NvSZUk/UF/XEcKAIr6vJi6+7t1KIvW87cbq6KMNb3nIc52JHkznJTOWuB3uADGl0ebQn
wmPi70XgAscYtJtk8MIYZeqDlybH2TRXGDH2XVQEKh52iYm4TScFnWPdzYWzLCrO/D6ft2FqGvBZ
BoTyfAENNjCHc5nDM3IBstK36yQkk+5fsqN9qMBVx37oyMnPs69kBPp5DQt8GkoZ6+GM/iorrwtS
KfggwgBjDlvoCUXofdkSZUY8OQDKCgcxs54OLqDBdgxEar9MA/gln+HHBqQQsc+tgzoZOm+2o4CG
9s10NWWv3PlSpKvjy2Kn+Dao/qkU6YFXdRyzs0S0pcfpRNqjw5FF2ObiAMDEgNCV4gRaLOcbz0BG
uBKvNLXjG7r4dkKc+bOCxOtuzboZgfHIfwlpXlb4OCJ4J9zzFh7uLtJdCTMGrsA6i8u4fnx9hxIi
MvaiPjk2aDW2woxw0psCQsDli91d1m2uvBFzkivaASh673mtpDW8ANCudDMp1KNRPYTkOcuZ8VTP
Eduhsv1Kqwq1Y04RmGoWiv7HJOlh6/w8aLvhHgWEhQs7AV6i+L1QLdPURIYMPN6IQmY3S9qw7w64
+De/UuQo17142P/90p5BFPc8nFYhtMdSyijg83brvsjIjtI19aCdzX2m7+N9Akcjd1MAaW6nLjtp
1efJShkFkr8XBkRdZiQKLm8Z1rFj8WTU/2T2hOU3mskeBnovRXWsoqHFy9NVvfWCn7V6r0JORPyK
XhN42Gic6gfWuz+ZgCYryiKx/saXAFUF+jSPS3Bn1R72nGGxoCXeJZgpOFv7hZgGHl7MsvUF14MX
9A+HoUT9LUQIWTCwQYNqktbny6AzZSSaAIO5ybzr0QLGQ03r6DbMwEfI+3Aj7p1nzA6D6Mj1EOKf
mWGJXf/VTqN17mzZ1DxW+tAfFHRrmUdvtOOw5gh11vy9iCTBDqM2q0bGn1wnY2ss6Mp/+ghmi9jQ
eMIW4HqFZm9ZUOm1HIBvkL3jygNUsq2xsapIQq4goMvK+KWTz/5Y+nQDQWmgqh9BHvb4CVqqoY0W
DkBqctM6kI+tSp5YgQxGBsynLfukkxtxBcpLG9eXCVIkKlKps/fQ5D84en0mXxpOwKMfnR72+eMO
N85DkGd5oEo2PpP7UWW3SfnFpLrXsQpHsEJ7+FAqN8GfX+QJmp8SwMekl8/UI2PzJzpT9fBRHirz
EDZqSgh7R39iwCj6E0t1HzKlOWIsYp06EUyDHEcov3jpH+NiXHC2ycnVPB5Esr5zTmAVrPOJ1x3K
OICqD6t80dsWPJEDnJQOqzuVirPoPoMOrp2k0pA9FvBzeEJ6wV0SKRmWtTbR9d0IxXFCXcdWicGk
hSkqJ2/gRB4MJEoVCv+JylOqoiOkFHcoZO21mXBVufFJQK5s65Mm2c+a0Pt66QKNBhYM9KJhKlC0
vxyVTjg9q/zy1ZgfqMSgJn4/GBWKXHX+guK1DaUhM/mNul55OcBk0SjmHqsSjmRrzLdUooHgnO8i
BS1zvYlb+/xRpc67LdIKfL66SsevWNKnZsq5S7haTwf5I718HwvPhp7b4NCNz81xdvnI8idcTD5F
03hYh9kGHlGQHtRopFbQ8gjTK5fL+s9UJbhHKINckbOlKhnsfooHeJYqyRM953vazzcUxl1sRlQB
yTHrHhTC78VV2ojRuDxNFxKVUe6dQQNoSA7J1oCtpqAvU+DFZrqrNzSr6gux0N87u4DqhZ7b3zjW
rGTH1otXjiQoCUsP8nRt6+1tbLRkguhYi6YgXsYBdfdLF559pzgWB/7clgq73a8nfu3eG4e5V3WR
DZVTArw5ft1z3uB/VQ0PWxbMLUjrX6i4mttnlZkYU2U+xuSZT41A0VI27vIynDNa7ZrN7vCIe3k9
gmizS9apdplE8KYb5vFJYgT2O7Yu7xiwGlGbjqiJc3TluzNFebzYJdhrvejO0T4uGrIfNzLGIsxH
7scMd+fOXy9wH48Nw7cK+zDaTq7jTNEbMEnQ85jkjMT3lgrrm37wwtolL+7szNfRSnExO9dQBN22
/RnqsV/SBqU56qK4CjMqclpSXog0d6sLWcrt+u3m/ZA9gFVp3nWbJOnSr08+mBtuRQtLCqLDCvCC
EzIUEszYTOvYMaJswSk56yZkN2mtUefnMvTIyyRYiJbeRFLE2wTY7LVFUovg38FhkZfk0sDYi6VD
vCv+sKSWEcjtcPJCld7l1awie9IJCs1nsnwKu3bU6q/juBtZacgh8MiRlxrKCIb4D+8B20zm50wD
kSUfgxUjPcQRj8zEyuVV9soYmtX1BtawwA1AXAmxzE70t6KOx+OcBA/++7oRRBB6vETnuaz9qpOh
MwkWD7QJZAsTIwiELTg4bBo4FUnjaocQvgWkBKLPkzwp29+iDZc9TDmTV19wO6tWygWmVWxMATXg
m7425qt95akdnGr3RJ+RlXvBRe2axoRaTBM0li2Qife1wTVzmAcuUlXOJeANIdBWBtUqRGcV1CIm
8DB8YQVthtiDzD2xaU73m/0ZuZtRx9IIrpadeND3Ef9oao4fE7rGA4i3NsEvh5JuhIIvhZLRL2OH
EpIwKROcyFRN+PARelPRPY3e+TmbCpgzzm5LsCzdIuOx6mN9ZBlgvwzJlVlOHGOvsNxGy9ZW6pEx
smB8e+5HKC44gPpY9cKzC5N2iiFiKmg/ZYqdReajsQZHb9S3qSacc6Winu8RT1u8JjU/C9QYhN9W
yHxcOYYg5b8L3Df3gBZZLkB1gbbIhUbFygXEXWS4GvuDNBBUJNWK0zCOUONQdjxnDBRLifMI93st
ChSy9WSXUNntYOQFGeBeqKyvZxORCweHboX/+Zl7MUMEM/JtIOAdRws4Y8mkxoz11m7Wku3DZLa0
rrZzv38rfDmiiEd2BI5p8E8qVSxPJnzkx0MST5Aj9ON8cs6hJFJu+9mrN5J0mYV3wMurmgNS6A9P
6tvvrySwYL6qXfGJWwdYheGAl50o3Ij1AA3KypwJR6U+LNzq5+10lccfBiSKoGRAdXB7OOwZUk2J
sxPJpcO62rLGwoC/X33ngR8s+4tMoabksCoqKGXyLZe3WTSJeXIk8vsfKK7OMJa+tQLJ8uDQTjox
rYnkgz+24UH/990KC4fMZHpQ0+ppUob8j0cKy4W2bKGu/CCKp16kd2JXdAbCQdFW5mgWEPjB5MIf
v9AMa+ZImzHM5JvKu7g8Cw6FbhqmUs0JV8c+rDNOZaZPhVv1wBficHyCuaHZsXgN88wtAkhLXx/6
SGLqVb+8SNxrHCvzwhz8jEDjUAFTBbeHpoj7I4XhvDzPxQTgxaqMLQi246szRjqKhUUhbgSwRQka
7EgJcFZJXJfhiJnZ9uGJISgJyFunF4WneibSylMOb2S+r5kQLgOh8KvnpiO5aPywYQ6qhBuvxeO0
CsB6mTbLbxc8XcqPe2lfC8GtqpWyO95llxcAKWTATAg4z7kkW2Y3qhWHJQ04dTHoN9mdeAlyaSBe
q+5q8rCMdNfx5vOhG6fU5mMiLRGbjxrjFxET0TmRXkxzHKM6PQnH1h6NnG3AuMGs2dHuri6yrcoJ
3OSfxS8ShLqmgqkmXkk7VPSPUQp7DS4iomt9XZXKgTQy98oHfVY+uMnai/CdhBGOoTYqNPQ+Ua8O
hejAU4YSLQ7SljRh3RKE/TUDLqNL/ie3ncb/G8jssKvL/yxppgB9mGXyE/kQUc5Ily2enQ9+j5aa
KqxukIq42xBLIdDUoCsSk+ML7exlJ/rjQlvF5Gw8VQRNHEmQ2GqUiy+cWRFLJnQelJpeKwu9CnEl
M4ObN+IIDFYSSu9J7x8qzqAdP0UIlsR3pk8Fp7jVbw7GyaGZ2X0a8suviDiWTkaGjDi2uJNnC1Rv
ryjkt/dIq2Y20upL1I312JDGwqG8bdSR205QJ9d8jSlblZOL1kbejO4FrJDilQzTtF+1yQsJa+Zd
0PrDIbegfQDwWN0hB70UnG6SPVcEYHIAAFViNRud271h5aL9RLhwQr0FLXeCiBD6MoAVRlbNI+o/
hIZG9/o6KTSBjUrCbbitlYNAAyWzhdP3XI5v/dPEpVdPumfwlMS28wy+v6oFASGFurwSJ3YNuG8D
WZm+kJhLxoH1S6w1jQCjC3E5OiZdHC6ACt+CU8rKydWspxzcDXEkrlbPKw8cGSIMEP1pJyoPzndU
o9ekXuJG3HiKHXcBrbxocT/AzqjhR26eR/gmXeRBbv8fxz80fIjHtkV7gb+yIYS6abihISq1d7ks
UDIwLJN1HuJ4jJIR0ajoCc9L/CmSLmnGpQs0pA8j9jiPoQhKqkUJa030LbXvAA4kCHFYG0lCXSqh
1jJHAAAh12kcoNa1Irz3/2mSiMJuvqAh0hduROh8AvIDveF8WZ8RlPTbUilr34IdvnZh7dNdwP/d
4z9AtP5zD0Ioj+cIsCKVuxNyNJfCnBmXD/Z2aTOoJlcLHOabcVdmSyrBgmzWkH6GC0AjfN6MR2w2
kWRM4xHbfr3a7FgVZEKy/B0j/8476DoMaYQhT43Mef8qkXWi78pmrfAIPn8wu8RUJTl3CuZRvNgJ
93x3GMigiExP9LSTxvBls43HGlTuieAcytc8QpXjmIPyToEqYvZsTujor6bxlz+bODL6SFLm8USw
Z2sbcPTkB9FlbLbiqZFPjNRlShgxUS36SqHYY5tiEuCZd7YaPIaAKC+Ip3Ell9QKv7HVNOxquiJ3
LjY40vZJkLcLMIFm3RCmgR74eN+cpHj9Hp7/IxPXnmnYYzri0yzYQJ5xEEYiqxX6eByupZCIivZw
nlmpbzT0fugvqbX3jYffrTZjU+Jrwnb1e670JeQ7xsiH5dHj94oIUrFANdbDbcEz/bQHCNwV6HRQ
cRbN2ZfBZCIZWiKiVo4VPlT1XWhPJe7H3rfcToWgrOEokYrcITSKKTpLh/nYYiwrm5WmD7r1qwoo
qORQNMAqT+BEKbQSta8/iFIs2ZzzSeIt7ZiFAYQKmF54uDFf0PPJdvCBHF3AqOfo0IpoDT6u3YyE
NiY2iV5BtJJVlzqK8ynDiJmQPVaGi17DEVr1U2v+ecikfbS1VudrhngrWRTE1VjznOw8I0bvfrYN
6YcD9ORwwzfJ6163at/kzHwfLwa0ThEEW1ZIFT0+jVPpoYSZhSkVg/U8Qkus1Ij+ubJUbglXCpX3
2ZV6LMrZHcAT78oseQrVDdc0PYfymXi6j6TZ88oLR7DGBUfbAlh0bXEgukZoT24xNnC+mH8toTj0
uelYr6Qg6KoCKqmTjQPyOQ/hs56q9nB+3TDYAevU5ELK1BklBARqNqJPO7L2aAEro2QRBrEi/xsD
vJcdEP5uHRzwbCojl8R8VlmWiTtMZnd648VKsKvqVJGuWOub9yHTUe4cA/pc4TWmbOS7UoQjSMqA
U1gg453XF5k2rYRm0QktwxKvgnx3tfsNGnryv3oMDCK93QV2bdzuvA+kaJ7jY/D9jI0yAo/8yLpP
GoYdsQSGD7RGqy1J3jgMKtjoa8wxVo9xmIrd9QqMqjDJNGEydfDXc+ePrPJndB4yiyxNZ+86tp+O
hIUUUq82+2v+l4d47jDy0VmKyPJQtFSXiEZj3TCYBj0twY0eEqzkG5TneeAv621iTVii0vs4cH4h
yB9xqCrFD0txkW0LZI0AXtofuU6wt/rhHkbCtWKqtp9Bd9d0i1X1WpoD7r8C5hLy+tX93+GizePF
j/m2Y8kQ7VORX3uLVX3tHCDC98T7r0FLKavHlLFl7jQOulnamDMGMIv0umlBTEpv/PYElGvcIDvh
juktGCvj5USoSUJWMQZiro4mbWbLXMdugwAHLCBlQbNvbstvhNM/E21GLfxPXMSJSbwCYZjKe1p2
YwUIbnHue0gPK4W5L470q+GRvY60e9xR1gkD+oQulQKBzjxNxOZSCQE0I/zuunatLLAbzt+5M9JR
cDNMmvXA+6fcWGJ+ZtIrL6cyZwCoVsKmi9dU5nKZu89CdPGlwt9QtGDpoB3r+KGCinLaCfmlirFf
NBEA1fiiUHZYUCcJH7fBs3LmzheO3Z1ylSkHKoe13NJmjFFGaqSU4LJIdh3TlPMs6/jBoU+i6bHh
ZbjlwNM4/sFsaUBUwwGzJE0+lHFsbFoj/5q34/GgvHpzeGaZKScXJxMA8+w0kbOrM+UAIhxNK8cv
vD4R2GpillBCJPduqTr3hNCOrCv6HKj26ey9d9h8xhIpHO0H5yjOSiR2f2OxPvd5thQ20IdC76Eg
DbhaBiEm0xn+5P5A4lEPvX9lwPgjjW5sGD2w4Sz0teOMhsySvosEkUAYc0EqBkN+pgYpJjdzUbZV
VUSFOMk+f0XhXvL/Sp+dNW53l6rjTukv+D/62FqNCnf6Xh3MOssfAPmvRdetCEQcLitOverbcmBp
sW3+LY/SgFfX+Bu1u4BzPRDM87U8ahIGSA2+uHI3fNgf3+B/WZ9BDtiZK8MKx/VFJVUORKjwZi7S
5kfe3ehN00NgzCynaSDeoPW+q2Qpzl14NR1yQkqAtq03SopSMSW8uTVJYmV9fhWcvpCbyvJOUNje
W+yWeqNdXIWhQMsyO/Tyhz2vBmCCR8NT3u7bxqfK9wh3H0yHal0r8Ff8kqOkBXoi27Hl9kMcVd/O
dG00Tmw8AcVTGi6NVTPHZSbeFSvRhD2qU8S5YL717RFkxMZu511kc2bCQQz9ZsYNRaekUNRV4uZs
k2tajr9BAPNK9K6rhoXIManuhGopmb5mS/S+QKrXUeYcNZyqnLoCu7sM9lxFpLA/o8R4RkdIoVIb
mU1pWOq1e3SiH+hD1c3GpMOwPGD00ZMeJmKSHYTM6BzYmUxst49JKHyAT/ZxED5Mj3/FI5HV/ipy
O1sHYcra1ShrT0p9vV7DSEsm/3FItF4unpI8RsMEY++09XaqI5GyVEhDtGKupAeY10w4n2iqLi2l
10Y3sYfj1rkXBAxt10z8gqCAqUjVnIDIWp/157nF+44fLhPInc+xPLFKrT3tnCNHazifJvxMLyzj
3T7Y0RgizcuSjTDH1GKxC0KFZ88MEwZll/+Zbo4DAI5DPREBfHGDk4zPReQTVm4Gb0B3x62DidX+
rprGyVA5qC1Mhi/ngLcvKulsRngZE4PnysILbfJ+x28OpLbDgvCWnlw6o+1yGd5UJ34+Hhy+4K+N
/gzf7GaOOVvrdvBb3Rqvy2JbFFSSfE+p7Yxfg2FrnxGE7cqPNBv8fZKq5YxosbhshNqK779dS58B
zwUW7wDDTeGQM4SNkDyp25OBwUW/La+7fP8+PHTOUf81jUJrNEwhLeR6jmAScMyZsDKqNhhzKhFP
fr8tuzXJHJml6YOD7hjOVxKibngjSalvJ4b6nibTwNn0jP1ZkvzH0DcUfpIIl+4f3rCIQuhcS6Mn
CePHJvrnTwD3SL9y2uoWdLxBzMVPhgtJ+wGdfOoH+S6e55Kg25nzr+G2glHjt6KP/OMOQtK1/4t3
65GIb+crYdSf4bWAykqmO3ipk8cWJrpopG4WqIX+Ch0Fzn+p0RdWVJ2JwMmHAplG+aC7XBEQJrtl
c8rlz0YBu8lSK14vEfgZOCOL/HeF5dXxmc32XINKUqdhfCovPZDEyx5+OLqN91GIJad584C9Y6U2
6IVQ3wl2+3fhOI3plYvCzDNveF8WngCOMlQkub0hIaa7Q0aSL6fch8MWe0sTdUkgMVkad6mp3DxZ
vNAAicz6Yhqfgsn5XYvnLeUk78/8qcXTh5WiKxKZUrqmo6T/D5ZtL5K4i+aWNvV7cmxFBt3pT4FA
cPC7y8jtGiYrJZQK9BA2MeNZa7T55HPW8mzFz7sBmamZ1NU/9RbC22rDVDQtvjjw11lZWlu2AXIt
r38Xkq4Te633DmLrGRJ2qKdsufqeudBNXcQoQMqhtwZMwj4ILTKXb7f7xkY9JI9SlBq6+d8+nYnl
btI7dYX1RxW840yMtGP+M1aT+I6sKQI/saRpdqHmti74Hzks5FCCPwul9LeGl70mCY2LmzDPRS/V
4/9uSiN5CctHhs2TFVa9JtKoqrBh48xHrAhMFg4XUFKfzLrpmMuWJ0XCFJ+N1iGzVUR0dljAVrJ7
n1GPxTh8JoPZ28RX9Oq40+IPJc3S5aJRK1djevNlMzDK4kWj6e1iOaPCvq4g3Gdwu2EG49OqJDfh
iMbCpu6vr6czmh9AERFaZ9oX9l4mfXsk7kUaNyvi9cLqAG2ziF60EMC8dsMrWS3fbKcC7SeMRVMC
B2dmoIuAWpoPmv/D/ztkrO1mUcjBU7JnySqmnS+yb1NaYdezK5xpJOm7KOpaWMwheoABL7+idUyM
igLtMSXU6HjY5cNJL5cJwRVD3eCGss0hFx3thFv0lVFacONYtw8k79Sz8DAJYFsAXVOiFDg6m9aP
zKePE06dlTuRXku1ui3II9pSxky7ipRyGu9jEy2tKwgYTFFZSgaYh17IUD19Et/RyFEUDJ7Ay6re
2S5VqPRP9WCiYSuYK5vgZwo5gUqcIGASnU/tEG2LNHCKcNdh/qU3+0+Xis1nwKIh0PBVOymIW0Js
HJMumycSCI/CKytTiFyoEJkEy9YoKkhmbw18xaCVD1gahqqsAk9asNhK6PAGlJr0oeJYkPIsfOd/
WwPRpWyKVv6z7ZzGyW3tWRdgTV8aW7KzoAn21YUCBj9DQCybDDDPetud5RRdyuDJJXwqXDYMvtpv
xvCfOFGDNubg72y0y1FYYZ3bhqde6T2GmWrqR7C2TxywA0D013u4ClaOUyxye61ejjauWdF1UJRQ
6hyF82HGww3+W1+ZVjObltPbNMZVi/TyTOFY8Ii+in3X2UMsNwGavLio9YxUg/YOko1JlxmgylHj
yHQpoVG6IdfCzFOMv5rwLiNne3IfIUUrxycysKHP1807D8tXNHyalJsMRvyNUfoIPtKaG9kqVkJW
kzBt338UBtj82Biek2AB4rdn8XU8pIEJZblDP1cPPOA7ABU4jzuzRBODppKB6jxY02ONJxONf0A7
7qD7RZ4OFHEj2x3dy2EXlN4nedNzRf+tLFcLx3NucdCDNDJm7ETqbkChBKQfBNELn8hNmFshI1Gr
dQWPQ0Czi+1LZy5RG4rz+mXcYZDf8iA5+hwSJFRKbuP+fPGIEfBSn+A+RGINsz5gnW21ohyOSFLA
1O24jGrGpRNPYC3uYPtUKCrrnKtNjkjGvYNb6j7usIZSywc/LDtZ3zpmGe4Mg03uCMwtXqkwPSK/
wqaMnK16U54wSYqYfgnCDNUN4UasCFU/Engurjh3+oIBNxaF93lZhA5eWmlBEQbGX5NEr0we7u/T
m4mVzbQ8a9INSfqsKl8ycYea7CM2XJmB3AS35GjcJdRcTdB5eEm1KC2Fqo37XA7QURt7uAcH7nRx
wlwcTKuYji0eY9yV/Eegbg8LeUd0C5m0kX2urNTvrasqHEX+eAp2S/IY9PGWg8YaaTETn+Dfdtrq
TI2a5GlhDYgfHKxD2UJ9CF8HLu9Ppi0GZQ2bm3Tj00ryEZqbz/yFqdv6aWldrYBE2NWlh8HMX4WT
cXnn/JwXep+qcFG4bVj8UFgwyEwNZ3TcDAnzZNrGt1tS0E+82SSYoguFgm5XPBvn5XXBquOIfcSW
TdY7x0WfJ0y+R4aMuqxXOmbGlPXifZYV6014WU3CWEjrrku2Huq9KemUGe+0jlzq8kVGYrzRsNKE
1T4y414gMQuT3wXIwtkWttUdf1yBNu3zsAcdv+48768SdKHGOcEgQic0fmQ3MZfWSt66kQmDzc2L
Wf8bgPHdBM2Z0FhfnshxWNKwIufYA3LCc9UCDeeGJeUwiLr0JxW3qjRa3RfVyOxy8droJSehuj4t
4jYqGl3DIzr6mX1M+aFEjvGVkEbCVi2Yb0Nauc6HPhLxOJTHmZHmRFNuF2GL5mQCVJAIYZCSPAFE
IjrW5VrEd6YvLyE/TbN7TQvI2WkilD5ixo590OdBY3OOUwdak2/NFiF+Y+mayxJlT+VP/VAmj2so
nTu9IZm7JTZXP8vK28KQzTGOqNd0lmz3+l4r89jl/n6Qql+smFda6qzhw3l0D79WW5LblE8M+XHA
WoQaPigpr9TQ5hsG3RkpmjbAcC+4U6GWr9cXbhkElAdb+IVaKUZwvFeStc2Fd399LDTQHfly7mwj
+t2s+d8LgRxL5emrcuikAavl6YEh13xTCUqMpp4iokKguBPNenw5a+JnD/X3ux6kB+UOhALxo1v1
DbJHJmi+Xi9CNNrHW9/twhyCsgd8lP3Z51zqLBzfQXko1rgQFutbfN9/Qy/eeaT61ewfdMwkDiKI
FpwIua7iACD8oIHwbc5f8No/DJWuYenJ8/+ZovuCe4NEOHpVOszp3L9ctubm9W0E/dBnQ9yF7UEL
pSz9GsWPxZCGtHKhqOURz8zVVKEz1OE3xX5OcTqYnRfXoQWRo0k79fc/Cb61wroZd3Bm/NQ8K09Y
q2cuQyKcv3QOp8opSHRkdcAlQpJxTiwnjIc8x5lowAuH1j41czuKQ+9qwpYSw8bn1HCjcGIMOSPa
rAtfTQPSc3kviAzk1CX7/JmfC+pCc3s6zx1spqKGD3YqR6nIfdQzZvw8YSsKe8jCYnPhH/NkaZRz
WbxY9mXeo0aJpA0DgSQJ5bkaEQJvhczGISY84IerFi/6ruST1JLzbNh5fdlb6OTNYO9uy+pSVQFW
c3Pu1nWiqQJ9dyjm95RbQkioso66M5jj+OAfECY9WsrXvJnxcuzK8EmxyCUbsS3iT3mJpzqNPCLT
a/LbmRRj20ClrISvrqR6Z9GIAvadV8ToLMKgxQ8eECvEST4QuAOwnotkB+C0h5Jfm3lu2AwPJfql
dkhCazrvcCDbCGGAURFteMBMCIwl6mjkgiOBAaX0NGryG+YNQN6Pcdx4McH509cRxplrep6/opZR
bM+HazJoz0Xi7p0WOfLPpzvqFDJ6u6YG3Ol3Sp+VjTUZW1QdYfmCbWe7xAH1eIHgyWXUQCsWGlA4
SnwMwLtbRQg7Z55+h0mxRX+MCtTQ8qVC+yj+wpy1Yuz0SLe7elaHgHEcXRmXgdr/3mTfIMAla6qG
eEwDFrhiQukVSz6uWIi72bcP06YdGJuR7xKjCFC/xmJl59EFXKuXGOTjJsu70Fj9R607HgcArj3p
++HanJEiXiSnNzG0jx8Gq7eBHttmWhOb1X9JdKRYjKHRxMrHWoAvXmi8OyeTnLFK814IVSMs8IIf
+pbTfpitSI+Z0Tsmq97f1B6eZwjjVMTY8KAmjzIEvUj7ABWjj7kErqLLhdZacdSh/R4QWSpt3xf2
hiUYeD0MCzAQSjCpYs4Lj6rrVBGs7NBp0rqXzLWXZ8w1RO0IJLpgD+H15qHZsz9ZI2B3eaihcuiU
OQ41q8waO2w1G1KryFuBrPZbuPtGIahuf+pgEHvQKUdfJt9LEoEZ3S9IkYtg3p19STm3iejGpOq8
DuFyyOdG9MsEV/reIsWzY6/kzZbpVq8k/C41y9DrtLnNVYYTwbeTWWcms2JyzIyS8/VNocANAPm7
ooJHNK9eDtkeJnAS9AIAlahN+JRNUiZLOecRLrbwPTfeyvkDFCeBVfek8BRpnDSbBacCRqk0dKun
4WevOuswad2REi+X0Nymbtyrt0D+qnpXBxhbWIseKFJqhhbpxl5H7cguDmTlg3AsZ99gaBnwp267
/EcT7czqxTsc3ZgITG9yluWHYwiN9Itr5laEGRAJj3a5xs7SI37eZpBtGWcW6YNh4MfyKsTbcKZI
g9YmsiaI0ssxRzXBsKpOgG3Uj5lsrPYtOu7dI9s3/+Tlw38l/W5VHValj47f6y0mma+dg0qjRDhC
w1k5hXUOawnmX9F1bWRRckrB9SSOE/Dz7nZrgAubpNwiZ2pYvlwtAxpknhPiJ6h4Stxq+aOhYe5S
XhcrUiCc/ls2aWAsKyc8wV9EZLyn0NOzAaOurpN3EyaWzWRgmi5kADqbJOBb+Ui9lWOd7T3LqO7F
pfEAiFY1F0DptBPCx0TtYrocaWjUlWKNqrOWVcL/dEhqvVRbfhBhpfCoKS/wSuPRFc61Me/985Sa
qOoVMAcolVDJMVfJnr3gX9uzRrlRftB8CWj8XD5Vk/Y/dpTccq4iHtYEGXu5za9cW3pfOMEPoB+L
EIghbU4UuBTUjfJvhkOspkJre+simnjWsO+f3JrCfuioGee/008/RdbJzs/SMbtJy8YelKZb8feT
Ov1wcjeaobPZk3NrQgYTx7kTJceNoaTNIKZatD0fwxfvwGwuevnqnHjziOW5ct8ETtUfjlvD4uC4
iEOMNQBa1I6aHxc/sd6HVRhNKBlKQTXUal67UsgDWOG3vCaSdNR695mX6yr+FN4nBfwNQYCIQZrH
dx0Is6Hkv90fhdU2cNvStl94nJwsl2kpH9FWjbCPOYAFzmzgKiDtvXWjTpAgDu1zxGcd1ENFXkev
yjIIYH5ttfSf3eBRjBYrCBUtqsdxyQqnHK0G5Bs8LB5zmIkEkaHKB2ZvyNvu2gdN9v9vWv7lhN07
EGacoe7tBSk5TsyDGr8hhRn90nYQ/qIFGXduY1FBN3EUy/C48BhTl3C7KxCa5MHbatBsDpNe/vdo
sR53EAkg4msxz4KiX4RM/hGaMcxQ9HKaUzBoEjC1hlr4NnbqLRGVDVPjjVZv7GMRpRvQkBU2qObC
tQekJuMxhKtIOZG8u1aeXYy918onKuJObjvtoCRQEHjSaykkoKFJPG9+zBSw5nBzxIqMd0f3mPFZ
vm+inSHQkk4KLshwBcw7N1ZxcrmqwzE7RZoa+2rNzn3EwO/e4Q/pP8f782epE5RafgfyEp/FyVJ3
UhtK3OGEoDLk+k46yDCPjaiyJJfSRbeh0usWT+XycP+dKS0o+gSjV1OOjLqPKo6JExRD4wpwwtr3
FGPJDLHxz6kzDBQ4h7a7XJVbbW2CD4WaIm4ujvgWLkNHZmneGbrl58/SDCkXLoPoLjwQYpRVlzQ3
K1WSiyioybzErdMuvB9vlpupPiyGzftOsuP0cdc08oEfLg+XGSu7MjHrp1IG9cBDS5g4OYpmktlO
qq3aQRL1j+1H1KNYxE1R1luJji6d8v58ifHgrcZs6ZmXnLXcLpKaVorH+G3KJLZffwu8lOLayhif
jWxcYDHRwvtvu86gm/bkv9/q+dB5AFWBZtXdgTNp4n/j34cO2VQTnMBtTUEoM7ZGpa09M/2W77AM
YC/NjGYZ0DC94f6T9idHhXFC/mQgqvGsF5yUqRveFs6wYg+pMULkjYlurCfmfrdUNuGzm0FbmkhS
emi2UtuBU/zQKr64V0WNazsN5k/a8Xva33PozgI+QfB/NSc7qpNokGs0i7el05TV0uR4EA7WS/7t
CxC334v8Oo3+Yq6F915rblTZMhM7Mo1CG5Ov2B6HJDSV8+3goRLUaN4JQA388l7o+xodGfbbjMmt
wLtgYv8ggjp/irwpRQdjByeSM6LWbo2Mzz01clHiD69lYAXhp4rQhIiAeOpNWsC8voMzfLEE1ib0
khBbKaroxHCc2+/4lXJ36mOdbQqdZDLSuS16xbciAaLoqIzOT3qNkKSg9gjXMoldMPxr1E/+oxAG
MwOZzSQm/FSPgaIZG7Gr3+30DPhNE0LoNZ5jFTsmeqoBCqwYOqskIKJjJiLX3otRzKxbrHEi5jdv
7ljZQ8B0egtlM96PPqOk/b4AbvSbm8yRQL+1yFfwIovZ0VA/TeIB+Zi9gRpFTCk6s8F69t3yl8de
IydJ2sVq1Nr1Ioac1tAQqkIpgaYeTEeTJdS5ceYxq4H2efWS5a9Qviu1GgH4swyTrJ62WBsjJ2fY
BIkl7AW9N6OeeHYppeKziLtDVZbxKKjZm8RaBrlV7aRIRqdUoGGCYZQoCCPVuLLrLLG0tnbVXpnk
s3nGgSEL1x0SHdTM9lwwxpsC8WtMZNvF8w0+68ZQHaQc0n/RuqppDj7Zy0uHUKx9YeNTQ6ROs63Z
yF5nINMiJrjVc1GYh9jEaXEu8/ZoLZWZtE6sU8ZgynaL57sJxUxQosjctKwnO7qxlkWV6xnKgddf
bZTUl7XtZ/Tr6xCJgzs7TheBgy9F4+4zF0AE6j6DMDr+q+MJuy7RuVdzq+Jz4y2bgPmzg0tc2JDC
M+PbQPqDbYrlhDTo/LGP6kk3dtcAzCWvCBAno/n6xAsToCn4e0sp3nNy3DYgTDgJ2yOm5EWf8AUQ
erQ8VfJvD+xgqkMr/NkOo+PbPWQyEKjXVbFoi+iundkFqxCVa5xB8NG+ufYxWL1hy8Fv/Nx8N2kS
AMVKPg8f5pgFW4s84bF5Eefxb2ayjr9k/QN80+X4Y31ZrYnYI537sbnUAfmrkVJF2uOKroykNePd
Q3KeOJGzQHmPEfVfrVE8rSZa/49YM/Ki6WfaRZ1fA4DX56xg4YUTrOc1733U2gYKcAsVxNKd8Oxh
3YBXwkZUvVgQkvY/wyRArL90TdiEKo60l9mMC3iy95E9btG3irc8ShtDx4JfmWnuMHGEltakWIYC
8ito4w8ObVjBZJlLxrD1GUt2VD7OPuDUdXZ3cwdGU8WpIu1DVQ+lYkWPg69qMwd32kVeUrlckDca
gN1P+kpuP9gq1ieI3jwRS7pI6YGoMWo4RPPoVY/DhT2ozoq+z37V4PU/hOspEQrovgoPc71qiYU0
fl7p6NoQWAiRAfKiCvTKc6E4hcucefAUhmbPLNRhLpkWPQkKB3bPsz+aaJkpxEByiMjJ1Fy5TNj/
RDe1hJ4tYBvwtLH2X6lCQStHQGQWtTIwHkoRXvWrzm9tWKol+w3BV2jZm70aynRxTYRIhARFb7wC
7rJfxLlydWfzrY3NKEKUOMTQOk/7LDcmp4hgKoFbX0T8mJ9jaVFf/qqOwcD9Pit11jiX7viMh9A3
3fLIj0JLIvqNX1pjoMsZdTcfkwMrWDHceuYA7XIlV1Nd2YqIwpff03N8kMqxV/7A3ysWRlt9L6Zs
rZXp0mDiy9ElSx8O7VP3CmHE9J2rJfwydSrTcu+/5j3hpgpDYikhbbxeNWnbMZ7veo/1XukbXZav
W3VTCERrCEdOWSGGXKXmg+Jf5BKps3FCDkASZ86Kt9xVNj8z/gxYCnzwOySuTar8E9igCK9A+Zvq
FT30QsdUWyDq202qS74KIqGIXkxMMnb+6NDU+84dX86Vtho9fhc0nJgdQcGxM51fqQ6G4Qy6PCTj
ExIu6HW0K8ifDYwUgDE0QNrvk/4BmOZv0fFTi27so8IwuR9IHK9Z8KCKXDEGyMZnjWLzI3NxvlrV
O05iMyY1fKI/Z15kOMMQ7N2/P5mVpKq75pMWjl0zz24HrHDddqCPxgdx6iFl8f+P01iOWLNENiyk
J5cFTC/Otj2AuVQil0vkiL2uiAbnxX4VA5MKb5dWcm9I0PaSwAuNl2eAAPyy8EH4PipuO28QNNEn
fjhzbS05c3ahjPDvnKcgglZzHCfTGQU25QtegIahdtEgs/Mseze1OLnwIGz5/Qo7G+1Tk+V2gKOa
kaexnuy45mkMBz9cQE3XaV8YQ3IsLtelK3sXhsdRiRZfZjNy1XJNPSkW92r6TapRWQEMuFy8wNrx
ZTXR95Sz7jA6yZvIyJrA8mRQCnX3z5bt8tATBfVZzf+WBp1Knv7cdbq999tQ5Fj4fkEeoUKcwffp
WeHQ0F6AO2GNJue4uZTKg9LYQjhbOGwsOYkhRyc0RbGEvzUO/pyvyqSH3PETgOSko6bsyOZTJnpI
Xwe9Gv1S2+u59UFhvzg/t7L9PtQ4W9/RtOOZFgA/F71rciGeB3a547claZ+2yZUoAwhEITL4KfhK
nvVhb7JMVJR1Kd2yiTazuBzP+09UgtnsG5rwgygABVY2VE9nYmUFpuvDWsovG7hR6lSN/4YVthWc
65T8H9dGG6D4cdH1Vb1jzjsSbNTnLsbBRtpnh8MneqoO57q+U4pS/Qj2OQWG6e9wy6IWsdypyG6A
Mdx2s3za+48O3XChhoRANMfa6qsrpULpOM06WwCBZwmgX57k7+BFNPJE+88TMmJ906FnNb2lLeWM
ysilfh12yJynLhLsRKLq7+rxe2t5ejMDjI/CUX2FLPtkdHeFrWUHEvXgrUfaVn4EdHxGnm6f/FDW
zGtEVndA6jhOrEjiYtAU7Vs8gYTmlRJLSqX/c761PbGEGlAifBMLADeD2z67ds6Myy/119O1zYQ0
gVmr0vC24WHqKES8F41ecEZVKybDBuPLNHpZ6oqsc2cNt3WI5qmgJLs3m4/gZNcTvocE1I83VR/y
+AalQk36+71R8gh/qCVCzAXH4FtOLhaFIr70ku/VmGp1gtWD9d0szYwlXtoT/EQvR9TGunjRnfIs
5P2MDecBx+Ym/sh4/K3gwueZlP6DmW2t9z0ihp1gkD2p+yQjihDj+jDhSEfUD5D5chf/Nb1T1W83
T23zzuiK864+X9+QBXdCGxT7M0pxxuSw9kVbYChxWfX56SlaBEFi1pMLspp7MZh6lXdhnI27I4Bl
aAw7obYaT0KQ891fnFIj1gIAh6ixAY61/4oeQ6RssrynkjdlTuohF3jkBVkKWGEG+K3n7fUA6U4l
JbCyj0ggZHetUnIaUsSQ2hcuF/AMeFWR/XmZ7+KsEtBuEbEGc9cyxk7jlqV+RHvS02ZBYpFuTKjC
vK4Q6Tn/bQvv2Y6mHnTYSKVDmEb0NxDxEy569b6CZyoMiNLsC+mFlE8RlZmnefHj6lTvMCrNm2Kv
tKf3KfNoF7Mal/4HApBobFX8WQHccnx/ZCS/2kiYQ8CoT/+0Bzd+Fui3foS1BdG7dryEqqOp/F50
1JHbFMF7fahzsQEEY+XLx4/CvMilaXTXWnVGPbaoWp8vqoVeLVgVbhY/vYSqlhdqKhNu8UmANL1o
LRqGrqiK4y5KJ/y3UKJitJGkCv9dItK0HwUTmcy3r8PS/1c7RQxrqAqJ5jKtNGUVxsEDeuZD38oo
Sgeg2kcvF+8qXDG6i2GoJut15Y41rOQfYf19VS2sSrijKpvNByMSKrhW8/1/jWkHmAmNiXsVt+6Q
mOh6r31rzwO0NmXDdK8dSboRAAVuez5N+UHZiW28xhz/mIEDXA/McMSNXfSzf7sIo7Go1086nh+r
H8RWmwO7agZo9eoZIuhYSzG/86quLVzfGbpO3AX8EoUZcoqp6KRdKS2xLS8GgHIIqN9rhTtVf9Eb
MEzZJSuVQPnt+EqNU50avIIFRZgjrBmoINwF2HarAZ04wfFltLS2QhREPdf63sBG1Rj7pvB1dahf
EBw+rR36W6UneFij6M9dJxAv82ItAysTrGadtkhsGK/xKPx2dUdNS8cTXV6gxg0+7IFzrF2/BjXS
tl9AvN1lVGtoeXaK0HETVXe+0ybuE+tqLqTOgM3W2ioSjarX1eZ+BCPlQCcpObBfrvOWrlUWYkU0
Ve4Ys6Bld3/z7ZQMGeoFvbRL2+ZCB/h2oeC6UgihlSlBddN3bZGBNLMMCv5CsCMrAP81B2bbqGNT
QOaohZ57Ubp+ZmyMDMxKehmOigUGGuXxcTsZkQ3ZTOCXw8pkZAdtNFX0KEFNLEfqtYIBcq0M1ylp
UeS6AI/hrxnIeKf51yPvvJnCKIUoth+9hPhzC6bBQTsddgcCw/giIoxJcVhMeVJI1M71ifbU71g2
WbRBodpm7LrHO7TDV1S2xeoprkU1E/ab3ReS/UHIvq4CFP+zG3ZnISUCSVFya3d8Ar7FmFfvju/c
Z/Sy7zfroYDmFvwwrnAI2Jm6h2iLiNePW5B4FRR27GZe6GSvSwA7i+gMNYQc0wSo/be7+0P0HBAf
CLOzpJw2QLIo3ir3PnOtKICNZYbdB9hv8pqT4Jcc94xB4PrFsu/QnBFrKvo0cM/6C7Ng17aEeSvp
0ihYXXdDmaWcGK3QCE4LMZQ4iE4J7eW9GX2vKDpryO9yuw9HlfxkDSvJ30sxMhmib2L+jDLj8UdT
8BalhwEy7kAYJsb0fmmDNWixyMkDbyzf2/uRn8Vt+WPsilTvTNC3JgrJ5clYzWtWVkKTSmgALp1W
vBm5E03ZFuNpsbp4tPsbBNaEfFVbhihOT4dTj42EhNknKeWb4Te1goL+NSobV1EOU9soeJJWdVWB
7+E+0ORKXxPzLLIfQDps1JmBO4XTkGWSW24jzy2wXZBQNmPkD+Ux9Wp+08cBzH/nat4J6SWVRfh4
sljt4eg/TiKia8DyHCePlsCoBa2H5GAlf8mQnfx9XL1tNKtZl7IhZHPqh45ngmAxRzpA0HKriljT
dcltSFHKQLP8C0ITH4YYN/6HE7PglXEa+Bm+YStq3G+EEdh+mIXwujUUzIKL/W0q43dcBesSF8yN
7M3VKSlH439MtMmXmWFUw1bB9pVmOeK1ufCF+/W1gULk4zgoMvX2D9J7czkHw1QEWDjFzFfORov4
DP8nGsheIJu+84VZER1LJxudVZDzMQA9bzDx1ifZcsVGMPTPeflgpMX1yIW25tkJvw6yq07FXZP6
p+vUiG2twPBGxrtmMVseWCFlp7APLwPipRrFeXEDmi8NRAJn7tVz2l9HXYffBbA/mUiKBl4CALlL
3vfAbQ2KFVfckf65jtBaQvh+YT30xWfBTaZ7AiuRjk3nWnzgckd6xL5FHX4cflfuTESqlNdt7SZj
OVB70xl8JDiCNr7m5lAgsCqcs/N8jlf9PAW67oD/l+WWejO0vt7+Zewl6fBDAX8rn6MqBdkjch1C
LJCTCtq9cFfaZSIU04M8nu65BSoelPrE7P09I6BJ31GxdGkiuRcICpMxVpcNG6NffSgnQHvnLOZG
N+Gve9fbUV+M878KV9I3dABt58NzPF+KwoXuazbA21up7saUzUwG0/5ayZrFDMbbcDj6KmY/h9yt
JsSJtHDayPKmUZc4z4lpZ6vUNwAoakxJ53BgZuI54N90zIse/56MSc4tTS2fEBpP6z0WNqIwGDMq
rEQoNxatfc/awb6xtxzICmXo09JcXPuaVi2To+xVyVi00JQ/mlRgVZ6egwWbisnwNrETqRGuZ1co
ZaPbmkyFFBtE3nlB7ua3ow2bNl+1B319aTWVs+oIFrbGudjgRsC3/OLO2MXthiHF5g3dSmHoxkPm
uRrBCGY9ejCjhWqB7fDTblQLTfz4jsg1PPLi3EbOlDJaO9lkm8w9SaiDl+WjOSAuHgDpKyVKWvuQ
843dJid/7KkTrEIhMIpA7eKqyX3Fdjq9LSWY9jpQ0gkwSXeFo+wq+qvuDkvFaPjGb34bstq3W2Od
DpH40ER9dW0J5KMc8fCm5GRhB9xw6EcGjxwvbI+nWQzT2etoRmttVuEbq4E3+wSFAgzmdLUD7u20
EM7Wuc82QxLdILi6oNsEhp0FFBm/GjENebEP0IMEW5NTzw5WlKA9ueBXzQ1SbOKCYf/rke/3Y3Eb
tPumbZuD4SUXD+iINPSzJr/zIId+7NuIPWJkwjGvg0lkPn4XQ7DwQh3V1rLAbZHjYqNjPeLgVyo1
4MjVDFiDTtREUtCVcXJ+eibQkGDE+mxh0cs+Joapj7yS+Dov27z+mBLBeJTjY3ok8OlZ5GvmgkZi
q2ZmbLKKqJTpGfJuRawz9FpeNARjzCoAoInt7NF3hZaIE0x5upnt+hJ7vHyT1B0Y58QI73zsoYcT
DHrx7pWmVTrQGiB8Nissi1pk4KYZx8VoxZbOWhd0/aqLhSBAeED/os0JS6sEehY4R1InQmTZRQa6
1n0TNOatQTTsUG01uq6PvEu640tqGvfI/t45ltH61pqKGARnBLTLDSqPwAKGY3J11nfylt75FOPI
zgaECAuGhxfPb/DJcmF6G+tPdFavryqJcQ2V7X5dyjXozFow8ixSHh6v/QBNwJ7/H7yQuaVLr3WE
iJavNKrpKa7FWaC2NUgUKIOSZQMHy/dQJ5HZFGXB2FuN0985eeRd1sGfTSQbAMEtTb8SX96yB1c7
ho4g+npcakESrr0Edf5WR3r/YkPNF7Owq+O3+A1Rg1TWsYh6vDozZtBbquQ8LSwGWopATfYKaqB2
ylvVHKzVZxU28NqOfeuWnnFRjdSRd/5SOA99OHRQ/gMrQQVvPSc3hthJxvrwClYGbnkXUNgivefM
ruV6QBAE7cV8sNlKnkjkQcordABJlN12dkGB4wds8xvi8mBQdg+MnOBoaD85ffv43VTyD8mDPunq
zHWT5hmZxjzJl1ZdFVu6L6pTyG5QT8MkiGUhyOJAnFxf7MMl2b0FBOEKuFxcWD2Ar9FtIWxC1zaq
dT/MONkDTY6lNqiWxGyuo0j6Bwwp/RfTad7j0fzzFBvlUeDKgtQx9HVKGubbNH5YhtL4QWVJ1e3D
qtPzuizRoC2dHK+YniM9Mxpv38nnrAn6x0r6Gq7CWhXQvWckUEJFNXE6iOLA2jsYVY9iID7q4bV0
hwtDwJe1Xf2jO8B9QHLYyREn6fyHuuDYO4cqfEuKSj94clxuGI8XRAEHI3WdxjM4ayrSS3fHhdla
xnje3sUrSdEQTg0XtDWpPJ6LDxenmPmkLgEbfIc2382U2j9yeGRgfniMPlooZhzjLIuEg8wf5d8L
jsKXHKb40xmdFMv/l/fBAVGbYpAAUSVoc3dUveRkxTAJU8bkI5QKED/2Q3cfKd6f8Yk+L2L0pNlM
y5r8xmSKpsGvoipj5+6ktzRNRMcNWCRi8U8woH7PMIYWcL4bytgd8QZjKrd182KA72n5RSKGQRPP
WB24FhXAZK3hH+/9Nopwt3oqs4SLhJQfziFAEVm87q1WSOcpQg0q5I1SfDser1FYxeAvzxTkOIBN
GYqUtOZmeq5niMxYE3GlWaduFCrgZHnnqPFK21s/gVhmino4BmcvXviqa1ogCx6rev3cFSQexwcn
eUxo7b6q3YCLSjau8xFyck0EgYe2dTfOw2R+eCiLHYv1jYpa1jcmqyOQeDKaFBDKbUZhyRU6SLfM
QDj8B0E7qqYZK7TbJwRu/m9GzuSy2M/2wW2lxh2WhGNL19sr8xQqM+/KS3FxiQpKMXl60NV9vamF
qcjWaZN5doN0ZpoUk0RekwS4bNMb+Z3NXxDcoZh7uIzdmLifeETuZl12emek0iE8xRBrM2BBpp4e
KTkGtyuYB6KVE48TYqi3KnIjzKjm4gasVLzg28qs7ND4xYURKWIX/ORAnnqwnAnMdXwMptVSA6wy
rYreFTTEmQ9XSjPyRKDppOFm1Yms1ON5SJZMlfGymskMCG1XahOBMSGImT7PPyLsN/sUcYWU51FE
+/qtcnKT30Nx8ezQ6Yv4ua0v9Viskr3oBsUsZBhCjj+O9luPPNgIzW3on4NnJDMC9xC4DqtSQtjy
K8sjDGfAfn0mTpWidyI8ldqobKewKVXIcSTVvjVpkcLdC6aegTFRDYZ1rPgYS8+CE8eQULBTYs91
Bud1RcznOullCy/UfTnGpuEmvpDRh+mzcHvz6KaV9hI+bn+8hYDBFpldigCC5HPC8eFTZDdS8TV7
u3VzEspDry40WHEUKazjxm6tNcg6EQWy1dyKWbBnJMYPPYxYT4XBdsNGXvGyWapPOpVyLeCJ344T
pqGEbPsmNtCW2809N2G99wIUTO+qdI6FfdOBe7mCrX13VdGmyjRy0IcpvYYgOZ2uVQo5ukm/2WRq
3cdHNPYvFvQPOdML4bahv/P03ONhyJ0vMOLlMhjpYUlnwsLHbTuMWHt+g+HkAvFeM61nqPD9/8Fq
Ii/2h8j1OdDM1Eh62WFRXnImcCifUGSF4yJ5vz3Fm9T1R516dcAL35ghGBZvXT5gDA01BMfRp8s9
OILm/nDm+LFJ/RXDpscDekNJ30WYEHl7PBSITl3xVkjU++kene/DxiTniQU3GCRQCKbpRFU9lJlc
0aFZrj2B9tmO0n/v6NNKq7tK5YJTeewi+viMy3I5kI+lzIWDZtjES9KHye6YviqI9z3STqIZxnNp
hHA7xf64JUe631gHazz+G/vtKpU4ZJGSSuCEyCtS4eIdGoxateZ20KVkTa7owMUtZKlgiWtqsO5E
esm+R6k/1q0ZPipOsN1nlj4Mn3YOmmzdeGkrIV+YTmQZEGFqAN/IyEYL3LXIm1JHM+qkT6XF76O8
rr7sftRm3iaPK2eNLft9iwKNR6kJaxcaYKx5JE2yeMoVZB4QHEhNugiE8qbR/JN22UqD7ppswQg/
6aM5lLKnMzaDMrizq1fSwKcyxGG18TsgA2B7PZY7WCxVKL+2WbRaX7PFRlgO3AHZfXexAvLn34NE
VHof8SeFkztooZ7PesxJq5X+BpUN/UnMyVmYp+ZR8E439OQGg7MhL8gghnO6AQgonGX0dbjYD2xk
/gjDseiGKKVhx6ZLESdZd31U5xWSuQlKBzA1dPP8Bg9IpsFhQm2hqi1RASm3x+3mwE3Um6BDW6J1
8ZTP0/GnuzLBEGZGUTtKg12sNzw7bOorEmQVl41xKeSyq1aTpNeKm88oouuDe2dYRWqL7PI8/Qdh
ttq1kfidZ6ELjjL7yd7JLfxmozYOM6uA58aKjpueANn4hJZ6V2nVsQAAnYdUJmj8DTjYTom28IJk
ol8shz/Tx5a8GO0c/J6kSs5BdNcKHfgiRs5k/SoRNz4X8fQavFFm3XvQZE8ISEGD6IMdvsyh8QJ6
LG8ec45Lm2L2oq9H/rxONCk1LVTmwMD5+I/SEn4mQUQrVygznYJH3czTDVtSJIvkStEwM++K/Ur9
L0nRdE18ITE3Tq5HiDgdIXuih54vLrJC2Gg7eWazH5u9ybl4IzQiRmN3bP8bCeOq7Q8kIAvPHUXX
kCFzDMxyN3kqos8igqT4ZYqMij5k7hj0PIyE2xTr87GKFj74tSWxwiU9M6co2hiwmLR0hcSmKNzQ
c0zlL4o620IUkONi930VacocXkT2au/J7z/7OPKdn7Ury5zwgIfugy99RPg3jNjxXTQGYxvKizS8
bwR2eg4d4o7VoLvVffjRgobiT+wsZU5EX8cw+6qX8at+mJNBCTImgAip5b5hWSVp9o0BHyXrTAd3
35+3vLvLChV+cozAvK0XVbugdr6wSUr8No9/bEz8OWji7gxyVo22H2a9M+wGheyU3x0yNSdiuQ0n
4h9DykR8BI91OfnR9LI8Ry8akWcGOkpOl8lUCL88skMAMI9kx1a79BIIgPtyqWNc6Jxj0uITxMDY
c63xOOJG5WsoRoHj5LgSyqmlkbxO84L7mVVfi2ol2z6tp4o1UhXrqC+ebTKS5U/+atRyinuXLP4R
JQE62VGQ9sLuvet9NvsnmNQXVbc3bAhBc26DY4RBYEiR5RnOUUD7ZVfwPuhk3v2EaZUjnJFX3qvN
Rc99XqeqdVdfnCpymOfYa9TDYcIdghPOrOl837J6tuQ34wleilzsDz2iWI1MYc3IuKbs+yLMeJe2
kHhA25x8cXNCK8+VHoPc0zXPSqWhtU4HUmo8P/TqSmDY+zNzRGayiDVIn55MW9ET5HM6zkUsegeZ
61E5V2MSRn8wOmZSa//3XAcRBoQ9atW2mSynNK0JaWUuMwGhQxBFltBpFKXvgVwTGtKT1/25vY2T
Ef49bTHa5iK6oA8xKEVsa2Qnifm0GZPjksFrhVLBEjtL5xOkou3uyFbcPazWG2lumNnnQFlu0G0O
ni5coVHmp7AtV7gyfu7pMLrr2vPjadxXAtuTGm5bIRrMNY8g9MH3eO8Nz3bdFhQaeDCPuCN9wjsI
gDFy0P7TTJrIbiEQ2jW5U91QK9CgeAGH/YGgJyiIBeoHns8EgtmQKWyQdsqjdPIyK3fm+MJudRDL
QrLKvia2v8XT02pU1reBVmMOB5Splto2cQysXHM/Pu5GkPIg/s0fSk3lHEkHNqNNxj1rZM7kLqlt
6Mhmxl6YJCZyw189x3MB1AJ3sMlSb21Zjg8GP37GczNDEPpNaTemNKvbVQERg//H+VqpYCZtoEds
ZE6jDs6yCDIEc1H2zrAUaFhvhmmg8h5KF8SNy8dTCnK176TfSoRsCHcOxovlBqnEzIMvnpixL389
CJz3h1eLCBQ8ZGCtnX6BkxbIuWBxs8Qhza8ihcg7BkYw5BKte0O5TC3RcVb5aVDVWdaXt1Wax+Gl
PNNFOlV34/nUAAY6MtUyynyhIbLnpD4XAuu6lQqcgzYxez0GloVQxseCDGYlwNmwGLvML1dgAY86
BM2oHwnq66x+yIF8I6Hh+bXsiPupdPNvZD1Fkq9Ot798PoQ5C9Q0HwsnSAM4bSsoh18JC6ASuQup
/qdyhIzXT3rXPABnQ/Baen4kV0hBMf0f19j42NOxjKPZyyE9I8+2FDEh4e6F0FU+YBGxaoaAr5iL
qmAhBRnrJjGEpcxWxLGAOByqeo2u+X30Py/6hj5+XiEdAnim9mJo7SxWaOy64xDiN1TPn906xSg8
F5+wqmD+ObWW3hqdGvPxpUTWXtBipkkYlxEMDvvQLY3l8LlecHphIcmqi3jE8054oRpADaKiTJDF
iftxNMskU21YSXuy07McU09Yey9DkXwhSBFwQRic/1Q8L35DYNYsIcthRZUyOYHYT87PXjz2nPgN
LOkCwSOi7y37tbs7wtUh9IfPyS3YqaV64XzGjm7O/zidvS3gdURG0nRlmW4P3Gqn11WD0M9o0uPk
EcRWrL9YEDxd7BTCIZTpZxI8EB10ej+9G+/DnhiStmnO8eJdyytfNM/7e4dPaw9jcHCbtp3vTcFM
KNUCVtZj9/kFutmr8Dbqt/FS3Kon4L3BnnuHKm5xXbImM1wNOEAcnvEZOhILSKlxI88mQApT9Sxs
/4FUdkTAyMD9QJwjiEQMgskf8HSNNYpFY3Qgu44Y1IyTSzN5d+N0OaalpZTQegkMuMFMUCxOsAeJ
vubm53xGdCzTNg8xgWSqQTofHTa/bvOMjdPqmTuRzhm/9Hb0/aqCaCtHTy9g4MvILy4qNoGXfPQ0
WfQ4F4NKs6mOmoikyDV3WPE+R5OTVwkyD7WVTmOtny6RAovGl2wdr48vvl3RsXFa73HNVIorO+qx
uEO5pUtz6bWOWDfwy+2Vy9r3pOYdmDzC+Mn+GabdXV/L/fqbANba9GL8vOEGI/I2mkUSWJjYCyeE
s07cm+UmMPOCWtHX+MxYIkAPXwciZtEA8D8jWGOqCDR5dSp3RPDs6QNs11jPalHJuojPHR3DswIt
9g2gz7hKZ2DWGuARUrnPOLEEQe0YkIPbYZ9G2s0+OX323qYxD8s1se/TkE3DphTy1sMJZbrP82z7
FhWG9B6rjW+K/XoRqtvgfjlgfwYWMhPnp6ZekK8RL1acNWhnlXVL2p3B+XxK93H9p1W82AtIbnli
AGwbL7KpnoYW2EvJK0QM/u9tY/iFKyVK0VptwKxIHko2lvX7Wf7y1wbnX2Mc2ndv15EDLnrK4fjW
sXyjouGRLELm0mIF+Kagzls1268JNYYPugw1au1ouve2+0d0gRsOJhkKwqZF/Mq2oKkIZc0dskek
o2QRLt1r8Km6xpXTHi/zY0Fif5gvPNNw5iHEDfxG3ENgxr+V+kgEIRE4BYpl4Sknm3Ya8FiSXiGr
gY+wZm5mgDxUCdU2FEfopoBfAaBmvtK9/Ljz9OGkQWkFPbbKVXlQgvDt+VOBdfpr0AaeJjGP9RNH
fqHzA5VOpvOXRCsHjUddk4xkVMq5JwmCTr7ZWVSGC9PtfQSvXZN6pAJ/BLtGi4+XoOihrj1JaCfl
qwXh6UwPYBWQMnkFe+Y22HKIMUUjD2vI/Kp/Y6DtWkDEjlMUQxfudEApnM+p+u6aKnmoKweG7/N9
1oe3ZsBDN3CQrmWKpaqtfsewW9ePYLIR6h4K4M0PcHScqNnZaveUlfMuJYQy2XbIxKtRt6cWw9i8
uyE0JMz5gXYyr0rOZRsXFSomWG636GTCgJ/YT2/O0a0fRw4zl02WA+EpkW0XsiyGCSZvnT2k4WhZ
YPujtaiRpbFomd1+UsXx+FPpTGpuFW4NG8BowNTiEw81MrULbkQXWy18x1N9PqvyFU8Axp3WhjtD
P7dbdWlqCUHjWQ+/FolklTUk1Hmcu3VzTk7dXgHS7JxrsHnEG6gCQ09HIyDx0zbGH6xKOrr7b54j
7uVFbtuqUcOyC7m6Tw16jdrksF+XKigqPn01apAvdXWhgpNNjKtA7UHY+YKiIsHuW+V9WqvJaKh5
sINbufrMxcu7Ox8GtaqBWTy106ogHoykERF9Al5fiMelyywWcPt+NxoG2eUcLnbcKZ2+Pq3LwKfS
gMVmnG1znIKryPj3nZiNuwz9qHyxRTk/umVJCHcsGny6d9Y91JD5keysteUpDcjT0Own+4jWEcvw
4oHMHgWC1mRWNrbu8CEKAow8uKTKjKWx+DcogRoc0c0ja+9kWGqmimL6jlUW0hfxlgpF3AJLDfiq
B8QSOBxaS3XPgYlHobx4B4mL8Xy8kj8X2QqTGt/k06HNmjG3Z51IYn3hUQAryl0COEbNaHKXRbRd
xHFA+FNAMGkMRpCX5CNB3DNgRyypuJYq2fiyHRcqiGGaTVuAaGVIIX5Q+6i+ipSaZncIkKKQ3NrA
ov4SyadSBN9/rS31jYXmmUGR7DAAn5EEZcDWngQ2dFsUMRT+cRaHCykPHWscEwGZSBM/618ILO9J
g7MagNud0GQaSms6d5oEy01gLQpuL/F3DrnYEiLqZSK862W4tRO2GRF9o3aMck/1HRrXOkDnshqF
FCJAKzu1aFBVLRHlpf01VDjk9oV+bZqmhimMAbUtagKZjz2BzqpeZQ9ugxHpRQ87Fd5442X3G2NI
cdiHSQewnyZQIRUPVt6rX+ovNuJfnFcXkwW9C1fR4rWQty3uxyazKQyMSu7zt59MIYnrtIgCH2gn
qQQ7YnbgkyHjgaBfEnqqbj0maE6mTSyXDMZqa1ShEzzvTYkIqCsMuO6dAy2VQIw4dwes9TSVn8d1
sZ55Hrv5xiMEZzfgEeZGRltHC3ELH2Ia1dWucPK/Uy7DxEM3gxuRKl9n2FmWW+TWnL+NgtYdg1JF
ILH6tixZfQmmSy2x4LW4kzCvpj6KcIlm8L3G0dnkhJjzKwKxyo4huj9hGmq/lWuxs67et/+gHZs9
MoR4JxbJ9O303w31xECuG99lQOdG0ehzlTdgqZAuqC5oyr4B+ulIsSSeRwnDsJGglxfymvznmJz/
534uLoWxhswJnBaTe7Yn8leZbObujMSrxkZInKM0pXLmf4tzRoyw0jDFTUIthUejDWWo+QjLhruq
+utSbOXaMn8LgdRpk8aSjjlNZYfSOKYIMyZ3xq/TgWbZ/Vt/bOmYDgWIg+GGozwF97yyjp2usXpP
P09jirXxgP/rmIdvJBJFnXgyWs3biRn/z+vvOUPnTwWZhTBPhv9Cr3gcmSoH/F7ViOqw0wL/NHpW
u8OEqXrjahxT/RJgl/FfX4CyNeqCyTZAC5/per+QgRbY3OGIbnLTkTUFD0pWwvjjgBBuoLgw1VWD
NLV7yAA1Fwu7mqo4DWGJcbclvj1DSTW4OgAYaarYF2qO5esRRG9wp2haISWmTcBY1emWawKMAgC6
I3TQSo5o6Z9+7F9OLlU++93+yvk0pkDMkteHEODco2V/49iXCmIhFBUmsP7CZW7Jka9yz8lIprKu
TXuocsYRFKluyhBpKl5uvdOD4O3s8rFV6bOGy7DJxfxQWZ/hLUUX59Afuf99X2W4P2lL9Ao/fFjR
gbhCR1nFqpYI7FmleSaH0iK70nG+2eHyEnrUfO/mz5uw8pgQwUIObPBlQ1uJ77gl5k0mfeSLkjzp
wZmsdNjyu/KsRXcev51LuIupph5oqCuxoqJSCZz0SwUubqL3bMTZRocXzpgc+SXU1an9B7qayMDz
ZgO18VQMohCHDs32HkFTuoAMZ9KRHbEKV7om3SZc1mg+7u8mvYknK8DHg27YY3gdCKOFe4aVnLqh
OtkIUPjwGmj4nBXBNK/oO8ACUzkkSKPr1ozlHygRXkSF6Nk49eE2mFDsfnkCPtFrPYE7O+s8oKst
OaxJqxQ3K14b0GOmcYZ/E6W00nmTR/ZgM9uukszIawat/3g1PvnKeeysDe3mgi2hzI2JhtM8nv87
OfAUBH/NyPygDPdrJ42Jd2rmN7TPwOHZIR2yiDbZUsNbvtTi2OMpuQGfM8wJZab0pHYd0FArHNsO
uIuti90O5Wk3wQZcEtmZhBhPj0b76FnIEUZyWdtkGVA9E2Muj4Ytd0n2IF+XuGonY/pOFSfyfgrH
/B+j5ym8+V1dpeVgh7XNu5uF61SOJvFUks+iPEicFXi3Xuq6MEriZPLNCuyxTRYIKrA81k5DnqTO
V+lA3fuD9Cpv/r4dZVew3K4OAGP33t6M8Y/9SzfyDAD3jw0uPPV9XFqei/nmiaNNAsC/dKgfUvb1
c4l/OQtVlgVmMEqctufz1hmkgMIH8ZK4duLevMN8aju8Q4oXlYMqTwuX/Up4+Kmzlf5cvb+izUxO
rFqjZFJLGTegtAAtDAqR4kiK9uxls2NPM8Lyd/TPvfu5N+sOMafJkru0Dh9QrlrlIWMLeWAGf085
UXsR89067D9bAZcEykdQCw094kmG03zDWLq51tdvYp8eSWUpOO4Bbxm4megATs4ld7uqCyYkJsfU
JR1PyGYSfjl/KKL4Ld20B4gk7mEF4aIfahTfSII0fuVfA76vXLEUgxmTxFWyTgnpTBvfew3WFrCw
EEJhfN7QHBYKR4yuqqbWA9jlV8MuZCvcMpqA4swbQgCeIqXz+jzRNf9hUPeP3aTYfkgJ6M0AbrPq
K8by2zB0tyBPMCTMC0xWKhCr3qfyVSBzMgI29hldaIHr9wY1L+rlOeV80ziQhACzrNms/3174wLs
8QkJlWWASElkyfvyvp2SC7QrXw+SV/A6RVWDACba16OB4NFuJsurgI2kU04Ulm6+AcmHnJXRAhWh
TWD5hlNMzABEdlDpZHHnV7juLBuh3Q4uThj2IrP0TBhRS5l11IYIfzKgdVRE4gPiwT1s2793O3yU
uOI5pSlsfH/GSNxI8nYDNKpqWDsPneq9BVpLzwfPWkBktoSHxPfjMYUrEodNm1rSUmIXfEYukdQM
wM8hviv7xqh50MWzCJhkn/pMqc8j0KTBGVLdfOH4FVyeLhQQrAf0wjjQpduHlXxIpjugL4Ufg76H
2e5tFr2TQ8S7v43+CCuhukR+HRUCKbnrEjorYBz2a4ZmUyGedfk4SnwJaXnvzlinMwpHrWsME3Bq
NUlDrV98+9JAWW/WlW1ZExrCQgoZzS2SKLDwalGPRPg08h9P/0U2aS0ODxQ89puyjcxx4HqGHPIl
I2jw2a6hYcG4LYwchcntImVMvimTPiWejQhtbT2v56akK4QnwNw/V7Ce/bIkpiMjMr1QXEhKLX/f
KT1JcrXGYXgDw4K/RohussAYlA489Pe8MkC9rXpb0ZN/qrxO+efCJHB0ofbEMxHx7vem/2J4jsiA
H8G7KffRVoxnRxMbNN+CAu3KwN1Bpetu6y4Qlyct0mRTVurF1uEkIa5/KKaVvyNFlbwT+In9L2ND
nnbQpf1zj89wL4jziOCDMO6rlVrUOPwQtXiPLKna7Sciu5cSBkDqXsNKzVRDYhkyh6Zl5Wnpjeox
RtY0NfxOioiSUtmNsirdwMssMBhNRyXlR0XRAnt9kEfqgDE9TIOSYXnRfAhlFlBpbzmS7gaMX0C1
9hT8q3DYVEjCiDsvi+95ePBRl+ZGIeHp0Yb6i9G8qz8N6Z7q0Jj90YxfRqJ6+GTmLjphtwyz400+
FT9ESDwubPkjrPduEpEr3uzP5e/oTdPPy0FfAQeB+BOxNSgPQSOc5hp7n2TULH8G7AH9UAyFawdO
YeB5jJlSnEeH3GVvXVAJJy8BssgvsPEaEZAOtjm72OFW9L24nsg4eP3Yuxj9Y9nhF7ntIuA5Y8Bu
xZMoXlwT588HQWofLffLswCVge+an2fmK0vATsCgDOXcqfUqTZC+Smnay0P1hZujrSpEpAKYKbHW
LiCtdKX1BBwrcj/4QVSafSJ9v/Fs+2p3js1KYVeRm5fOxFhlL+qSDV7OvsR9ChzK2KWQUw/1vPa7
0VNHtoHV7x4gMMP6Dkf9+5Cafcu3IHsMc3RTmiewU0bwhGlz7EnVT1NsW0iZxfEh2eWg75jepP2Q
hH6vF1fwWdocacaS1KnYqsR/Wq1nQLpigRWloeGv2v0mUQMDGtEQ2uFAX6QTS8nRRej0xypvP0hE
oYpe/fX3VFeA0+PAZ0aGhz2c2tUK62zxxyY0OXYIO3a4+7Eja0KiY+uyNyCDZZPk6nJxENhqecgA
pNztapuUOSkBzXu5OLZ4uSWYfzNbv1QTiCHWrmALfjKXBf5zWVEv54titet1oe6oowOzBgTRRQ5j
++Bk2OCU4AjCP60EhXRDZOQ+FhJSf0EfDKGycx+rGhWrCZiy9kdqdheI5rBsrBKAh48Os2zCknHo
bRm/42NernAvdhGEOpq2H7G0TZGdPBsbza5H6hH2kUfz6N793XRJ9WaRwYVwvhAxYtDxnplFapco
KNtEMsri8v1KqPGtIavomE/Lv2TPReSNx9P9/rnBaHepYXeg1pi81Y631+IsX42NOv/TwbEphFk7
GSDcwiH1c2eQQ0KsxFf3Hw9thsVmpIWVEGo9cevieKUgQ3TBT0AanQJQvSDp2MKzlp8Ieoh75uot
2NpCQVSqXw1trY9E8OU4V0OJ3IHR3LpZPryIu9X9gBykhWRzKGsWfqopeEZljPPoIC6qI61p9twH
cOY8FAb1kWuWsIbnU9gAqB/8JQEKRo76D6z63lgBST2hvrKNlI18oX6z6PjfqhPD2O8wmz5XZaZR
9YDiN8cdADaF+DVHJanvsR/zS7R/AtWht/XX2scTRfFBHXsGo2p8jWNymSLU2q7Y85N7dGqH8j1G
GYgz/5BImkHsEIzN1mfTR9XV6jtlyGVZA0EMJPP+xOOs2BnOMLAOyaG75l9hPvje3AqstllS1Us1
0b1PZI6YCrAPuSJYg+LFynbrA2ZE2q5k4wsuCb1WtqbxsxLl62vkxQ0Kwnm6Cn+0JzW/uAeLPGkq
4FDKAgoZa9UJA6hzLXB42L5a5u5kM6syk4tmfrFDYe1eNPs9BnuYudk7qxC1QQhvW3EZo/nrorzq
wR2p+V7qGHconE48eWVcnSCvq+Y8OIm4qUnsF4QdoMAmUgE16ZWZ2q7hDCB8Clq5mIForw+lBzon
YTIP1RyFJfhBdlZ8weDmCjxbAW+/phtDgzbBD384tchUuZNiHkZHZNEYqaqxSeGzYYeaeYf/PB7W
Fte8Y2UdCOnTHNFEOcqJsanXl8VxOFd+njuGFJKn5vALEyE7vLwUyjIkMlbUlOWa4L/bjBrUvTNa
NZ+9NjJfA0P+coQYeXXm5V72qFkvVMplP1SHiBrfTK4jpylLdrv8ZwKznKlhwVPmownqtWCkOWlT
DaHyf6htaqbqdtRlIu78wtifrlXFdqZWowB42cpRlm5QLL1w/us65VoxqTSUHCbdyiyw6v4ZTbPn
zbz7/oRgLhbcRQnvtO2/5okEXRxSfS3XX6CVFCUO/srwwJfqMe+ItyyNvav10tGYejN7JMpM+fcL
hyPBXz6e+aZ42v+z4hH0gJ8wpUXS2olTOH139C3i7+gj/y7r7WtjN6mNhfTMlL+xWzHAIvoh5CG6
Rup6p+9bmPNnR+1kfhqrXS+O3+OeuwvCp0y1bi9Gso4lmXXZW5zF6AOJX/CB6XodKzam5wCbvakP
Mijt1uSYvorBu2CmO4/rfV+4HqehUG77Jvn20SEYvhOsqTVDcgkbQalewp8krseK3ZOHFZn1udrm
Aef4dKmxlrWe/Z6yf9DaSeNao0pH6Im3B9sPWqf5+hnhJlxqNXdTZNAB1QRHYWDmLZcnyJLZJUx+
nnRlBpeXFA9NkdJl6E2PJNf+NKT2oK4ns3Nv/FvyTYX1a1XjIACtAyz8P7IuVIStusRDUUGMV7Q8
gQNv0Vvvma6Ee2jeeYZCbxGvyxDHlArWkvCr3yHG21yO4iNhV3f9/oVjoGe5vwgkTPDQT7e73++H
NP1Xzhv69zYgdqC17oQc1SEfy/2DX+QdG3Oe+ERMzxfti6067QxrNhVCl89kQ7QNxTOOok537KfZ
3CScpPSYO/f5Ox8fyL49QsxtzJN/HR0J3bsiZKHJZ3WON2GbAxen/OttnyYNJmU41twwza/B/hxE
CM2Aa/1a7pcaxiN7fXtj6UpdrMYyyQ6xSyNtcefne/tGGDKyH0Pg1FNvg2b0Rju487/savLMrZYR
oUXdYsJ9DmjPUhuq80VqUe1imAkqFcCb8HAwYmobksNDkiuo43aKrzARaA24s76Rg0aBXV3m4avs
60Tz8lVl0axU5TszHgtm5ARCNuiMAADLWqCP7Cu5Ge4DlffYmt9/PsUCZnkTuAfNtcIcM5BBVbhY
wzeTmio/DBRmBGosfCe2gvGmiXyR/HHhQ8bIIyWl/4K09cNsf54jkaMOO0I7vSN9odu82Zw+yWVv
pEKZY9zqPVKTjzJgoiyt8xc6Wfc/jIx05TrATA8fqX4AaS4Df45BzB9nLdQ5zOI1kOAIMTug6qh9
qNEemN6alTWjeweXCogCahAb1Cjjr+kAP7RL+rBXvP7a2511r4xxrLIsBwsIDihBi4wTxgi5IP/S
IXoafgCofHGM6liBc05Rf0QD8HESwwONGtABtUqWokzP7/9UXovaTPE3lDeqlrLePpmKjJxW9OIg
NHrrLSMMVUkbn5ounND76Ko3mT3+PAsr8dSt4v6d7pUjKoPF5j8XtLntRsz7Qk+5JdHmIQFVVBK2
aDSCV5lXQIZYy0z+vSNN9kQYKtoXi+OQsu5GCnlDuNyanraMq7l0gm3raTHcU6BSgAf2UVV7agWP
7Aci15zwu/XfhyIK6HiKZVqoywV0D86QhRQc8Ylw5w23xwMFOwZHYf/uZxl0P/xKq7Bf8ETZ2dxp
y1RrZw6Y/X9I9mSkgdi1JZD7X0id0QHBertnkNokmpbYGEwovLKY9NQzoH9R8UiXtcInBMewytkC
ZBPSxG4r3LLHkyPG4mhDoOaM+qdvnVNOf898tckcolhY3ImP/SN8ONC9scXmep3/+bjxZ3k5hfEx
IzaWx9N4YpVC/MHu2ei4dxytnPTeo0phx5UgdeT4wPH634Uku7bFquCfmzWmDPj7Ee8LwK6nn6dn
9qxIyjjR+ufGemlpKxmIx6D4QHiZ/QPf8XbKy3ZFcvWXSgtrtZ9Lg4LRYxEai+8WzcBc9jsJOSa/
6QLPU54PjgFK6u60VGxkwLaLR6BUOzdGv5XIJMjFJ5EHVBBUSfDTA8nk2PN3Z5mufhjEpETnhGaR
k752UZXax0MyUJTLC3ynMR6BAQFnapU3xTWEAxYUfA+26YgYVFK/KohULnYebdgf6Pus/DZEAdMV
im2e0EtxCvkz7GXoOrUpn8HFOtdpgcr/Svueu2ofmEu/MwDe6plPjm7bDQsP9zhOTeQ1ieR8VY0w
AzZTlT06LDqknuwYXjYjMKikD3rUWvfjdotdme2gFnLBw4la/yV2Ho0gfdcct0VfKQimLY1NforR
zMZjdhM3C0PQ1FXJvNgtsAQR5gJEVac+HnqyfcoJoV3puGfQNbnvRiXVwiMntwEwT62Hn0TFuSTe
FGsrvA/ZN1F84EZym26C9jjGEtCD4hn0aI1ok8+SKiICLj4c1Ri0kWb2TjN7q1vCk/gmhiKVL64/
QJA5Km5hgZuL2Ff/t8kPJIHSKYLqQF5CR3Hndttzk/YwziNeJEZMwEQPUH4FT9xk2CyAQvwlNK8C
OIx/JRtUnL2x3rjzT9+1WGAGjzNxSM7PdCV7TfG+xNY5pEDzsDS9tixpVVnFNlCIarlN9rZ8JgkM
/uk1OWV27/SfDQlVuKIIRqJuukfyYZegUCemTrotW+FC6vBVJP/3/MIn/IYcf43OLjEhaxM2QZxK
wG9KqXZQ8pSOOir+C2mz5V/bj/V1zoCXlObdlEoJfJDV6RNGwmiT0pJ1Zlvxmc/wn/NvyuyfBnPV
oKHPdy51WHNvjyrfUJqlnCVznlDH8gC/OWDnwNqN6GYkrlxESeaDdcMkjmhfNtCVmWe5pvteXIK7
zW0WyxKEiCsMHJ3FZrL3h8piF0ZprXnTnkqL0b+Jyadx49EsMQAKQFjhOShtiV6vUbLIdXPS5RGD
p/8j9PA55j2RpzudULFhkYPuZcfocbLwu1h+Lxp5lmO6BiCElnr763yd8/wYnkg6kEEn7Cr4vKBe
VQIgzpnPyzjkT0nXUlo8/ryzSAlxfCzqUBCcSO4i+jwPbU6iquFXi2l0VV+UQFqSADb2VTAWE1at
QEJjgAY9xYQ9vCPAPnIBEDVPgPww/40IUJtyhLP4g6r4e1gJvz2C0Q5Wl230NzVHz4CAR+foOpv0
si9koiyZzAnfkI7XNESuIEJ3p+foUymW/17GSM10Sa8D0srVbNYiT2v4F94LHf4q0q+fd0o1EvX1
KHN2mBDRHRy7eRaJjz5BfvbLK21uPNt132bG5rI3xB4M2/42dpxZQb11enABPCD8I9pulx2fR0Tq
QwEjtWOui/4io1ei9ItwNQhBPi/xtFPissVParHIYPNkfVdJFJo2KHgERJBc6YSwejs98iB59ojo
tstFbaE/mAE20izXjVTla6qPDtzkjvn30GskwA/+3YtnBMt3Y/Ml13FboR+q+nChhBqgOPtHsFHj
OMnpTrvFznc+K2FTFSNqBUkFKxUK24OgUikeijYo6PDZlFam6UEVdIlLFPzDoJEGrv8r0Z7q2GwJ
v0Ap/nQSbjU1lytuzX+8tGEtgWwuzkrorzuqR32QeohswRSkkIz6DkK1kBz1hkYr9TfzU6woFsT+
3F3DgI4jWR+kB1U3s9ES8wTyO4D7ysU0rrlB6Iz57p3+5fGqzEMTD5T1ZggoyDa7rx8kHECruuxD
jPcHlu6XPovKKTuPMnF0kHGrn5X0AMyE8CWz9CXgile3ty4N+kqZhIoCGhWPDmpEP9jhC2YdUP6H
40J15GH4VXsBedJJ8yB/al3YojCo3HxzNRk9MhJZQP7Eij30n7VNtNuVvCgetZSH8Dnvwb8wvYa6
qUq66WXqaVEmmzx1xX5kZ+cjF6nlt+hZ9qPTBUQF4QlOwzgeo+YZD9WOzpvZfJG/HNMNtOkzZ475
1wa8wGDNreYLXYPLbD0o+bQmSkxm55HmoXVk+Ih3AZZqRv1ANURwRBoKm1eqQUZ7w31Rl7lZM+rg
nVGfwBZM64NA2NqmoD6VMQsfVagikb9u4kopYmPX5dfVhIHCWuqlh8XVqGE2c8k9I2i182mCEgCL
rRYHr8qVbWaFfCNSilegereaUeSeHLg2FuF2iN2dcp/TF5AMr0ucCFuDbgaVzAzXvM9QREK763bW
Tj84M7OxpJRQygzzBSMKsTuXioAoVPsGKg4K/yFOgousuEAbOWZD2PFMCTHED14b0yyA5+Tml47p
15sdC7+2zkBDB2J9hK83U8k9WWa6Fz7McWIv6Pv451aW/+1t4Aa1qVAyIYiB4qOOYBO72zJrOnTO
iL+ZfIhWYkL9VFBfQyrezqgZM4FDJBgSMnX5mnIMKve+aYO7Oaz5sl/CXRX2oksbhblxWGnRYlgZ
oEKMlcfYo9n1c50kS5WHNhr0c0fyBFo2gCD/YXlQhy7j8i84uE8LNylOteH/2LerRbM48unt78w9
UWCO3ECKMViNl2IgplVdNaEUVTl2xWiU4BkngndfkpWp1XXj445D4sdf9wJoM76KwgDqYZVXOuO4
DVUcwD6ys8TTNMS7kqHJZKskckAnc/pWLuCgJMT7FvVtTWndvfDBe82/2+WvU1yD+m6DpLJ2fbwj
MD37cxXOkTEsJB+BzX3fAEA6T+fmB5Wz6RqWD4bW0kwk8xPRMWIqCqlscg0yQpV7kRqvWOSOy6WG
le/amaJ4T5KpvBWFsuSyDGIV69l4V6dnQvnOVjzzMhXC1DO0s7+PjFb2TEGY6TbGrb0h4dKcYiJ9
9d4A3l2Hf5pCfkZ8PYirVl1oExOsJoSfiAJxgOG896+QGToZEKJxEvDlZeDU3+MXL0HcUb0YjMBa
7eKAsq/sLZWAgmSu1m+AtliD782rZ8XNQHcqv3J5I7zHDRsAonPODARkV7jjfe7jGDYRnbR1pWhr
8930Eus2YooLhKazrpWq+1nS+mAoGa0wl2qEQdbRAsMD/npX7FlgtX97eHbef6uSJFQPjkf4YdUy
p0671yt3qZfFLiQAzCyA/c3eAGqqgEkq8T8ICnsC/lvyRMNmrM8JC4rDhaaUcMIvJo6I+o5kxJux
I6JAFxgDxIwlbFUoEJ21uxY+SZlapWDc6SDPk3oiaaHgpx1Ij7F9RbLO6p23Fy3Phc8uQUNH2Iz6
tJJTihxLtJKXbrV1TqUCKUcr3GoIxyt00V7s9Vc/0r6sYGnBSArWLwTB5px0g1i3Co1k9rkJ7X96
alLxju8nwUNImZoUyNdA0GpAyldqKJAOCUYE47Xouk8agddUlyWrH0bELkO2wmSCMBa1bChgJt3T
5fECkPYKyOzQpb8P+G8djdWf5pR5kURNUQRidNxCTENNcbbHZ7Smk8kHuSzZFOe5xiG/uv+xy/tm
i6EzP9oJEsuTHNNT62Qx/Ctbs0Yf4Sb1Kbth+vhXTTdbQTGBg52PymGPBkQ88lyL1PU+BTcLeAQp
1OTonvKQeV6MI2YfC5uCC99kGH7cXEM9O21EFmcqrrfe3wX5e1zwupO0lgxgd2K+tb2gA0ddm19L
jD6SNP8QkYG4+9PBc9D2bUGxyMdzh/+6DNkC9j234Pg0tCw+FkSD2tgazZZGHye7gauUebsZrM9+
flG8nV5rxpke6lXjgrqh6zgD9pIqcWzAaRSXIv2QSpnUJqujeuZroBXmfqW3lv2OI1GzbQ9eNVGZ
fSPukYs75ozjctRrHFQgZ8O3MBXNtqe7Hezav3vp+4190IPuDbNiaNbUkl7ZkodnBJS0KTCx2XpB
7gFZ06rjeC7G1o4EAryi5koHqtWrYle/Dr15UZKKemUGIt/4np3tXO5j23IBUjmjToFKctPpqcWa
ZwtuYDPUndzXJfKjLgd38Y2aHxl8ZUoYg+pwr/gdFftONOmb1O79/SOMKqoU7geC2/gfDCbAq+zc
Vebzdbq5JxpJdY4duTHg2dKtE+jGFj3VOcWQA5u3lshaZC83BizbXGmvl9Ip93Lx/cJ/iH2bikm4
o2/MBP44pZzy31ZICu0l0+kA/N2yGxMEBCLbK5ifQfOKEG+VYM+x4rWYQWhdb4uW2pm0JCoRT9+v
p6uCrGZgmtKjMhNUOCPdRxLvQtWJYdRI2Xo9CY2nQ4nOXOH1uJybey+2lOlI1DEh5OhSC1Ydf1G/
4mZXchQftUSMiWcmUKvu03B3IyGs/0jgU9HWjsdbfpLoaF3z+rnekbbl2S5cAZ8lkEtu9jYIPyre
LXo6l5vkUJPmYy7Fvt1qgQvQ5f0oNv+yifkAw47m8FLqlZui4FkUU+KXjNAGybuvgwL0R8CicGxW
m/JayrzqGwIrVYMxfJ11MFG/LeRfCPAlQKMeYeYG8ZXhDXlYB8cGCQkZL7zR6qAdLCJcy7iF8GRk
hB9xKZIgLaPicMwX5EvMkya0qs0BfOpSZ6D30UerhQzC69K8OWAj1j20gENZJMEH4ei/CoqR0OsG
20AY99p03lowNQkqg5DxRXw98pzX1CO5KCKHDVgMvvywTTa33bpOOOUPaaExwRdcQ6FARTAZAAYE
gv/+GpvA4QByEJkgRS/dwOtR9GL5DV24ffOlhuNOpAM6nT9P6ruJTX7ycKyEIiOJIarzOTaiJ/Aq
BF/xW7h0DnkJ/8P2GG5Ecd+ikoS9+aoqhNbO03MPtKl3sqKArmCBX9E9J+I+GNoWZsYapYSZ2k1Z
naw41LhojU/t+Ejwtlfy4XmGzRPFBAAVCJIixeFUDQNn3I8FJCTH4T3m+onYJ3Ih7zMBHr0omVGR
Wu4KbZHfUauSQDXJ23xFevciD1+7Gqb8mZYxnrkwplBN7LrPMch6/RgHUE0C2/61sh7+SVu0bcAu
HoyXd53DceBom89CXNhDZWTryK+LR4DIEPGDF221Px3vKGiS3apGONYKPnPa8P38+o/22PESglGM
TJueIaGDFnnBpU40cQahXu272qAsxgy49GHDGnPf8cExcZNnOUL4TL2zMaxsUhwgyqmTwPFrjQ2F
Gk44eyzTegS7b5r/f3Si5w3+AXgs4PJpitaOA0ngOdD4p46S2cMh4GIkWUMV6uITdhdah4EPfG/5
pbLzY6NwyUiMzNLYyrVPNlOY5NoDGOBgLYzt8SudREwYGZJYv9hCADl9BCxk7QqW6TZ8DlAMqGT1
LKIg2Dg6g5jYbYcJJKruuvcCWICxyX6uFQuAzXEcaH7SLW6nEW0mFe0ZN8HwjMKu45/dPr3NTxaN
f8v6NBFTslhYHVkccNmTAib6OOmS8ogbv1KEKWsbZfkk3s8Zx0wswnryHLQcvYUC7OOYCTYWr6Mu
c98wqZBUuurneeFGngdydF8DnWG7Nkr9q3EH6zr9N+A4j5rQ6xs4gYbNGul/3qAZ34WH/zB3Eytm
Cq4rWlYcckxSeD/TbT7PoRIhLk8wXL1kAHesd1yrvolTcTgOT/eNTDLjmdIOWpjSRbt3Ug0pkmG5
AC3lEi3gpjVvAhL1CuJn0gU94qqdYCayRmdvmmlAzR3YbVUaUH+h+Uv5CPAC1HWccF8yu+kCbC0k
xYOEhxlzrHQqO8XcgBIoCjdxxtJ4RFtimk43IXH3sXJ47LsKjglWdhLBVn5Y9qj4tDTmYZp9+dDL
OOpoHGXF31wHwiggaHPlkHrKJP5f21MsHP3OGKVNEi4m6TN47/PFI/fat/gVKM2CV4rwGy7N3WY9
JfLr6B6lJoQ3qoiZF2piCDKdQ8DReI53BMoA51ir+ndDstmb2zz7LrAFFs2PIGrzjDZJlyrT30FI
5zwMSZpiTQFObfdEwb+vwyKIPAdtC/0OlMcA1DoX49uYvCSn/O2KkLAgHBG+gKNIG1eETTTkka7y
KEg2lnQNz/sZQmRoGivq1zNEogqT0EhMM0E9Q9aSxt9OK4A3RwAc1MoYDiuUFL4w80oNXy0ykbOc
X1J4tI6A+SHVChfz8EyQ2FZaQlMxQ833txk1CTUBtyM0ooAN+BqAPos3iODHaHvy/LB36Ze4Ac/p
EfH5VzLIc9QCLD1/x2uZ3xl4fBks64PlBwbuAK70HqdNY8wO0+pbXFaPeFhh2gtEJtv7MYIGGbop
qnTq8CZ6CDaC/MNrdovQA16KZMFlQYabfmajm6uYfFn4WYRkKceC5Ne0BMDJjWvmdURhwCMBe0c6
w+6TRD+CXHHwS9KGlXV0hzOuFZo93VL1cHsrPXZEBEA8NXqs0KpTcc9W1pYl11cGAzh+0SUb2J3g
oz3AYMgX9FDT9FWBlkNeca34h6zLseLTjTmcNetC7CGKDCviataYPOdy1w575XGf3Khmy76Zd3PR
Hk73pF6uk71BquPxA2P6sf4eiXH2k7OlZpPBoOpcEADDgYzhWPnNC8lRDkZ0c14LNWBDbRpm80c9
Ym1D6jY0i64tJIhenUxzD5CTIAGl2lh6nLXQGlaWg5hCCjV2mrAqlatWHXPqXFL4RPeDLhYShdzb
LUyyrI2drsBLkczS9KilO1l/TrfxbLC9n0TDF+cZmeaJrnXTkgfrghJmfsWfbJMhwu3yNfntpiJ0
ssBhFBjVyj9K3hjMa06hwc9XicVLvaPCuc0WVyfHS+7+QrN3nTbaOeBGu7bLO0tpu0tLELyi4zz5
nyQ2j174yI9RRRTova33NY8dGnQqeK0vCZv8+GUHCKMn+G/6++shbALGbQyjhh9sAtAwWTn+sfqF
Sj/pPFMrbnPbzLhD5797tarKka6nSQZMfS+45JclBE2/0Te6+1dHnTNw5W7b+Vs5camzc3pm1j86
aWygbKjJdLUb9gZIhTvrU+hHo5OiZNKjPB8sBGpQAIB6N9H49sEZw/fQy0c73gg2K7Erd3jkxGb5
LlrH2Eov4C7NuXtjnsI+mw/zvFxXrCZBWbulZJrGNnAegmMX6KjkTwQJImBmjYTaL4J//Q/NqFHr
yPd9lPzDTi46oL3NxIwrvJt/3mQrAqTwuxMz19FypsXiL8PYAHxJof7WpE/377/NqVpV3qmrXwh0
wOlKCVIfFtDpDiYUWkCpzDM6iuz90uTHdBAGCCwcdtsRBixY81qnWTXW/v9eYYzWPhrj+anzp6qa
TPhRihj4/VYv4uBn0R2q8ifMN8j+HcKyBsmX1ExRhVE3eCarXwOlBIo7NgVhqNSorowf2jyU6awT
1jHWY+qZTbkWXfz4lZm7xWXLvcuDQVC8yAycbG1bYFB3H11dYydUSZRGy1AiGcfAvD6LvKZKQ9R5
HGbijIqG2+pX4xcRR8mwhU3oExR4fepaSC/O231yQW12bOufQMrLxyQV5g2dHNY4/ulhuAoBOVzv
q5rde6NfpcudS2g5QMQKkB4XJzf+CfpEZUCLR8iXHhLFrfhZrGyYwcV6WIZa55wcE9QvHnFd/MAD
zXHgr5rA4JZB/SxLxLv7KeLcnhD1Lp/QqS5LV2TDOi3NaSRaZsH8GdcHHFqkeIBE8JJ4fuTsaOgC
ltCkrI01WPoGKISO1gPSBeLBFu7pnQbryAA1nqhwJxBAIvc+Xrfks7Y4EyTx4cS7xYzQECEZTeFJ
Tiz493zvG1LKpVoUNweoxiqWGTt5VkxD6JUiONEapNs2QNnNQ8dwHiSmwUG5cpvEHS3PgtwFLxsU
1qRyC2uHtRTkT7pjBXxiYtLPXv6A1gC9ciSqvPjcK/M9zGdFYrwElOOy/uKqCvk4ZnhT2NuMG6cD
bB8HxuSulyuEo/G54U9MRj91Dy+BEh3Nwb4QO/VdHPi2VEM5DY08a9lbnhmY0/JyH+GEIZO4AaQr
RABCZvOoEFGqQq2DVmEdVES2fbXlEmR4y8D2MAjU/VcLBxPr9dKzEw8wP5/gY2JGvQtBuGCOu5TZ
mRFflLxh4oZKivI37FOWx2jVNu996NaIvy4570di/NnhNF3+y7hzAcQbOZ4eNXDDVRPTSe3Bw71j
q/l5os7tus1ai73OBl/0GYeUHupGkzQiAeOU0+r2JqmAphNBlBUMjIKEgSRP1RugXtEy6APHZbZh
eE6xZdRZqrzkfHryh2012I0FEHg/3n9D6JcEsXWBCQGH3Bw8uZ7aFJYK17wXqMkLfJaT/qDX9st3
Sf3cjEEzwoEIk6XAQZuJ6VujEH9J/k15HrnCmGpBbUdY8H4RApWe2kZUlU6/q19+uezKKXMYQjoR
cLoZ4J1KApuq9FyAdPrdKA8eFx6/wtNVK5cnRGcIgIUVhvByDzbO/Zv9e21/bpE9m0SIMslgqBwF
ER1/S9EZf8vPRW7JNeOHsfx7nn1GVaODmKUPTBi7YhX/S6+TQ3nBzo16jHDJDcFHGOH1428PFHnZ
Fa+NeGkVQyU8yaH3t9RKGOpgLATz0XJQFKKYzDMofvs2t302z8cLQSbIzilSBo4/GSxRwPf3rhdM
m1YAJUVIIYoSgCjWRV7jCMSmGNs/0XgeEvjC84v6Ogxno5JyK+Q7P4JnhXnMw/uu2ydl2jCmVtSi
ZIWuXkykCXSOEdv8nd/SkpeSMiy87VGJZQca2kXKneThucnFSifMqMVC1LQXMkkY4VgTo2U/P5uf
BoS2vGsDalNbEou97c9GSwjg3tr9oL3es3KOP3KMd7Y3tBRkKjEbCTRhTKciHaa8b/CJTRscOO22
UGl9Z0btdcfxMUaT8Ihz+A+eC8aPKgv0XLm2Ha8g1lehoYl3XNJbfnfzF2FGoVkzRX1zuyILq2qw
mVB1eeb1xW1blJ8FeejRNS+QWmLm61nRLMOviRN07tgXe334hsiktOp+3j0E8vqzUqs0rQET5lCu
y1kOFuTmC7iMO5NnFPDfmu5NjTTQ24gkeksbqb8ftI4Q54a36IhqZK9+f4na3zmXrRsNZpPpgAVt
B7YSNOXhc8RsBDzNCz8y7TWcJkdQdpak3jZ9eO3BHsGEnXzmASNMG5mZ57GLtRPWYj0kP2Xqypt8
Fc/ym0C6rudgqWCcfi2SgZ9rn24ogJfZYGmQa98qmF5BtQNnqUtR8kONOXoXSqPSt9sVJwXpTNbp
irrWee62vsoF6gaBLi72+cdmDP+zVqs/LIxpfs5DZB0yRFLMRJVttYOAfHwUk7iI9xZtrNpVEfs7
IUsgaK1zwAZQUHY3jf/mszoP4j3Q3TXcG4Tvqtmdjl6ilXiT/uUvipY4PIzz7Z5Z2cRiK1zXksi3
AHSzdeYxHjazCjmFcrmOZhxFnkGKjY2m5nGOb9fEgqDqry9JeOAHmlFgMtl/oE/q5mAgmFweGEkk
Gt1GeXdXsVQHrhJYUA52Y7Pzz+SUAEK0R5z+w4njxE/ac4uuYi06OtV9s6ROgKP8kArl8oJ1YI6V
voHsjfhVH9ad79S7E/QEN8dMCo/QQs/9d+72DJ5YL9iCKBtBRkQrpoj2yWR2/cA+dTZjC0VSl8uk
Ox0mJIY9HxixKbt3tHri6kU8lHqiQ6YpuuHiins/6iCjyGJfEEaAj87ZtGdhO7F8JiDdasbNl0ue
PVoJ5OjFZnyYO8TF2w2tvV84U0fkezSV5M22FZgwoby6t0ZMwtPpoU8lfjkSztYsnNs+BvycqKZi
NYPRy54qqZh4QgpJYy+AtlXVrgZf3s8yjtDCt4r1AExOtffOVMJ3Ai/o3ad9LdgulhKIzVobvrEk
NTYSDGtLGTX0VUmJHRRZywo6PfU8ZFnKqhgqWztc1RiZhTbnqwUCt26/ec/nAg4co8XDSNoLNyoG
ok1Zwo+z1k2gEqaLVey8O0TOvZ8RftVXvYOe6NOjx13MO3a+VN3APeoBLHzXzLsxDYsUR7Zz08uE
RQK0UPXAL4kP+Y1DaSPLJTLuARiBypTRcJwoithriQYem3pWogfK3JYCf/lS2dW9fpy15cwnzqLI
8cpHCr+qLP56BLFEcn2uxZzge7Uswuqs20DfyumKpz0wg7QUluM2jLU9jPff66BZQnGaSVifWIg9
vJA438ccrtE34fxoxPGJJB22CTexouT9BhuFQ8NtDFw5c+XDZf4rkByTwzrsSpzSuqDVQnnyxMjr
aV0xtSf+RxAKaFETptDvNevoPQJACJmYdmTYPXUI6t4dzfQcvwD4F/Zd94qPgoTJTKMBHKTtvquf
gLHg4/pa9TzHyCzzDdkz9sRx5Fi4IEJWrqrr+ERqXHUFRarxiC2/GLPwBgwbn+6RJFPbFcUXBiIB
L8cunzp/hKGVJz4S32gKoLkW7Tc1x4NzjGW3xVmQDpRK5bZta9QCBkSlbYlB1G5KxE3BVm8DREyI
/iJqCh33NOQ3y83xn36BPZzOp9IBi4yHdOVlnGzkmK0PEKzp45nkyh0FvmaoUI3aTnNxi2RuzwKS
H7emscIdgDxRttc6iPgksR2ZC5ThxR+1xTjjLt5W/ycI+LFYZ5ly2Lit+IbXgqY6muaNX0L1Wm0S
rx6KOAO3IbFLT2DW+GPTAPWk9Y6efCqe7vbmHWDWBbMEz55xvsGTkbIfVU2HnYrPH0eQ/uBUvzCA
2jSruCEh8DF4Rk0SbPe/FjCiyd7PMHwptWxQpVZkNzxP5zoxL9HEcaZJbwxaVeCmw/mLbHWvN0yc
zN3V58iwgcbknBJJjP7MDiUffZAA9hsv6K9b23u90OUzap8ynsNnuxEp0BgJ4IuK9804aKEwzInj
1Sas1T6qQCSsOwCwTabWv65newi56JKCHUCiRkKRdnFbGho8PUFho9ZfiG8Ykl3rNGUAt43Rb8Cv
7++E3b2vwLD9GjXGaPc3yYLbdQeg8nrp3OqLA5lq3z1yuLugp7E9jZ/P66z0E2ADjlh5tPKmz/EX
LqPMbtL32vmqL8X4kzVWVtNl2l6MBVrT8CBRJeEqH1OzX7S9DtPdSZcDXMACtjq7OQBJzzEAv1vI
9YH2SSKGa937IzcRYdW+T+c5N/CeyZsFbozsSJBvo67JE3t/rwahe6yGDoJNHuJWv5f7Dj8lVvY0
yeSDxBZiWGEaxwug4mvQwMOnOK8JWPHwm6EcQmPlrCGwwaW8BL7QEklWOTsleiLNy6jQbv2NXJsd
Dru/aZWZxbBYW8yAtboR2A8s2Mo+Aslu1ds90HvFIkmXx4AMeEXLKRaOZGlrEhzXMakeTSamI9wW
JG6wQ3amJnU6AxlHVsgMxE1qOjmeHagcftwmTexneXODWgaiReBXEpPI3WSBRP070mtHJrh/YnVO
/dhl1oElTHXSorAfIlnnj7vjmS6K5f/NV6BFDdATUbVPwyMsIVr4/vOT6iOZ1YoildG3OPdC0JLN
fAjFmy+nar0S9j3mgzq5xrWOZc5wGS5mdw89iyQF5dTZuFSb7fpQEfK5/c4i7tV4btJqYy2AmeMF
hRMJZz1VROLz+0Wpi+Q9pnOwkwpQLvcWc1f+Xj5av4kR8FDObiL8k9KHzwZ/+Y7bMmcaxZh7W85X
tDjmJeVEQk6UpW8K3VANATOSNMgqJlI4mpgcZFBEzieg6tc9JWcvXKpGa/SEzOEvcKVM06Sf9ua4
SqRAornrHGIintD/S3eao5dbA/ri2l/8NUjIPFuHMWHeQjgGEzFhJp8LAUlwP1M6jG5u+E9QYzu0
AwuOqX+va+YRkanj2xUQCqxZU7kxp2BYy1qTp/asPfqA/sAqzqobux3UQEE+3ld9RjPdYsLlEJaZ
kiAJX3Jv0vMWX3hEYITEBHoF1wvgjU7Ddrk0/QGiLadL3aXzhUyMXfk5XqcuUT4c5XBIRCudbKi+
LT1Ic8NlAMtEUId1Y3bvaFSUFtFvRT0dr/nJ2nxn4+jUdQdhwF4tgIELZI3Lh2aFCIH3/KjmRTP2
bYqczhgLwHlqshJfBY/lCZb1bWlxnSZguuRH8APQggPyMUkZ0CLdjmO1Fvb3OXJa/Is1RBzLYoVy
E/IqXA03+ahrlpAMF3jyRLWzzgqGUGk6C0QnujMvydgIU5mlh1iy/4SgPm1B4I1vwuI3mhib59vf
4EnTiACrlABJuaulk/MAX7hykIAU+xPwOPEeIZF/cyQCfZsUzzH7GMsAdG7uKBnYhlApyd+xmSaX
BU2O2726vC+yZdsAb0pn1kxg+Dj/2r8D9q1OJJIRe/uC0n59FfCCao1uLlNjspPZlOfATDQ2cWd6
uwGu7rPWKDZ1KM58f3782CTN3bZBc8CJpXqgsQx4llvbBuhfFHepv2hvf2QT5hXzemVT1kGhhhXQ
Bu1K4wujw1ssFNn+Z4mi9aLUTqyIc87XZ4Qb3rFah07kL/Yf9nFNe22XNzB81fbeg8vjUxO43rUY
K9XYpcTpL2y5RyXnAUV9G7dfA9+BtoQTyapDBX+iKGArA8yn/rTUPGs6DKeFrwCoTPAter1zgzkH
8Btid1kTepOZ/BRgkWIsW1zoP3BCIoZT037TQqI+F7DYae+nO/bTi11TMhVshspqVYt3JGvf5W3I
tC/D1dJBRjOw6vRQ+iMRbzzLo2Kt13VRQH6mVMGRUWRUMpMI1+1K4dy/J72teIEDxLwUawm+e9KY
0R2KSJcK46fgpAlRCq8waALmFZJZvrVTD/ZR2oyRGTf/GMhDSc+RAg6hux3GrCFraO/qEc4kjrm1
4VXMb6peheqjrLxiPn1Mz/7vrlrYrosulLfImfybYaypURHdfVvBZ8wx4LzxCcSAKIjVxCcyWURp
nPWWTw4G36TIey0O/B3Y2EHgV8l80Ud+BOLMJoE3eO+M/Qux0z5GziG7Ooi7hV757hDZqO/qYYnu
T28m7Xr6BMhUmfvReO/gTxcv7GdE0MpmqzxSxRrbsTHJf4bwMoeW4/G30HyiTikhSmb0I3U2iJyN
c/pfeCDoDFVhOrrw1xxxR4abmlJK5pJzOVmNzwudxissxWkwOfPtA/njRlx1VFfbySZI/M5dVVD4
MbuZeBNERpq3Iz6ojAYpnq89QESq4VwSSQPSwc8I+Z7MJ7JHTiiCi8eBnqdkCEJ18yhf8ZLkQMK9
jR+VeMIwqcnOv2lC442Gx8eEY6+omYQjmC7fs62wNjx5Hjw/uMXFTpJO1pq52m8EINMIp+LQ4uh1
bLl+WSeRMQV0uNtH35i15tOUb8MMbfL/l9TwM7n923BdmWasdSNnvnAkJYH1Ls0whkLVpRDHFOnm
hSdA55nIOnCldUKYhHqT3+CPrc/CA0Vmd4w+IsbhQ8aUfM2NDIlMCpAAuW0euvaOgrv60o+3mz3K
RI298cUNSYFUInWaNxInKbSjghHNUQuqjawYBwMIsJ3xuE/6YPVP8oHAQULMae5HBUJOQ/2cjbur
Mok7D4ygeySdzPQSvmZjDOsxlk9H9aGk2my9q6FtGPQgq+JWhmrHSJWgrw6bV1wr610Vj6BoY9gu
2fWOdAMculZh//+nYZwSi8ZQUF+Qd8PY2wRKzSeJRTFCdgxwT7lMnfKMgtuNKM1JucOViCcmiTiq
ge4K8VA/8StKyqY2Jk7eP0gm+Np4HFO7hiCGZgMLYKTfNS3OI/PDRKmi25ypNV9WiP/wWzWQKBgm
xhaHhtNdDG28x1e5Rs+4e4cIMRrbAYH/PO2qW33WDLKitt/igkdtpg3XFAIavXqarjDlRvo1UOkS
SLPfeulV1CHyFPyWaHoPv7is2Sr01Zunx5t6AqOCb2qFrOPmwjeIts385a43O/nl9K0FnktuL8dD
riOUcqpgms0d1BWSgCN2ySgFAWj2h2g3rvl8DsnTO13PYB4YwvHcZMNX8aMHdjxr71jnc2sdNIb0
LFqb2vRBHiyPZhpHoD+/j5ycpMfUmQnAjQ9b/O7nO/WJo8/b6Jv+/QhEUGMzg7RLigsmPm411qQT
dc/o0NTflh3U+01ZTx72pnmIM8p6fvT1z9VHxqxx7MhKe4wcYhluKNOKqFkgNy5WbECaT0+4IPSK
0myNI3L3G0OM8rOTjSe5PjxCeIirv/ZkN70V7/diHqll87BZGDkvwmF83z6c1lBUURrS29fvBV51
qNX6INYP81NZoW5RLwQX6+sJiOwgvss5wye2lkYNHCmbYfEx4+qWgxwm5FCwWRqWnv2MeqM8giJd
Btwc5/zpCDJiBBdtpPPT2d4k1b398GOfqC4LkoDv+h5kGMAX4IXLAX/zADGi7P0we9WaN5lGgkMo
43aDfap0effoOx815O8hEnd48C97i8bhYkTlVQNWqXkKSsHfxy/6pKUXsMaqV5PJ8hGm5goBbeo2
jARTQxq48ueCyKjRBHLas8lfrFa+Qz/e8EtdE7D3lAqbLE8uULGSYDgC1yBjkQd0LqzUjf1A/UqW
SnsQjdGX72nvcx5fRv8+4bsv1HOy6+G2I2PDIfXrbSfXkFr3P4N5HPFlZ65hQGqTrwZfHUqqacXZ
Wv5uXQ2An2DhbkldidX9ZmzIewhDC3et/QbH+iOZAg6srIxNpGBZbocjIAqI2T3Mms32KGE0AxeL
hsjZPseYgNyaP18C3QzXmXMglvxznnTa5FMkH9N3aMVxMq4VVeVX2Hz2f5DjXyg4a7qNRsl3gtGn
4t+8guN9G+iAyN2WLNCcDmMFy+BC5p7bqZrogw/9FumHWkUgh3tmfW44rV2LvwyhaKozVv9Y0vsC
xB8iShZ7zV4bLVtCsoZbwqkQaKLl0ZbEkYI1HGbask57qy6ZdT9I8HymchOPkWi+hnPG3WSDiGiq
QrbymycwQ/L5i38jPxOBVYklgxN6/T17Ei5ILjtBVlLH25S1SI3LDYS/ohuDQPNDjuT39Z4sCZfq
lCxpM4CKLOYgeYoeGMm1IGLFl1ZyYsnHpMFJmL/oGonm5ulRYhfS6Cie9vnyOTjCSpiZ2ugcqbj5
TsydxaU572MfQiPfT45dG4Eda2eORlRXqBVobNzZzdGfjl4UVm5rvpV+wVUiz6gehs4JOOfcUp4C
FYUh5n1ZLW4+wooRSB2c8uKZdJcJucaGC92rRaakWKVSE2ktBHAx9ZOm1CaPtBOt4pACxEwyemrj
+3/DTp0URq+c0nlQ5ofi1MY0agu56Mr4UWcK3WTswIkR+q7FX7gxmBCB0YIdT8mA/oz02hYX3NHQ
uHgXWJeYWuz365BwwH0eh6aqz03mLgVwBB3AEdx9mNoWLdMnIKlLZNCBwAvqz2y1Pi3neGh9E3x4
keNY8lU7DrvPoFDBJnv6CIegdjm7LICWgd+QRZSCpZAmA/EFpUxqdQXz7EAj+Ds6MOzGWxOA2o9b
7+lXjZ6CCDorTWVaOk+Q7/C5cpWHJn8bRVSAlT0cjbAjmTrVBAjviprVQCCcnj6nWaQn7ZZt2hit
Gca17hRFWO3UT5wlL8l2vnyrAmOsL+VYv9bH+RbCv4jm4irVfnF0/Aw6Vrh0hGAa/UbffnUup1Az
8UE0o5be/v0W8oMQFJWMej0WGZ4rwfztvlqt7cKU0nBMklv4XE1OjYP8Aag1GjaxPPV9/8ewW5VM
3Z+0r36TprUk1w3MGyE8Yrlg2pVs8TLWtHyftIU+SA1HDWDfPdyxp3MqeSVGPCUhQf+MKfu9v2LS
S1J/k6DPY2U6M81PWr84Q2EhMuT5uDfdvsDtK/Cl2pYZ6Ww59NaXbYffqPIZyYjnJlnbV6JMV8Z2
/18JwKlMBBtR10oUIC7+saL/mzKTGCybksvipOJN4Yu4IbPtl7sG/ePqM4fjAV+AEqJf9STST29H
Y8HRy2IKgrViZguYj/E7p4pf7rraVebCzNMWPjdJPo1fXKGW1OPGRrTmp/TTlh49R4DBkBSyB7go
LEk3a3Dwvg2vzZh6h1r8n8ET2nlgMXPDasOXd0DAfBic3dkqZqBA9Xc0Vj3sckdzD9RLkc4jgJmq
Bklv2In2nr7cE/SLYoMKwRAtzyCBUTiKEyXU3woYq/quEVzPgNhg4Por+WWkySBGeKU1iL3XP75B
71iVxRDZbMao9d/xjqdj3ak/Pel0OZnsOUhXYG1LGvEvWrVq1s87H9m4zHLDimEws4IpAjHJTlHx
3UGh6KBZlCVJUh7QifiOolQEZgWY1HnFpz8G98Q1aBIpCTzLzbEEgWbYnnayI+sGRhn99KxTEKt1
YHc0ZSyB3TtkkOs+P4fgdhdn+HHlg+aXzfqiBteu0d8nX12ZANQMYphJQSJrfYlALt79sMsEaovK
XFyxipvxpiPZINuRkTr1f6UcnY7Uif89Obv1FGuaCWosNm5cbyoL4Xg868eKFzqge6i0G2Krysy1
uyOQNsIJ8rttF4IaY5SsJsccZwo3uLX9AV7Lk/atVtBlSXTApzWTY1Gpo7b8dAddWu6Z59tUbWHo
NpbSj3O9Yk8B7e/q156wFVujnb2LWDbDo7IphlZar2NTy3EeCml6bMBhqONCXZ7r0RBg/bekVmvD
4cgFUvjivRYTRlXAi8I5p/ahp/8pqcHC5P1w4jYfJ2jmFrmpjglh4ISjZch6ofOpWcmouZf7eUwx
JCmOC8PEAWDIct5HuaMaFxHTESHoYKyWUToBT+GwDDEeEg/0XX3Lu8CVo33M+DmM5tYXymvUqrPH
u/uwjrMP8aYd3+8y35GOAW4FqFn+WJDQThIH07/aA1K+u55KIueIc5zBJ9R41SBFgLJSA00FmTbK
wK+ka14dcCukxyEdtbhiUdo8RUbmGgkaMRUGNEi1gX5MoVKoJipSx++HCW7H7laT5hc74wZk1LRn
cVqLC/lrerHQaZi2eJXnr84OgO+3c6jfnFS1q/JtF7CfFuFsdxWveVuDlvd1fYE2kF4/jKmIP7NF
03yn864DRknJkqbT8PnjsB4oGyvPgNJNA8q2WmtZ/Vy3kisnp47/kcK3WUK4qIoWfT2PrDHknKD3
AGebeD4jXcKog0h29lfGRBIp0Dh9+K6EoVgjRj5bJBs3m6zD5apynuDmXK57Bjzpa8d4ywKGG2HS
o9UYXMoIDx82s7dJtu+g/XR5jkD3uH2FKNGTLwB0TcExt9H6Eys/liCPQVMAD0nMs+nvcGinu0Fo
mq9X3pPUT9qRDaUMg0bAMAvrNVqds16FlxYdTjlX6RLaLB70G/JqlTAV982O22MQRuUtv4u5fOwK
1EPD1ZbFYplMU5cCExGCHeJnrf78VhJs68ei/SpOSof+CXBjbms9RVvNgtg34TIb0277rfDaZ7vw
cIRr7SkLS0XirrvzZxioDHCKWMPIMw0chb6dIMlyeDLX5WlJUVqwprbM85jU5e/GGP5fkWI3VRip
STUwlNceVn1DblOGhBl61zFcW5MXG2O53acO4nHmQR6OZGqhTTwkMwqkRm3rkTdjBV+Wdin8s4me
c9GGMJh7UJob+xch1K4E66KLtRDQ+xKPWZmybFY6SZDC9FzsdEPnkPydzZ6DAO+dPnGoAyjyZUsd
sDQ337Qm/RxP/8393D9psfnJRaJ2XSXmmdD40Z3YIctdGzjvWV+NUXQUqQygPNO4hzqxQ60ANDWq
wXjjPXXLadeJ4Sq+I1u2J6jpz046EnK0ROWfpbDQbQgET96ha+alDhTkvBqbCCf6QdNdGPjRycz9
cHSO6unZSGxrLSuWp1V9RYI6e2nU4Q0Qv3g8VwKYkIQRotnetMCKaq/2UhdYWm+bNCj5Y6oeu+BL
0dPzO0T1VKg/FQb721fVUJ5xK8diKNksVMSZEzaXEqxTmKeCNupCxfG8x4Umxxgfm9dTe0970fTL
Zy2mVekWzaOchKXwtH8agWCmz9Z58FsTqxtaPwzF403DMX5mr0nAcILc6O2AcR2FjQ/2e9iy34Ko
a7EN8it/EWJbm5JBI1HcYycmfTFv8Z2Vkb1t3pqbkzrTxSwBcN6+welqPMB9WYUX9f7j2OVCZIlp
q4C41C8TKDVlTIZAuaQDano6YKDiPl2CtPmpNbC4/Kn9L5t+1V0PkoAoGE64zjIdZ0j0y97smpZs
IHDcrYs9EbeeUo4jcxXoEuuEYk135aXNWmAsAv8fG+JjcyWmP66oB+4+C8G+oSADuad+EpKMTd/D
NrTpA97Xvdq2clBnGS4avtwhaYg5jQXvKEE3B8RIOGm1zLU/VFxxUyq/KFW2rU6337GgUYMey+Ok
w5Ip9D+zNsSneoJkkNlK8C8zDbTraXGSYBCS60T8K/Bif3xG2djHhFy8TuNyTBueKqcNcj4Xe6LX
tP6YsVIoBl+ENJ/ivMrHIwKTs9783slSSNKul+KkWa+opmsobslVyl7GlnSIiu0RomxebA6CMTu6
MUCZK/axwjFOCyEbPCGqXOQEuKJyA86bK24FPdQ5udunmqG1Zrtfu1ZeafpClEfzVVhZ+T41gD4w
jqAoVcbgG6VBGRSIxgILW5kN2zzNpNRIMD09UxWwPV2epgSH/Cgmod4OsB+isgYKd53ZtP6NQIph
1hn4EqQ/2rN/V+dI2SubSycGwvzEL/Lcja/vxxxeENqNfO/3VwgSJs4U7DmOZ6QpVl3bVPgZU9xt
uXWn5N8pJRhWelVvkXVGSy0XGTnUVkwb0UoBx+TyKLMJ3CromMVGV3bqJfJW5oNnzhq7CAqqFBxA
ExxnQ7+wqA8AdnwJdpKqN0Xzjk1ROiZm3bD2Ipvo08X5dnI56tMJisR9KmSCQc49/HeOpynlGurY
wQffPbBCAOpsaApfOSxfxxAYYFdjcvnHZwxLCqqqpwUqpBEeQ5bB6/6Ye5g/0NhBWnqDqmWeREHr
UOaD5JWCWJXNw9aVGt8eYyqRYEEcJCdsQnSMO/diG8BdDg4SLIETE1/yZMVk8pbUgDCQzC+aEqB2
W02jTZmmuWWc9kD+rPj1TW/tiWOX9NfCH4SNW9NMAD/pNDLMdzupxkqMwN+GvfG/23nt3PXb/RV5
d5HWpF3ayENECPZf+Pf+NPPdzL8mQzGdAYeye5n01Vg9lcDNz8xrJbDmBr3tzDZ8/EC4iVoyzmFU
k8QvNaR3nKlcP/UbalLXeKAG2e6V1AQwb8H3rET/ip9XsNxcpBC2on0ipQ8Mp7XwWeg3wEjHCfNg
ZULNbLvc5w6D531DVPE9VHOoWq70B1oHxwuAWuO5AYoOtj9xR7m4WW0jtu2+F4L4rNxmNjNEpZTt
Qd8yj4Qr93MW4cP8qXUou93Lp5wsY+9LAP8GbFlM3oZQqC8VLFeznWZNFbWC9VLc8a9P0AQcEghl
daTnnh/fyNQCzRVN9cfW/zBAI+4I9EYoxthI+q38d91Kf7we2eU00M2EOVVtGEuHQwk7LTMwyCiu
yrZorKal8j+vpYs/GZ/YkvugCGT9XQixKP3oXk0EllieFO3UPugWk9/wPJkDOmSSTWXZCHmp4VYd
6tnN1x4P+PaG5qlJ7f7hALZdlONLueU3i+iykamWfpo+bul3f1zOP2TMVzNXdjEODI/RIQC+PQMK
QYid7sOZC6t3QW8GE6+XS29XzBykMzK6eQQp40bq+8g4rRZBRqzYx8YbW9YsCUFnRJFfuHz05X8m
iF4hQPQY5HbWQZPeqCwswkMn+xqAtCD522f8RqFWzxyiKvrEnaNxVatSQd8jB5MKXG/k/bu614YH
PBj0CTdsoZQqI1SQzHVFPMtzzXazRJrEr2/ZQCX5/S4Ek6cw4zOqUUe8pKa4tooPwqV4Us5+1fTA
GG7AUhw4p2+kdW91860DSX/02cE3TYh7Tj7rqF+ARShVzLrmEJwZSvRaPoygK9YfDcOxpV4BVmP3
5H2vaV59+iIRpNM0Snmd3tstOvMpvwkgAaYfAGzIBzc2zWRTYUWgH2pMjEixEVTGK7yDE0znAwRS
i0m8eUh9X6KU6pTogo+9fCNllXafiY5nl3xDt1mM/PuUiRJURVcG8TB5T7UXoyCgsNlmkBhwvYuh
wc+WtX51Qd2It/z8tvKsKitS8gXxbQR+RMIz8zfBabWWgEf0XIiOCaO2rvlG3gfM6rz3f0M232U8
pPUKAXiPF3vZjkseAsFlZCJzLXOo3QojZe87YiCMTdDdITssr54POhuANSb8/i+kyaHnUGQ3IHA/
1or2AZ/G0LQxlX0hks0R7XlQhKI+bFuD6y2aVFE061K+z+TnPpVGCOPJCefEHfN1zzh7Dnw62lpV
eKYcL9R663qhqadfXUaYNpyYIcT6dKNYGzB4KHA4MGNNoUQqJQ/zPLQtl4ioYb/wksSz4vuObKo/
/92Kp5+bXZnadhZLYS+ju8U+QW/gLZTVtJMu2KHYWO2AFNHOCsbGKv09HD0YMUEDrGceMVMxW3iu
HInIyvzUrLqZqF8fCi/s7bZHkOLOl6LqP7LLndmZcSKX++ikP3YQqovRd2tw4UaVWLVDSRIsRH0H
XLQeRDytTJlIYP5CMhdFpZSmER3mzRjYWZzWV6GIaf1QEppcPLZ92X1qcySzkCQAlUURoltXK+vo
weWOwqWGe3YuFYzsHGObUP/jJNi4zMWgHG8PEqVOGCIZlyDfuIlMPTIvBF1MJBzTGA4TIWo/R3Qx
Xk1eD7sSROeB8WUNYb9VRsFql9+l3DwSWnvNKl66+TxlVm4CotmZP6PehRmG/a6zqVURFSrDEj+X
FtD2rzMTLJ+vmVzO83u1IdBiGdRgAh+TLunbi2Rh1PP37iJqAmwlCt789DZaVaQv/0atSttSeaKE
XsBiztpnDxk3IoAj4d4r3lXQ8ilgpN2oTvehpOGx5EggiO4E27a/YSS2fNVi1MIHEqdCFil36qRx
p06KLtWDEaV+a4B1Algwakf0imhWDFXM5L7oMInf3f/jYmOc8YOcQvN6RcihVkHNbDYNdVEySOBO
mUz6wipQmeI0oLRt/SDLUDPirW09rgTBdJmNSmOIWwz5Ki/bP5UqCwy7B3j3sJoaAWoTjv22CCTD
MeZqorKbrbQ6K+RsPOpsy9ryC3nA/qQ2IaxsHUWkGOssVUZGs6MeqoYeMx7fJDxFSqbMVPCSOfmt
QUhdJRkwuhpcHki5LTkR28kYsr0BHYOYCGjk2d0YAEB+hQPBWyii8Uad9jZJyuVD9ygHtXidmV2l
TN4LydSfFl7GTCAKyycTXxqt6gpaCBdJgUsuj6P8l6IX+dpI9vSwEWg5wAFAUB/W93jFrj9eJFK3
UjCwLrncdvTaFxdfH4ucmJSKbEJUp2cVYssFVwTeJpR7RzXWQy1K4/W/b/E+YYQg9qHJJJMgns5J
DcuLMcEiQhYNcck+yUviDR2LCtmJmFfFi8IDLYRozxnTHU55BZQ+gyJnWXmAl4y7B4SWDNW8TMrd
gPeTKt3kve+IPHGOc8i2ude2jZ4fdjlebNbCYCV4J7ktYhmNARXEdK/pU8bXW1iWhbD3OYC4aD1u
0ZdakcfQFodTqSKUewWvbvl3wY2SF14VGgTGiP2bbNwQmC12keEqgm7sf6YaW88aMVxFk47F/wmQ
V5TdizWAR23EocZuc8JfifFsVVVpb+5SzCetBwI5su7gACiCZROS2w5LPOb09DL9CLD2t9cWkFyl
nj1rnxHKNHxam3NUkmBk38wg9KyTyy86pEIYI+VeeMxE8TIqJarjn3g0siwYQdJqA351+6hfxV0A
5muifkilU5igPObKrzGV30C53FrOfjSONspsAdhw9bgKnkCJoW6U2N8jWkx3wLa2IHvbMaYCq3qJ
du+VJNPwy6yLHYrqIRpzkWr5iLMjR5veTYpTcLX4dyuGunxtfsb8t5miGFjQceVYNBZauh7vSgnk
a7kEGoWzcG+tWoQwnmYv4znFB3rYvg0VtUn0PQggwzhs1mpfSiLGYSWJZWtXe3NjEA7YGudhWnIe
IGl6b2ttoInsWZmqoGTUSM36N8T7xd68KqySBovv/P8j16hQnLAclEWAtF07zwTs7H5Nz7H/Nyqv
qxb1kVIJ+5rECtyJQA1nGWssUZk0RzWJsIEFzEMglgL/vtiukbHcfl0ZqDRRHUrwp+juBs5h6lyf
oZK2UA8lsHJjwae9JX4Ea5AiZsarjxlu/Zl0bK5SA2yp+eHW2NKGrJWPi/A9bdvKrb6yEMouoJgy
EdrfIR+zr9yKa+jc+0QTbQ0l/ylqequ18daM6X962l2yhHQmJAQaEaKvgXmMtRcx0efQbPA3Oc+B
5K07EPeioTyWXztIuXKrSzU5lVNvGXYdQczpepYPpIhEn9nXb2+aBNhNQJpNtQ8cKnbnNfAm5HNQ
7c4vtmkYkLxpBixToDVY6Rl2W9LRRUkNeR3wB7pPEOZlfX12mRnh14zk1nYl+rMzJy35rG9ohu2m
OolxpZvc8+6yOuKmwHfcTtb3seR+R+L9C2qcyfEDgI26hEgPuPRrE47NZR8Td562PHv+uvBGc+7o
/Vs9xW0ajBTdIP4xOav7aAuVIWPLecKEAr5EjBNk1Ds3G6V9Lgq5sUHhkvehDM/gnG8cUyo2Jhwq
9AYx2BtJYzh8ZqWyDD0Fjm+ir4qZXBYHmhQhj+MRw2qU6E/Y7j8uXOdo2MmISoyQhJrekqJnk6sh
nRhVxcp7vHndkKWFVYH/+32peXFtk8EpeWZmmCBtVwEsa4pmioAST9QrR+T8nbjLjhrSikSQhJQW
fosu+YJZS7cppSJcmyiOmGhsfGsaXbPpZidkvlbLNTxe7KZm3w3zjV1f25MLUJLGS+jJgiDUU6hF
yPef4jprfbXVusPRyMeaqL5wG7KHEIbse80KrV86X+pNvE7YVwh+X5ZbUbmtQizMByKD7zUA6Sjb
5uo6+iexo5WcoYKd1lrwriM6qeC3QGzLpGFtTVMoZAXwLn0hjhswRd4JlVFq0ZoJYyKILtQ9IPEo
par2HEWSg2FVajJfBuak5tmCXonBiaEQmkhBSE3eZr0fN83fL+obMEouzCFmzc4GQknaUnUqbqFO
jQJM/mDbdh6NAxiDScK+/rod755w5XhQO7v5Wq+WgD4IwIHF4DYKH5Vpu8tlmx9NXhuVdxBg1puZ
fYNOkKlIZugoYKspopACpWB8mwDOGdu2oe7dzwz0kyH/8PA5CgmMCZc7PQ0MYK+/XzGHsE9bPOLk
Ctcc10fym3vcyWpWts5lSPulT1K1j/2QxiZIIt2qW95Hr0G6IB/byJGiG/QT7Tk+g5LbH/8cqe9V
0CN4WKdSfChvwDh88zBWB/B7BxTRQ4v7nL7pyBp+RmRkgz0fUa6ndaqJNu+zHtEtAguvqqktVIhx
h1pF4VN25YNPZinARi26XElMN/7coUBmhLjxIJomA2DhFr4N0kxAGaP3YFVwb4NHs6IELxDERe5x
ptrqBtCn0EDOCLMXtI5iHHgtKwF2laCJXoE/YhaTekDmK55Vt7KaGSgcOl4sjYOb9d5YjGLzk44n
Wzq24a1Mho3MewHO5wEgWBW7GydtM7ctTOq2rW5wmjw40VMG1doXnyGSMXOydi5ETefxVIJAVBjf
FFtca2MAy8ZCctpxw5Ap6YkeRcYRot+YGkg3bUCyWCo9eUFL5MpxTScKzV/YTcnnQU5cVcakYSWc
4AoRwU3TKfUloAcSpFyfx3+qoV7rcwis+i2AmMHySc7ONyF7IQP87L8T0Il34r7Mq83OpJ/rLW+e
aBiHwYnc8yj1ZnKcco1HcFmHKQZStJQ/CbaECGA4LjdoVW7CvZF8OWWyuqxZMrVhF1hK9rMGYCxD
2mrqweOfql/9H8wHuwu7pVSzVzrDqOGdpe6YgCEIAm2Cud1LG0YAGWaFYy+OBmHqOnuP9wjxCRpw
GKzGSpvpTw/fa/SR/Fxva+VclFeH23xgxAlhGVicd+gwFZSDDN/8uxjPcgEceFVDkuXUHfHr/6iH
HQEvkLnIpGJka0ZFMA54LbWZ1mrqhQJFhT1LsYlXepxR4sG3adOFMLQ0oMD28SRg04JNGd2Gp902
H/L2KAf9lHDKGgPD3UlfhGd+wC2VlB6EuurX3dKo9YO5VQoC0beUC/6qnvqwWDAb0cGK6eKsrCqa
PWXbGbtm1qXE7SFwY4biJE4HndC4w5QZhIGKY2K/84M3+RMhq1DrG4lK7/FvK6izLwlR1BMaouWd
6CcofpDuxIXHfXVpSxj+KG5Ar6OabTo0GpU3FT7HDqsLC+w8VelQIXyzXxM/11xdw80UP3ZMYYGf
HwYAAlmQmC2jDKih/hngPUOa/nFQIqYPWf/VjUWo6/h0bYLGRbHWnbqa2VdkXX4plepUOF4C8EuO
syelSUmGzD1khhmVZVN2WY/3PcYF6WxPiFLGA9gSsWqeMiPiFOO5vYTuLw6DKgslr3Hei4lKHDkz
7XKRatPfNOzMInmjoi5FoDE/mnKUfrUIjAsGooB8dguWnlrJdx8FO7VQLwt1l0G4VQiJ0CUrVi7/
CHdCrKLGIuMGc7QQCd/vCCQ6R74/Eqd3XxKpMVqATVOjV0qNPbN/ijYgMB5LbJQ9mJBvWSq4uGEJ
nabo4Z4Na0XewX+WsAI69w0Lo7jUuRpp4zGqOQqJYVzz61La1+gRNntmg/9tEba5IT6pJ6hpjGrw
XPY250mSBthdOPpWvO7VyonUVzn54Lv7QiZIF/oxryOKjGI626jsDntL5B3K/NH4sOzvrw0K8bfA
w0JhPsdln3TUp3ZilmL98VBZXTPQBEQPQ9bjAeZtQW42b9tpixfNvwQSzUgIn8cHS1xBIdMbWpGd
7cDZv9swFOpFoXjp58w6fuv5r22nww6/dIu0m9VVHeN2RCXGYZyX6H+aEl+iAqobdPTmsereQNhE
I+tiGe4g2Zpv3f5A7NniXbUxrttLGspsd0QbYWVrF5TW6/SkaMQIcLY2P5E+fzw8/H7yJMWGPK/u
HtKCnyVKpoCv78I8LECsNjmqsBg6gCn+VPmHfCp7Vu9/rQkspwhHpqehi2OmfvJuKghvn3HsbD2w
The0xXWjaPc05T8+2zOyHzkkm6DOYyC369nhpQyMXjOMQeZAJC4DKqcoNznzK7wQoJ3P4uzxpR6R
vZo7300n28D2GWnJrbITh8/FO/qdlsNka7/zG7lI48F3/2s29TjOeGG6BHcbEo0L3zSw6epGEvCq
uTmhb1y7F/S59dK/y88ch3xvrkomFH1moaS+oM0fqn5NoUYDtsKjxiQ4OU6a+7veUhoTUWSGxCpb
He325480pqtUVyB1Q3havrbUr6NlHv6ZdbOnh/6hlyVYyMM0Zjoe47lnj6ELY8l4HZ4/RH1hgsxg
90pz1ugPnHL5C9+OFyVYTccBBcX6o/dgS086z0OizkojATCPLqN8dGwojv8LvLcOyeiUgXbgbfjf
3cqQBfBcbgdYMFQuYYqImGmlxPDTtpNW79ICWH8sS14BEC3D53QblGOwDJuIUZZd/oTCeggtDq8y
CzjMhYmtHn3DiVNQysV8WX2sbkdYHvRCf0luz56E+u4K0MtGzSJwKNeWfwbTtKIvUaGZRLOHeeWO
y26XJvXAvFanrb0JhL0JNdHyRGeyxdW/Mp3j1ibOfA4RNdlJlC4qj+cTzMYgzeBLF9uUTr6z95Fg
pYfBXAo5E9LUpS9U5EWsX1FEoawgiOQV2flBt1V1EanKB/JFbjkrz8rdwly7JC8cao5+g4CZ/3vD
cyrFHz6K066n6uoXyxBYyWXxfk5TkOaWFZPLzTBqNAvJXLGwPeHkA9Wydp0KebRmB6MK35WdKsUB
1Z7kmqjePNoG3rCcaBIFz+ye7RvhN4lajEfwZQMWn+PkgI+bDPDnj1Q1nfTOk6JeBlbUG+FLgdgg
bqvqKhpQwpWnyelZ+b7t2lbGHC+jY4xdfLzBM1UreVBRSWX9Vo78n75WHDnR+T43gpxm4tZ1W8Kf
hf9uoeAg8HpJLR1qNnl481h4F62dHQOSvxeVzC8nRVOoH8iFO/mnMYWJIp1p8aWpOd1rtbaHa8sz
klJdu9vSnH5iypBS7RDM+fD5ULGRjzyEdtXS3Sob8BPWvIsOhQJfqNhvX1Tpw1DHHJ1zAaauzqt9
MR7hdYNfnoOGlepNQ6MWItJLUtOfL31q/wg8OvArDIP7d63ll35qCLeOwNjdUUeysZJh/Z+XbCxn
UsEfGrqX8z5pySUu6AjH4FaBNs7yj1C4P6TiYhZ7cuDit/KOggBt83wF3YmlpsYh1auGR2UvjR8D
vlxAa8vR5DZXghgzfJ732SXOWhjpLaY4GgdoPr5iTObSmheetUrAwpoTrYDS/eGYwdsOEqc4eXW2
rbsRIRbcpi2u4CdaJu5G8UP3FhcIuWx4M88+BOnNQLNoF1n+M8cWOskCfhzv6/RRaa6cbjQtX7Te
vjkW86W/C94FSLf1Vp9JZmMh/M/1yJSOXVatrHJmartE79JiNoLqLqdUiHlzwlc5ZOfqYxU2JKRt
Z3JsH48tee8CXiPPsjteayhjWo7ZmaxfGZEb53k4XqVOfmDG3LhiLLHzKzwLW6HWEnwEfchQK6zz
kXze/7nyB4LhCS0JchByU+IU7T2ODbc9p8RIMjHbVm5cYYQjQgKpV/4vyC5Yuu3x7u64FehuRCZS
SmW81VL7djpUWwJb20oY6fM8X13USHbT9KrvYBpwqbAbz6HyfZZj1MpY71hr//Ki5JhaXblezDfJ
oVq7uWJI9Rwpzg/0EBDysY7p+a5RfOMqC91H7tZJ9j6qX+k9TV4fJSV7rp5OviPvTWSV0JUsgIBe
DhuHlvlqk7Qp4dF0zknMhEU1Lk9PNviM93Habt5Jkd+u8Id7SBGxeZn3HapzEiFv2VKKuf6G5AJQ
jKdZ6oRGHL6i9i+brQJU7D3NGGrNnCAHg0w9XPtE4v9Zz9hGpg5B/UTktasI+u6MMFFu8GVBsV/n
eM1YHEHhiopYjzrZyY6geYG3GqbC7hdXtXKY7J17X2ptD+PUSPvk6tjrCqhAC3dMqf85K7VR+HjM
ovObgVJLLnjYPptRCa7wybwkvuAEfKdnyTXLdHiP7amK9rPqpxkkm34YfdRy9AwA4RTC3hXpRKZA
T4xuIPr3BvoLTxJmMbh5cAIWRdTaVSDsfC7wzgYsWujVp5IhcNnxbbAzEqqGLLpJwEZPfOD0SyJv
km7WoZhR3AMteAmHZvGXkIPNH5mu58tsTduqo5kQmEJE0ozVtWRf8T6MbbrsHLeNjdycq5+NQIri
2/aIwBeq+T0SSigBIKkrPa1/V1HAjI6pbWb8m9q+O/8/seKAPDgNvqukabwybc9iJLtwiHXskr7w
OzvThlIDFZlzRAbPI0eKdVr9y3fPWgGeg/iDdop6SmzCkBuRHljxZzP2wdhk4fO4p34qC64OB38a
NneYRPU6/qbXyN0naHWWfjTgog+4iIkdmZ7WlL1dc80YERgn/QWEv+yewRZySIiTLP/1JG8NQUJe
XPJ6OMVb9kIPuBfQ7m05+Dp5Al8l4CGPsvUrjVK8zXcIpi2RHCLTcJRAc3asLluYnl20VBNjsPCR
HtVucGsi8zPdZ3I+4Bc3ybJWT9p2ihbCAf9ZgRmZW/ANFcA94mhBxRwMWQ42jrj56djm9OoZTt6A
tD+7x96YoW4zWml0FEhnzUOchsvQixH/GZs/r2U2Wketo7Fd72EkFYki2JFmH8PoG7TsffD7JlQo
AGJto1mDQFMv9snvyKZ4pTLQigKNgVohekWswU3PACF5/WbQBueDHCv+lFcqeaONlSt3wTi+shHD
Jvh/Al7S1p1y66uav8OYVmPvBtu1phHonERhYgPUkU+mpO1f7SoRJksUb5O+w/8sYruGIU9g4yJG
elujyF+VawOKPlr0S60f/vEB7ZgbJwV/rOKNmK8aG+OWFwxjU4mi8i6L5sxYWNTh525FjxEJ3ops
MiVplYhAo9t5ifP0OLbR5efeLW78F0InD2CKv2fnhCI1BGb78bSM72qkjs3zNAsfILf1QALDq0jG
XhTVw7muaNnCGRUu9lNcSGDK/Ocftm7jd8bLyPPUwvZWnb/oOMe/DxEDrmjk0aqzsEO1702umMyg
uLoL8B5SsZK+bKIQzFbI836mdMzyCLtoqEXdxacgS6jZWSC0h5K7y+1r7b94P+kGAUB40TL/Dkpz
67cF9XQLYYTyeMoggka8Zgw5vCXcYClfDpTbc/WDA5c+miH2VYksSy9+Nxk2Jvb6AS9byAbI38w4
vefFSQ6A3vR5Zt2UJNMyUssez/K1hC5W58FIlQmIt9g2ixb9jZ3inj9GpOmGJ93DnPhHjl32mPmY
Ex6RvfC7/E/HpHYNsJP2bj1sXXAh9kT/2YrdhbjbyPa8kxiq7qUZzgTEDy3dP6wcxZtCqXSxxI3Q
79agehlJcYIED9Nsq/jzswfByixwnNuxMdGP++21zqpiyKlPuvUP8ScXSNds2FPl1BXTDd3AeXtX
013INSlvtXSTctdA9P5xiluRD0KvM2fFoT7PGle1sJzghgll0j9lJufVevMUBsURg9Tzb/uoLS/1
mmtS2AE+01jnXvqz2RDH9PttaDYoCIDrRMePnVwX/2ocT9k5X2cgKucaDF9uBhQwLYJrxl8ByJDG
w1SpwSTOrDVyj9bFRZEYhHtX4SPbBnpKxknV7LXv+alkXqzx9spzvo7gV+MMUHs4TLcYCnA1D/CU
PJXbsba5gQhzuVL0szdcjYAeoZQDtDqd3/zG8fhvgAzzoFbKLMfUXmlKnL3r8ddhuH2MewtY4Rod
AM1qT0SZkZ9UYoEe59gWNRzuo/APsoYkw3xCZ6N3aePpsp18yD1RR82yN1v6XN4R7WYaYckpJ2kc
2dPNhDiwi7hJQanC+O7GYIb1BdOkNJhz7fsfFil6+Xjdw1Sc7agJSK5feIQqbbrN/nv7Z+SN62Lk
xri612r3Aamc9ibqCmVAdDSPZm0nEebkbpla9tqhqfc+GHQc4Thb/cddMP1TtfQPAZUSaapj75s/
NW+vyDku9gEVgoYCvYeIM0/HbzG1LhOBwUbkQmukzNGPHLSOaBzF+eBUQ5s+3tD5AZs3aStvKPWa
Foyl48J/bVF+QCq3WZRZyrlG+rNJhoFlIms02HGyx093AV05rezXEuaFESqdw7nV9HjMrliYXuvi
7rMpFoTKSC5inyJSoxBL5WAIbf98LywxQtUfNKxOi05qzzKbQfPqAXYthcmECYmxdgljQ1DVR5ie
YYpFq7UD15BL0bibNjEwVYiu2j19XCshL/45TIUDDjZVneZpYtilb/wE+7OOI1NWBkjS86+NnQXR
D/b2OF26ljRxJoZ1GtmhgeiSoIKxT1Ku+HPBPrNGQNlHSjTOaEd8x5vqK6YzRx8F/d8CmHTlNP+W
dVw4CQ0VqivHwNIkPtmRqddOPe3W5vAVSO91wb+PD2XXuKeXNz9VNq9q8b+FqORN/MtpiZFtNPXc
+b+TUCPoLx2PFJI3rDIdAy+ek2J6oKwZdGbvhEcmPFuXrY1JMlCBV+19g5ABDBtaQ9A1jogTqDTX
hiyOADVWOZBK2ttDoSYHgtKf0zIHVStO36IpMT9b07pT2jQVfxh0N76Zw3P9HTHrjyJGCYR3oTJU
mXDVTiELZec+6Y5zlD25/fyWuY9C3hoUP7o9sAeFgrzOXBSYRpCnh8v+Ut29t28LcAUMHZhfhTEt
SH2pXKqMZUn/ijz1UJ6RC60LxCugJPjmbEwWbJZoQmXnmoxopV7YumL0B254OrPiSPaHcQSE5xEO
/TINj6i9BRGEktk5U/2OKtOgIQjLHqKzC5Z02+bqLMTErLP56MR4uJWRNC18PKBAOl7mrnD1TA0l
yDgMifBOwAmxOmPDu3k1//bNEuEY1LjrfV5cs/+hUYw2OwJYriqb/TP3WDuMzxc7/nj3eDxfEAut
7PXXmCBh5ge7TmsgiUHvb2spXllvL+yKXL2F1A+iVS8OMC8STbYsdK8Ie2CILEbWxGxQA2HjaTLO
1fnZYUcn4e9t++paPSZb/CfIrVaL8ZX47lYlfd2uC3ELXG2EYA7xtTdCNsOUV/8Dhto4FNnnNdDT
IIvAn7x/II4Nr8DO5pY/Q9UweZuY44RSzRcBxnsCEzPhMNxxSbz4of/ndZNZpVWBF/HcwobTL84f
ClSyXxqZ9cylMW+uYcL33CPOIf5g+BxUPcX2CYnUTGIGhMJbWTFbIIkYfAWjYBmg06NHSiIAp6Jq
1iZ+6zXWkJO81VjRkWGRzUbBIHvBnw0bVWPVKSLKVQr3BpOSACTKKMC7idapsN/NziTSdvVCFcdG
6DWhXjQlq1qatwxihvO5JIONKJWh/kEvnvCFfyzq6KRLFPgqQumI+Wc7c0P43Dal3C4Oo19i6xB4
qg0EdYDiUT4TNf8uutWfTDnS/9nGUzMe2RcrrhK3+R29FnSCY0914KeGfGR/1lWenav9HN0DcSmt
hrEC2nMMNe2/aWMDmwmSWiAd0067hl+a4j/0OXqQjY7rBXCNFGCrJrUSEMJmEWBB7P5gg9RoB+82
wwuofxaDg+0KOBkI6TCaW2ecJW8fKR9f9A0EcsA/m2lCeKxML56f4BUBmcGlxBtxQusTO16eIcmO
wSgPBu/65GS52baeWzg9VvREnmSEcGlcE3GZhByRYga/qA+Qgnk4FFJUKBD2H9ei6Pxc+xwJi6rl
O5/3MpJJR+Md8FRLu6c+c9XX63o+h5OV0jhQqihyEYMGLhaRqq762iCa/bZpCwmc1uhnDsxcU3e5
E/JgWSnGQZhmNmSPlQhu9+86MkgxJRTWxswOQ9A6mm5nS2twlQg0GxvDDQj5X1vMOeVW5Pqtjsdm
FeFceZYCme9IZE/4iZrT4tKa2o9+0XI303kLiB8Qf9X4yW0qKf3gSMs/Aa28djUI2SyENbrN2ovM
Sf2mpBpe0kk25mYwxiV/MOen5dAxfZVgpAbdnuHmqQlWBSHnTZ3sub+Ac7FXWVfuJBTJs73Kgl2T
07pcoZAR5t342XHYGRcZUgoZi+TTQeCK2gJMnTWR+HlQvVklng+3sxg04294IAF2Unrdw2sAeVkT
/RoNwfPDqhk4Fo/Rzqv4mQd4q7czQtiFDZYEVe9fEKlHfDun3sNWUByvl6suMDSLq7iurazms4JJ
IiuabLEbOFp8B91bnH+MPEbyp1crDbX4lRg3rlXL0VKI7uYwzEnbM5MEDqvK1oDxdkOrFWkRdGn5
LCpoTxy8ZHQ8hxHbDIw7nn8HCS3vjOCwrGEmC6/IwOy8LxKQPvYSz0EGoyUmKtnmMQAEp3B0VZCr
ng3dPrMvTefPzD0aGQySVRuQXdKHKWy5OcAXB31pU69SvFYQ4zWplwlP6eFTl8o6VkddbchEWPZf
832hGuZxpg83dr21rdwU3Yp0mdUwAX8EaYW6/GSjMMEguMXqr99P04udSCcfAa4veRpN8IqQGsP1
k1lvh3OV/kPXulnqa7RsiZCHG86Bnm6kYDTBhMi4Go4a7pV047SRmREXVoMyOoZ+xIUC4Dh1o2tK
gZtV6vrQNOeIGrmHHx1FPR7eV+U/gFfZVkBR+gD4+m2RjsLab23+s9rrUPH8f+5XVwkjFxzDbZy5
9VdiP5BC5xiNt5psfZcNxdkK/8lGTxZ2CdKFLWSbibr1gaqxzg+T3ieuvH3Y9wKMrQcq62qdx+om
FlroH7I9xd9SbP840zNHwieKWbbvV4X2plmSwiTtG/2WEc+R80q9hEpaswUxLmECcV+NJ8KAUvaW
qKLW5UTOg5pSzUHI2eXgDqIwWo7vm3VgRFOOixJvp568bxKtilLUC4Y+2xpPDDV+aBC2A+tmGFjz
/b0AoCMabjilr4M4aWbZoAlNmcmE18HBO+d6Grx06jqaBbQU8fy9rg9tylmF1IXMcI7x+5a+GVPj
HT6A34QfJG057qe/3TmnMPLJuGGw+TJeYjEyeG8nyI7g1HLGNlSpWEv+EMr04UiHGqq/InAq85wb
Frim0wOUiyPFH9EjHdzxK4TSnuo/1c8a5QZE46oROFXPbUPsZIHDYdF49cw8J17Hpq7URZZ/h24U
/aOPZIFANCAVh/AfbY189JerwwyG/Gz2zr+u0GMDFQaUEtV5QoNneykTBJMz6t59P/KLzuHiMAIm
bSGiQ1kXePYycyhkJJoHDm06RsioE2ueEohlsShAJk+jo+Cg1DQN41b+L6Y/OYYOHS8ajB4X9qu0
Nqspzat3gVGQ4tg1Dxpumnp/zIg36aVr72FZBWrfRa+brZNXbq5wV48Lakpe0p+oMj+t1AFWXXOf
EgwgDp+vbyXH5m7cnofT2Ghv/hswZuYiiMCxogXRqFQP3mRQJ3OFRZRUjW6vY6IcDFZ6g6DN/n8z
fuoemHOI+38KoSlM1uhGtnQEUV9HpBITZnebIvo5q+O76eNoqpJNkFxLRw3lKTgcuUWAZXQ9U9qf
YUf4+PoCeUIYAbrmXsfQY5aZQZZ3+EhJ2FKrt0aPMmSyZfgLqP09M169Fg/l8JMzux659Jz1qVcU
UIffnk0FQVJXTp//TxTBgPiHGjQ8/kPfRtlp9QcXFiIP1JNx1p7rL5QMfbJljnh6WYt+ocBjmzWH
01WJV0K/g/YTnZLIcvE67zer4rbxiYwEt9491QtelDTGdcPPJI/lBJH/9K39DqhNemz0kZCf3gjj
qNm4mhNKoiJ2RWb97dpkaSqutJaaKDYsUuf8TstPE7kxB83bXWDA4Du5XL0MLQv5fAPgi0PDIc3s
ITiRyTovGgox1Zt3rnlolfvst94HLVsbhC2Ri7j4a92T0Z7V4pgVMGk/lZgF+E05av52DaIVAOkZ
Ysxw5b/LOyI6PmN44YeGc73wJ7r8TtAEdQw8ijTGLvQzpA7+6TFkykt8lCCWIJDXMa15N+UxbN7/
n+G8jfvmIT2mwaMzMuJeunBPykrsVoZwwK6nCEvAgGmlyaBW7d+VD5D5GcvAilZELsyezBGWAdo7
ksbbMrwwTyDRv+aNbA/nPFNmNaP6F4ryUIsp0CIpREu0IrsNJAWqNwi+3mc7btyuXqtIiHOTr28E
E0Bo8hYOa6vUce8u2eYnoyjOqTOqmvN5ZWRQ9DTfCPvx9kcnUHyth7kmh2ZeDZOmVQc7Nn3OHdrk
oz0DBCwxAqWIE7xFR6AWdgwFnz5AhJvWQHGre0L1Kkm7GTqC3JgM+hGQU5sD6yEBMxzJZH1qqFgk
WI/bMLdh6UrTC9nkY2+3lZxg3qZEDcf3EKz21vshHCwkwvJVSO4dVNoCZTe3IaVAJQDK2zBzq5fP
yh37QoDG42iTtt/tc4TMQOkbRuTxVcBO36gBMcSvHxCryv61odCI75cohUtc3ipEO1ikZwu2acwK
Yhc6xggp7P6ALwM296jXfwo8G02q8Gq0OdQ7YioVYNuYRb96j7Mb3E89278unVXnY5eyIvH8CGrr
TdummbQ+0iJPcGObOsBfonHrcoNBwRY1Hc+wIKEXa7Nh5S7pgMlfpZeEJt39I/x7a5ziO6MXUzKa
xTuKq8C0XsDJlOzX+dJEK4GckKblGYJSuII4KVYu4hIynMkdH0mlifktTVQWvo2Smzyqy5ZAsc0H
TuLPX2jhY2KafxMQtwzTX7xhysYQEXjGZr42d8YE1uvEE/IOhpCorbCjkweURtg3OF9cEDmJ7yT/
EjaJXKBDf3Bcj24vZKJJfVfDsdr8AMkO75p3jwE6ngZcK9BcOgKZ0RUIpWNMWNDKaAOnPMjmPxWy
E19UIWGPlqFLmgpE6dtBmCaYQlCmHFutvbKIsaqmfSxYjGwJhMlGYJGt5gQkyhG7TbNzffKxxcif
WrzXb22JdbC6RJdiZfvgVLrEHKZvkiQ6DegMfa7fBf/l4xIuKJZDo2zE7rGFvcSU0EPtMZ/gkYui
5hIlq1Qr4rxlJy+zHshsfdEOOTtaII8oEktHvSuiyqGd8FF1NMLt1hNC2ls78ME+xh9Z7ST5W6//
/MEeUxDenEgeW0FJ/RqepDR2VjgfOtf3g5uxCJTwY9PnSNgEMivjCYeRSIgenHJtHfNA185lq2oV
EkEb/zvKPOLsvAFLiDkab4cb9VU/eoQ5zQbdOviEZ+GL4R2iLWFo/BaRY4S9++DkhYMPrceR0Pu8
9HnkNmoCW5IX6FXEyzh0JhYdZY49v5HFAnNHRMDNBoGSG8SUQ4e3KNkaVPlDqlzXUvMWixJ0Uxe+
ZENlqya0wU3SJ1H92l0aUVrBrlCnsL2R0NK/0icUe7ICiVIjtH0slakGdJJVmVYo5YMISdc6yI4p
FEOOGn4P0M+r5RjhKh6a07Ceu3nDxM2yaukp1oQybYDhEBOJhBCDuBzwUw5Eqo1xpFkUh7bHKZBk
0+nD7ORQsvIOcviAUcT6c7fLf8yH4i3jSld5YpuwCZVeUp2gGnVffx6MCVA3C8vY1Zeeq1Rg6zyO
rctiEcXYrFWuTkXO4epgQDNJlKr/rI3A4pRLl2HNqJ/nlQyrsPwu93uo+XQd+uXS4GNhtwWaAAOl
Mq9SqhryDWP3R4uUzKv8nAfxH6K+ANUpMms77k4Xc2DlrSJv3eEcojyFPWpm0jb5hCmuhVwdLASf
DGb63p3YqXmtMJPhlfB3mLEi8LrMV2YiAWTZxzNQDz/5sRHmZ3BgJNyicSaTvXxB5IlDOETHjiIu
elAKOIiqzIEgdUjwyzqevMiaGC7H1gEU30wFMuBnTD9q7vwJMBYi1b50UhrmBfPTA3M/vbvZQ3Wg
QBdYm5yXU4rjhXvGbiLQbV2HROlQ4s4G+5LLtxxWst0sou5OuUEHIq7Lfh8MvHizhowLJXBIrRL1
yDBM4rkXQx6rCtDZId9RowF+9nxxq5RTcdcEL5XJA4u8DcFlv956M4PWX+HZVTN3NZOnI636KIFz
x8j1XbnwW0bJe1PxGJNnIIsVqjkZi5TzPZ/gLBmSrS60KcwFBj34Wkqj/aCAHWxSoLdV+E43kMLG
GDVeXPUVvgB9np8BJBc6CP17bFV+GRwEURFZPgWEmiwZkTsW+jR6NtafPNvL1BxOjZWR3BaynCa0
sFVIt3T/2E9c7qGjvwh45FL1GaCQe8TlzKfXAq8hldWH58TI9bn0UEUlg90jDEK0boGRU238AXTP
SpeOJva+vtMf3v++VxmhI1bnMBaCxNRFjYWmKPe6zi6b+6Q1W3OZ/elV9+3IdAqeEmXiyHcPlmb4
AXUukA0RrAwceCmVVFF5UVqKpZ2F7X7JvC3blvlp5P2Xo+jyAFyNNNMCvNym5JbbrR8k7XleW2io
H3FXeOC2OZZfB5Kuko9UQAtH0/+b3NDT40IE5AfMlwCNeJA8b4bjZqoIdzXueNOmV68F+/2t/euf
jCSz8t0UdY/LdSXwnbgSW/h/NHhohu0g6p2kMWKoAsxSYZ+dTiNgWy5qNu87mMp4Os7/kSi+7uCq
yY0ByjeTllGewqYhjLXbpjIuesb2y3jD0nRFkwa9JHrbPfCXQINxMvQ6/Ct6FC+vm9TMNVjwZaAC
iPKZqb4Rm8r0QcgeefomO/j/WluE3Y2sE9y1E/5o3/EEhvSGSYSS6E2dFOaQ6mx3QWK4WgvnZOPi
Jm6DCMOZj6HHi6ngYzoEovmzqOQGYCZ7IE9+I1/c1FKhLHvpF1qJWxNbWRKjv0bmJZ5/HRi5JYsp
PiyvxqSQyajX6YP8soRC/rpcslhgmlLT4DD5sfxbJZPyiXzW9z68kKFPjRRiqFI0X3XMaG6Wg82p
ns2YDBOIu1Std9HfapDYiuAoQQwu/XHLFSqfNwAlYZZ6T1ACJTWQReimd69EdOBI8gIqXvfYfLwd
bEnftJrQZmCy3+0im7EQTKlDjW/mlJRBfCPeDxsxzI/BFHNeLO2DqkvG6MJ8Y2c7/omJTtWdB13D
i9PBTzT4RqYVJccYI9i8CcZ7r6wDPx4P6XlpGrAhPMDErFx+XpNyPgLCJ1pvRBaQdOV6IdqYnXEw
NWfEMJmWFwIwEeCBIkQg7PchNNE9mD+UF0eA+IiTk5s1gvNRqfxH4IuRmmdpH9+4R5B8POMeuQ6I
Mk9n6JRtWGmkzGXaeWPaRgZmXafBG6SSlddZ/wKPms3TAg+RTsxG6TrVYjbM4LBbIDZjNAgn2HA0
uyBcExBU1v1O7YKAEfME9gG90HBprerHx6ms3qwfrajm9aCWCPIzF3pR4VnhY+9u7Wz86oa2aUV6
W5fVvMhvzfR4T9gOhIPkoU7YL9N8Qikw4l6ChL0SKIL1E8sgmxh4nfUbZJQH9RliZXt0A+V8KAjE
Ag+2Me8r2IAjVOYgIX8jCQBLVObChKjnAE9daP2ZIsVROmAO2jnLzlldJ1vI4CA0jNfMSdI+jySX
A7WWlDeslXN47NhIJsEopKVr4GlSYjcfYrRDHuvxsqbK04cSgEKkkeQjK8fpJuwltBmDQCPfRL2K
mVTs59IT+koNXGntUaNHeykgkMaGyeOjZS8NxPkpZQWjDgdgRr2IsZ0QQEv6xztqSeGNNwzFDW/L
aQjK6Mv4QUTCdDYV6Y2fBi6a2ySkrWpHRjBOMEiN9mmef+R/CVz8NupJ/4/p1chNHGIsyupwMLv9
hJaRbEr8xz1iaL61xOvr0kX8x/6rsDyh7BePGLk8hoYY47XqO7iPUGAEgsQSVOQ4Xm+RkiYPfj2y
BjFNTFqT3pYgZDjZSfNMQq9hfRMBTdaYkbhC6jSleOdktE6dSmNIAW71AI8d15/7wn4owfnrS5YO
SIPovV+MYJEIurL+9J0Pe8Yq42KK4Xh2dYqk02mZJZDHFc8NvcHsVxmmx2/7ETN9NGMew1d2jaIL
idq/QyMv2Y1gPjcKWM9cZtRd1Yj92tyPjVmvKfHN6qm5m5pfUaJ+MBFroBYWuEyZewXtu5MSoP9D
o9OEqVtU8Q0ppI6MHNDqBqE3GNIngSj8wd8XH7vUB2anOFxqxyekHgdPJDQ5pc+IhCA/v5XtrY2l
eomcF1yHBDotpZG+Hwhu5D2fX3I7iLbZekuW/k6dBLWYKFvy2YMg0QirWiJrT+5FsSDwTmss0T9W
WykhG9TBaVJ3y3eWKXB3334GiEyXqyPFoKGbRui9I/JPzTYG/SOa8SiTyE+gsTMfWKOqg+RED+PM
anRiJiy6YZnxFmjcF+fPD5d4B1HwdsWEHy03aAgUfdTpMuQekjN2P/SErRbb8p37I4U0F4yRNXxj
d7m8dMuNTItiwo1R2IcMT2KZnnGkU8w+sPsmofTvSj1JDxj1GFiS4fDs+MiIkjsw25h1J9EqP+3e
l9wdXPqfEMX+CyZSeHfc++/vaPyAI2xBP+nkqUclsZCQY+6skmxpFPNrja102jIqPqA4KgeMcBIs
K2ZOlUgh3HMENUTBmLdnJtuVid+9qZhDF0sOQZpfHKsxZ17YkRZPZER2YTB7FOmBDRUzYhfa0+71
zNm3mmx12q5wwPui31QYy5JMx+RPugyLnpa/vGPLuf93LaEw3CckUhl0Fy/eCA5K/eVN1kaV7dxs
d8DRdsHNw16t3cgtRkGbH2UaeTBMS3gWAt6E+reJwtnHfXerQ1O04XNvr69bTayS5YmDmgXWLsoa
42x/ejY4KxTQUjk+a+deL+H09HYKEs/rlmDmi8fZZMU5FC+3lmm2NRcbrB612l4dcrK/sq6Fd0MS
Iu3+TK6pBk9qoM+loDVV+928n/t62qH8CxNdsFvYpEgJHZ7xjl5Dc/SiCd8REe3vOPT8p9Ats6OC
9Q3qd9axy1mwLiu4ELvrLO84i1pH8VnM4ifSoL9+kFfueMKxGXMpDd45r3Pt9C08wJ3TAoGC3gif
s8lCOdGPahctohWzbQ56yUTWm1hLmww/CSQxS0GpaZB3qDSqEUUbeC5steuEagEgKL3eW2RohEQM
FS0oByr07uVZGPzimSp+XExlg/Bcznt5ctSx6bTBNJUaD/noTo2cECi/vZfmRx3mfdPgUNvDMOnT
QzOt+UuE3K9x6D5kOQsC0gcvZOHqmTcWu5CLy3WI3Pk//2tfmROXZxRQACl3fiYxuWtXivr9aw55
kC8iEJ0NXKvPieQkTRYgvd3xCeGDj53UklXQB+pUCq8yJCf020JiQAF4cVPfsV+RwJ+mLh/58lWk
eZBCMcdtJ4+/A2kABEJas+Dzmw03LVMzjaiUiLG0dmWIfKnbTvwByQQ6Q99pEpixb5KGGtX/aPjO
HyV2TK130XceQ1kX46HPgb1+CFfUGIBznJbJWTypQ0necQGXlKdOeEkncj3SICA8IrnuTK60smq1
L/DfRuPUa800FENfHF9rQlLp6KByk1XSFZ/f29ttqhpBOFXCs/FWqyRY6AShJtW2clrDdEilQEpr
anoGJEpUevJxkcDOEzqJAJpx8ujQtgicnripftzUh+fPjp8qhhZIlntWlbNxTEemF4NqArXhwXWv
MiQHzNzzXsN4kBMB4mJfrQfh0OLkSdOzZ5Ouz0iFZVqoZe63wQU7JuoX8lNwMS1tP77RI576ZtPi
ZES0AS5+yPwufJ+yfIPflKkmtgz5z2oLCc7YmpsokWUnOFR5U1CBPHWcPDj1pXm/kaSDBTIpQu3G
htZ/J51+J367+lzcilCFSo4RK2KMY1cyeKKIYYiRpYBMI0dRVDjOfvRN86KHbWUsivaCoiWNVlC7
Ppnzcl9j+qkrQKyIV3crgjli72lwgNMPdwo8nW1MqmjFb1ewE8f0w8xomwbgCoOlq6n8pe+QZolc
brpP9BviwTpVhYKRx71ZzFWt2H6FG7vQSJqM8b1hztY3ebt8tdCY1pZq9kkq0i8vcDp8PK1K4v4J
2+NI5RlXmYDW5ZjJxN2X9e6eKK4+3Y5fz7V73IJETpZdkkKLxF1JWSSn5pITy5k7AJ6qx+lEcgn1
2fYeXeag3H3tTPZkjeOIMk4z6fGIzHdr16AzmslCHJ4e8MbBlmovNxBS4GDXeLsfPQIuSvzhb82v
ixP+6NTayoq7hFoh45Xc0PPUIagfxYKr8I+UoZtnT9j1uFgOf4SYAwoHW1D3M9byp/D0XMM5R9Ep
s1PvLSxKOneuvbDF/3xzKbpi97jS82wBGXJYEOuVN0naVIAzpR6i947s1y489k/rbuQGGmxJJDo5
PvIN9xP5C55wFlr4Z9CM0i7zrQ8xZxYsPFVPfAASW9C8k6KVzq/f2hcPuL60B6+y8/Rkq6ymhiwU
VwP/lQ5L2nrmaZOJodkhAFCWM2cMDrtt9Bhy6ZeIKKisi+zlgYLRXUr5nTLZa0iVsQWy1H4op5MQ
dUNMWCqZWvzMw3ar02vMPlwIHQbW7AchmCU4DBwK8ZAv9IfD5Ran76fKKqv8UTUM4c1rGL57pX4D
/cgVwlG5hOwzzYaZhJAfQxfsa74Q4+N9OY2MIepGAkrunC4yiCQDGR5yPdY21SyId2vReTZ0Gg2g
6ycXRerpO9X1k6jv9Q0sBzKu+gST9F2refvrptdy/wELJKVbD/9mypTWAKzzOCxtxtf+rTkgRccy
0QyXtLw88+09Fx8ixk3ClRg/anZt3oZNEAOYNZRS0lHPNi8VvKR8avYZK1xQcfN3JD3yYCeHNISz
+yZ29Nnn4PfxyNw+OTgx+uPIGuh4i1J3F095AWq9Kl+wNvOVqek5b8j7NYlp0XxLRWsDyAEIiwIX
rnpqbxdSqzgqjpvLHhDToenjyAC+PMljOO2v+00c77HwqvrxNxe6PI9hieW4if5VG8Pu10QjrSot
KtHPLdRKf8dVtzs3crSbgCdKB/4EBMQfuQEZO7J4TPnYHu3lE0ckWaroq37jHCcBVp2PS8C1rJtw
c9avr/HmqdJQ6O+R7QRzbrl5KnvI9qZE2c2di745kiirofb2TQ14/K91BIbqhCj1jOax5EOihA4G
LBtdqaW2xBStSKgQqk3DVs0euJWMAAa00nXei0/fqQr1EdpPQKziKfc04OAFCyfYeiOeQWVpQ3wm
xq7cQ68jXJe9uVWTJt5TJ7u1eUNMZBuUPEM4bU56o7PofI6AwPEKc0EupJXlsVS1u144jpQ6iOZM
fVdaTKAIIj69DzA5/Os2aZ6J0QLb1iZFRFQV96CEESAw/5HcRDbDlZn+z9hW3FUBmkQAU3nAwPuQ
4h3c9lQTB41TWbS0444/6JJn3pZjfQrH1RhZvzev7o0m5a8jLUusmqmaUAAhZZi+k0PRseJih+I7
+A8r4enGSTp6IGIOlCoKT8Gvf/9rLI3XzVjuT44DTarsi++rgeCGf9lGX1El+cw+o/0mIBOb68fZ
SiKOSvo4/WDJeF7DysM6ofbu74BeSdlrDypSA6VENcTU9njkK4kcceQG63ZC4iMCOPAOU4Jjw/CS
u2LU3vdwVJk5MWZCLj0WfHQADsf9dPQbwiSE/CTUybgDeAr05FuXArMMJX0I6Ld9VWcRIKn+IMT/
AaECFP8Z5OhUqu2XPKZfeD5lTIPtnA6+uJ0kT3JQ1uReLs128kYMZif+psykfGAofDyeTIdIw5oD
qn1OEUouRYtEqvpaDz7yvYY9gfbxozMWWCeOn8RyYIEz9TdpxTwtwZ4M8iS0Ibj9Ewj5sRjER6ZU
TEc4lCgeHv8TDhALsrUWo0j17KeeYO5BAWbfESUIRE0Bu4uXEP/boudqfgjcKGAWAQrTsSwMCYfP
SIvJlilmugMmo2RYpQ1hvYNbBbvwIpy02PIzGmOLsbDsa9QQVuICCrq0jg66goEqhJ3ON1woFF+y
Sf62NjT4QrpHlIgt6bFZzH2ylO02pbCzslVWzBp+JdePnvBT09/AvgVCNZEecKbtN73vbPegrlt+
U3XIm4/98IW4gkfGKUhBK7U+qxn2/H0njpbyVMSQgRtkbrYDFYL2R0GUWmwa1EcdwU8Ewmikim80
gqxWCAG+DY+jviPcKZR+06U0WlSic1rpGpRT3i1h6lc6IHIPmpXJ3Pgh56e2kF2JEXb0e+Sb1XmH
WZhmeFSpezWE/KzCesLdNvpu/q7iVuIgEsIvN4ampXSVL5PMNGCohBvdXVQCrDn2HwuYhFrvB4W8
FG/8CnJd6163qjfZjGL+mfm8d8Z7vc6c5Vil37+wlSc/3uLK3jbmiIQh6/uxWDBWv2PK8Kim5P/2
45GVbJiwzDqEyKBoBagFzCmuZ/Z4zJwBfsFpyd0gsXUYOof6f0Y1ZDlL9uM5ngzZ7f02g5m2SGPS
FFnI67jbAuxGbFlUdcG1FV+b3eix1FKctsN5FZjOePyeWfFNOZZMZpaW2yvB8WCiub9LKgCqeL3J
KL9oFJ4xk/Q6nMxP6/KiTIXQCwtQrvsx4Yotradus5WxlDkQ0+kiHc4RkAmRlRmRHl0OdyZVXkzK
F+cxZvCSX/7VLwsQ7CjjPtSI+pASHy1PB6MvMT5Gf5gHKIjgu+YS5FhjpV4ZoPzMuqRdxCR6HF89
hMpUBjOhT63KtIfbtz33YZYGc3tto+5hN/0uAtBSeIZvupcEcS69lUjyeLQQGSKtH/kRh1h8SSe9
U/p+jnwqJjTDnIT+3ApWb7ayBA0du50swELN8/1AyHBUM/2ZpxOfWsCNKfvo0fFIp1a2VE9hFBXQ
Fxds0XUt8dBKl5pOpI1ui0eZlPWBUMj0o11Z/QA4/0DwuWyvkkSAzFG2rMWIPKCkl92iHF9uFCSl
OYQVbEkEVNlPw4PqhIhEh1chkwZBS6HZqOv3fYUaS47oHbcgzW/sZqwa/O4ng5PqhdKBdRL9IOhv
fdv0oHI/3UwInlS6G+wxwdmlfVJqyHlFtMFC51gSqZin7g8TggdRistPMg3bg3SvVk3voSlJ7Xlg
v+DH/f0bVAiMBiefMExIjunIgDvurdVFOrh1w/bb0CUtxv9HD4/MOLELpuMp9b+xS9zyqPTH1b9x
G/PnaiQXWbQRNmknG8yNBMVvJRexsBprJu1jMiauvg0N74OHnPuOT+oD8b90MeHnSAu3RnMF/MN8
1hp6ejwRBRmVK9ohjCXXktVCixUTsd0SDulUZWEKSlT4o7xbtgLV/RlDOlzLFzDjMGoVe8e5vZzw
XTLjq7XoghGR+6xlUaXCVN2IhWPUPdNz47+nkJhksmp7UPJxQ+FqVc/xGBdITWShZQW48RRBdQHS
QOeUm2AM5uwlu2QleOTAewdfXGwDbAUZqmrh3CzG8QVv6PBKzN8isOUlDzRK7YeAZzHTpXHNqtj2
PX1GcBG5tNfPplRx8efkTKK9r6+hLcXvNVPjNhVE6d9ge/syt2/6L6n7ELCIdmm8HGerDVu2F8d6
NEhIRPh9b5US18NFOo0Blk5W4PJ/qXBOzxQkFOfp1rLx8iy2hfCCKXzbQxDlZLmmzH6OUfyr+hr7
A0mNUwVeYs7ZoEPk8cQ2LzJI+0+A1nD9kp3iZfl3PUzkeLB5Nw3dFfCcBTotIjhOhxg7XD2l/Fvp
Bj5/V/NL6OHTKdXjUWvBA87eB2/l8YKmSLtOTP9Bw5RZfN+EU4ckKXu3HIeqslQzNpwWuhGXe87I
2xw12OuL8f9rZuf9Jd1njUXwVdlrKi0pjcU/cRS1lPpPBrjMDcILNAgmneeOjnPWYj2bJ0ZFQDtB
EqsSAOQRwcwBtTAm76fRi9UwnowUZblYUBPY8JL0pQ/8aVYRVtFcKSl20uBZhZnKHuAWYEMcmimm
DQJyKfDR/tuwKLH4KR4XqT+DvXiLGTyENwWbm+Wztoq6OLwhw0/PHYiJFcdJXuyH5MDXgPXs/KYT
5DRTzH02lAjtWu9a0w8TvkMfUGO8tMXR2g7vrmTuVykj9eGws+wvwj7yubdzgyNpnOtPezC3MX8w
+Caa31ia2DF6gwmo15EgyuHm0nUVlGVqgQwgqi2Qgx4O0gsrfriwgbiNbizUW9DH8rNaOohMpFKk
W3CVxgTrQQETBkrkAvSxKrqYlMJR57qXBdMtUKuo6hvJXPadTEByFhRtoUwVBEUE/SN4dnAmy+Eu
bkob2ecOFzzedQSiiiUCFCdUBUkiNENm7kuJUTPoAbrezW6GystHpSJCxr6G2sqfHcbA8DwIirMD
osH+wqCFYRs4NpmZalAufbPws/cprG9A6DxI+c4wWlfjorN9rLLerXFJIi20BgbgegVr2E0kRNBP
nokbHsuxa8y+9dpVSGE9XUVFYwTAeEqXxHN90M5jQrm+XJ2VBdfQ+9wcxw3LaH2D0We+QrecatQI
4pusojUyKRFMdJ5Xi/wvL/S3TcgD6xHiW6EqeEXnmJKPivXxPp/yjnpK6t5R3PgVzlhgLNuf2w1A
7AebFse0tU9kuWXKEEhVYHXRZc0A4AFjcJFQTjmvQIoCfe1kETTlI3425x+ur2YdNrB5bUwEmWkY
R/G6qsHLCQHpA0mxLhctJ7uhdJfSKByG4H7SD4CJKHtozeVf8bbWrw6YgZTKJH+6CbbuK9UDJXny
8a0XIkeDiGAvbZvuitAl/zcfV+RZiV85uu3WbGIY18Ng7ql1g8f62aA58PSrB490YfBw7CjiUtsr
+P4rIVMIu1MVwjZ1DPQcqI3YtphlY5pL1LnnGeuzCJhl9rg7QtRLcrwmDn7x8mTCHNyc6+ynr80I
HJkq053YwysyrQmzimfAgU5OXxdTwnOFwVTBBItq03LHa/okcxtWAfLQzTVh14CquYlmd8/hjawX
IjmYm1mQ1eK0vt2tY6s1xIpRkvpmO2rBPbAZEYiy4isTRcFgSfLnAaJPMy142s2Ri0h+uzAKBC0E
f+G66fHHVLJOA6vGE2su8HteiBG3y0wacazLFGRVg4eKQ0qoPsXVO/RLrCIxaFc7kSe6e4rpbie2
6e/YdQ5PcMecLLy4nOqkb5YpFcHiWFDMY398Uxs/Wg8wgVsVPke0mY/BzoEYMosufG/8F9cWoZJa
MGKy58DXCWTzZH3IUcjZ81E7pCqCu0oFm3HKWRNsEmJGnm1/CsomeyktariESpvS2yMPA08kL9k/
/8Z/hJKol7jc9QPJndbk2neqeTwNMR5diVt8v0L9rgmZp9LLAVVpYFXBHAXBKZyvbi7g7u9p0gRj
NcFx1r/116mMPpREzLttwv8M0e89jBcikLunDggF4lreszxLjiBMyDklVCOORaRiyBbdmd8IoZ1E
Mh2Ut4j8cdmBoiXNYvGmk9AoWSsyt8Km0RQbqvSRea5kt5Ke08OSbtIUYzCvi3T7L96jp8BBsaac
mx8B6EqbyhoW6cGQhLSeIzY+veNV0h1gLrxNhDmIDijp8w6NpUqXwNbxqt85+V0vQ343gIP9JYWj
1A6Ci+3ys2PCrsxXWOhicwX2GFDEXiUz+a4iFzDAjaodybRnV5piLkjJL2Wlf3LSKItMQZ7s7HTc
RH3lSP5k7tW54xGWj0+Hcgc8SAsIZXizkkGgcTnBBD5eg+JMKu/TCp2O03gUzszg4HVKjuSnaaMg
vAoUJslyMVmNIbi/Clh33fjt66ZJJKEATnYkkOdKHtTg25nqe9U49py8lfle0zAH94ISlTmZ3MG/
9tyobwBQGxczyL+h0fEMN5yCRBnelb1Cd+d9232qg2NSgl945qaFwbSkSQw4W27DiiwbhYh/hLoJ
K7m2fFvk06/mMpsG6fXN6NyPN4oGVLOm/EbcaHbXyOMA4sy3MscGs8GcY8KrBFHE+TH5Co5p2Ub1
QYz+z5zXKNIp7TVvHPJHEcq26sEFcKuPvAEKewwB6OK9JEiLainr1CeAsge7AjjPU9VI4TDfutBg
PqXlRtqvzpFvclA7RhZaNMtKTcYnJ7hMEhZSTwwpx6ncFqgJwtPJTqygl/3qQZcc/a6cZ8gzwKCm
3gAwIcKxibjpUOZCNvob2j9CbZnC1/HKre9a1E8YdnmygrZwTO3SU0jiD4+oAzn9D0pr559+GBKo
ti8oWbrsd9jD9/ShzvyTcHYJ2OdGC3HTBWtws90qsq+G66rZXd1YYwkbWw0rb4pxPqjG3mwo0j7Y
RbXlB9sGyAABaAw/qcEsd0AeHXcLvzTccxz7d72zPw9yeSnOf0MFohTWmVlIeGNhSmJL+JZ5qNBG
A5a8d1V0ZgsKYQEpwh/RuSaq8YrtR2tPnzAZ/36H/BI4AyHxX8rPjm61Ncbk3BD22wbUoXNqUyuD
W0Sks0D8Rgmh4cAI2hX6yk1KX6Ccwm8QhFFny4RL3h6T124RVSUKmju47xEOyou5AW7MbjSmsDHA
2V1Ni63pQDG5t+3xp1KLFLf4GoTGohhzfbISWeiQfz001srtFFJdku3X6/NnCFytWNmJCJXYNKsh
4hf1d347fv9vrxfIVZdPLDlZaWHbovm1l2muDWsOSNG5AdNOVgmUXWA5hK+rWT4kFMkBl7Srbq3u
9fPKoK5GGj3H0m4oTQCU1JtdLpXAfQy2sjMwJQ4fJjkY9AwY1/hiYDvlZTP1yNw31RkrwUMYAfzM
cwdHuK0CwqbSKic9YeDztvVHfwdWysOxc0EgstZ85TlQ4eHQW/cpgtdSbdvrnWdMJJzM02IH6o1f
wvmKw4E6+sbFdKNbgjdZYhRSJ0y47PCNHTQSyrfsoveoluTJpd26mP8YIvXpSuh989tPO9Bz8rCw
C26MTan/YRQ8kXpN+9VOP/RksYYI2BQF2ZdPAxyVUNKWuDPBq9VuNeMzUT6fwtqDsQuCLiO5Hd55
SN9bAGj3kskyua6nksVujutiaIPdfpnakhNb4AezYDGprsczapkVbiyUwNF1A5CH1X56W/n/8CFH
wet47znWslpL4lFIhKWfXJ0+bxaDxWSmnTPxAMUxaINEqbrBtrIVG+rRB+KAKZKOvE80lQ/ASoUK
VtiCn6Mr4JwNJwhLVm2ituZFxhi/rNljC82g2sray5YXO5UAxxzKyNhyFYixTF5j7g9Jg2FjJnfG
oGM66cP8n3vr9R/5mIldGbtg6rzOusLSAFvT1NSeRLoIUOcvn8M8YaLfHK6qdULwKBxxoF/qHPqO
MuILdCzw9kXOyRbW5A0Vlpn7HrY6SNUyUCUF3sbtIn+vW2vOK2R2fRbDV9s8w4bSz3363dJRSIQS
b9XpUhihHaFiqWk1IwIyqxErYRZcOzM9Ikz6LoCJya9WeGxH0KeVQIwjo8cn5XQVJxbQeXOdclTp
306T8zcvS+CXrE7eNU5Pe9U2ME3ZLcmRtBOeAzjAAvFxDpj5kzZxb8lEgW7g44XhioLR4oJTWi/K
7P6kCPfnflnocPjLfU8A7cmDEuCzxw2WbgcGCfjgQ8xf1Lrh6OTz2rTPrjZKzxn9Sg0vriIjw+jT
QUt5psYRxKQtspgVsjm+nEDbWl+87VM/8Vbjuh+7ruJ0mJ2b4chAqg1dv18hH9AhCQPHRszDhYlR
3NCF8Id4ayuYfjj8ifp5Hllz0fTOFDE++2PFuRitN4j895GqB8FkCxd4wHISD34RYpC36XU97YAv
bvKP+mTLDvCucIYbpVsY1KuFiIrlcsrufIgV5nGs3usF0J/EU864IAJ5Q2iFf5OL8uMJXPwsX1SD
aAs85o5ndWqiXzRb7DbZC43gpNiemvMlrkS2l30tKJ7YzdQDeaXxUt8HoMsORU4+KpnFHyhU9dq8
rmF1TCy5ptzKLVPSKMsobB6OBcXCOmA3xQiNSZ5Ekur/3B9Gtwx0+leBJlNWb0hCe032/osB6F4F
j8MoWqGKIMqwEwt7cp/X3h7R8UO6KgC01KofN/wh2kZCDN28BX6AuZu+77cOSSOeAdtf3dhfl/X8
piz3cyfeTn929VPzrXia0Mw5ttQRnaa89Ez2VzAY/F411/6regUfoSiBUSoM6rhcBxx3Ij5MR+cn
xcIw3xJYlfLf5x60yLv/X8V5tAQcfvrSwjYF+mEdrL25ljjmrq/1WMykJutierLBJDapFzVHsRtD
/ZtYRGwzsLJX46BNn1qQJJq5vazW2fakNnThfj3BJGkJ6h0bzBkCay8dysmdCd14W44wO3Hp7IU1
/SkYFF1nJdaooE0TsD3a8zDIRiPupI6Kr/HQm07bzVqwL3+37Nq9oMRzhrnrrZVVvNT6UrdPBR3f
ryB1r+dDBKihFxGE2Tl6GbhxzzixE7KDcYVPtHUEsWOrfOhiG+3HLbh9/l4RNQ5RFd7i6EaztiQh
nt+H41APXWyOJxlHjV9Tser0HATTZbyTMFKnhSsJyq/0HGVe5uBQnhnxBS/CFph5hiFetsY31YrE
ky4pRLBD8bFdJRooRmHNI6g7raDY1I4Cfls7sUqKCQwNm1JEP4HrGm4LkyK4L7dkiEwyNsF4gkzB
L/5+PaPYJCClPmknFWNuMeDjxUz0P1heRSzeAlSnoaZzkcaOJL5Zd1rL3AHd8dvBfRA/nKT6gD4l
0Wt37riMysZoNSzzffd73Zk+11DBraIEt6gJXyYP3k4oCRtj08YxBD2TyFmme+0qsZWFf4Ox27Ry
4Rr6D0XnTiw2Ptr5WQ31Pz27PkAiIzuTbDzedw52Ze/y1M5o49AYX60sVO8W5myl/uKE53dWMUZ8
7nRy8ujhbSFi4cQJRlRhMjHS4n3HTWoGuEifrThW2H0qAALqoR3CAKiMiIjoJTvCWiRcoYSK9plu
qojntR6tCQJm8Z9Q3OtuyhipJxA2btywG0TtTrCgqbevorNiBn1yj23t9fX2p63b50Yt2NlEWyEy
PXjWp9BhXXEXZymvbI93GbxwQIHyVArdgznkQUQna6AJgA16AIx1yDAia1oy+/+RJ01XqZKRlBSg
PsGnPTDaXICZYC0v+hzugUFykDhCu4ioAmj3U90CBZ2sOUnhAoSUPRY6K66u5EH+KvgTJlE8Nts/
NJl4gmZQwGubCReDuTEDCuJyf06WTSwyqfYrmYw5gwyAZAoo6dBb/Nntu1/K5rQATgwYW/y3J90/
k8eaVViMr3xO1HAM6MlT68WugcRxAXrKI0Go0qtT8QisGC39wYKs0xRhipIRNFhONPXQL/ChvXAO
M1qo+NCEWQ1B1b1/ViZlZYin5ohzcRkiZXRZZbOPas0yyn2fuubR1YqlxIR6M8O7h8/vB9PXkMpS
AUAhGiTB6WDh6CuLLlhDzMH6QBp9+zloUQitQWST//vPuEGU7bsaaWoKSYpoavx4aW2fGh/EL6TX
VC49+s+FAUaCoEyrlZSCwlWMLf7MHXb+reSYtc7fBWTe3cqZqiaBfNl0nDyGLfXvrQR+EgsJeldv
SfPr0sMrFlHthiEGS/zOTmtC5WVWMWKO4ShhJHNjqUyN/d4a5QMwu0D2+iAN3rkDKh57oWFqKFC3
lE3WpNjNIgJrgBF3BPgrE3GLobo8D2ufLESiAm1cn0ajTu/GS40JxUtFcQG6b3asDMqPSPJKl7dR
IWFxAFImdcC99Aaej5JfMWnYuUCsq774sCbjLi8VTbf69Gm1gMsmLlNPGdQOvydUl/yHxvqsqXTr
9ZgCnTS2BhU8gIN0FTKrRXqat8Gku6E0GJa3RWjW3n/qGPUUyJgPC6baTUo9h//dN3NFCFbD/OAm
UIp3jaEtld9jEzof+LUxRFNgQM9imSEeMxnpTAgjjeVxn9D3Dm2fdoJlNAwSqeGSvgSvLeE2MEVW
ZwzHxC1BZ9GY4XncO17z8eX0ZEUHtg1Y8Dy1TmSRM0mkUf6f0lYvRPzO+hDhPAmFeJ/3CMfCJBiV
laG/20eLauh47OjNQCidSbkZnqZkPB3dattet7aUvxoUqWILijlC/aho3Un2OwjMkBzK6b8mPSKI
45MkygGXvBoS2yKkMSB471FWq4vhlmtCn6CEZAMCRceNOGV1aYsPqMPIc7Z50EsH1IxTUsNf4GbU
IK7W0PVeN3iTTVC8dEB34cGTez1ttoXDDwZYQVB7uCEvVW/ASUDBCozLUCPn3ETItFyEAoZpiTs0
7zj0U2+SOsiOi6GGRNg0+ac2U2X9hLIs2cApOg72G6/qx/j1xScQlf+bI4LZn1RpXXFSn/9lmkER
Ep1MM6nmRwVA8YI8+xfVD3IpiTobOjVgYgQtqwSKwEUKE5FO0g+ncN1lFxSLaeC64nJWPsG8dO/H
9aLf7WaH0YHfQPfli3ZvlJ8dtK2B/hIs1JF2oGbHmeSMr8c63PJF5Q2kirfoNSuMs3prPSVd0IiS
nCfwRhP5k001XeqCNQn941+Qwm+TgfYgaCtRoNKB3aXRWSwTEKco+BL0IkWIW6Yf15T/i+5dvXqY
umuMjPlIu4zJ2q2NW1gfW20ZQgYB0lhPx3NJ+LLPS6fG94Pd4xnw6INjK4N008hkd+rgq4s8UpyA
5aey56Uovx3tJSlIToouAXP4icoTy2oVZXzBKmwMBCfK3Cwc8srv1yv3P6kEAgNINdZcKxVZRcMJ
PIZSsmEAnIP0tc78y4AtRbM+3AjXWfuTE+yQtCFsAGGk0MU2ozNeNi9yvldRrnZ1w/NWPq7CkhOR
oqrUBtIuNgwkhidp/yeqlNmhi+DI1eJ28Gq7q7Y7zzfzLXG6YQV+ny41Dvepw/URcaBrpolcRxiv
B1BrMs8efIAEaEhMXfNF+WlUlXorhbZiK7mRUwiwrR+TcgO5JxEGTOR4LrNXjQ5AhX0aznEb4vVI
g/biJwGZdfs3ZHcKKymbkwU4L2iomf4cJx/Es3QkEouUyXQOswyBh0RfeubmPym7nh4q/OB8RSLa
9xUs9aIrXihWeV8i2bHOC73Gx88zMYD4BJLRZ1Y5ELDD6z4zlLKzversUx+i/Q1ULYqCYEb1yCk4
xU8PBfC+UaAX1JkqZNjawrJhbM+LNTd4lHbcm8syVlhfZVCMtCniyNFzmxFiPjUGumATWUeIQDMG
ITFBYaQXZBaD1N+DSBZWyKWFu+Ui37osVDSydM97M5kUXcGq2fd4cj+mzZeididhQ2RaRSXgfxxC
g4AYGg9yg5A6bOAyCVWGoYZdaAfEB9a2rOI2e25vrnZlibJNdDNgfgDu1TEJn11LPyJJh3/hksAA
4LOuWgMNCDBAKRNzcQlazJI1fNg80ibN3CAy89dIWQnFStJf4jlvyS3kHrOQqdN/1ZeubeAwuHur
J1bYBiFd6R9rKOZJwq0BFt0lXCko380uzJ8Ih43jKISTukTjbsSFJIYT4/m9S2HLaiq7rtFph2BW
yqtLAPH8LgdubSubuZ49/Wcq++qAW1gGeMwHZozL71MLK7YX+O7JhZaX2UJhs9MSPzR+4f22GuXw
uEwYRNOSJY9/beA+7Kvx4vu1JUyKzur/FO4lFHthJxzEFCPw00huzizDZBW8h47Ke2ZntlDMySvn
lPgtvwOxKE7yNNH1zzNORtCK3LR/qeaocoPpIuJwK0whJgjyVWlUMWWif505zrDxZOZ6hVn6qpF0
f+N9KZJ5lZ8Hc793UagVLJ53//hehHecjgZvaK868ZOMoS0ucVnubev9B+zT1I2vmiVX4w7hWntR
Uqq1aNuFRu+Jt1tu2eUHDhDrKQTVUL6xOBhMfnluraovduelD4RRaPgcjKMdZ2lKdp9SPbZifwWW
pXfHjbFFfYaQIIpvzZdef6t2DnQxazIFjm90XnjTJH07WhuX7vAOi/2lzFHstye2QHHWyKmuimi0
CTOsAqFRDIZNZE22cwayKh5Eqe5/C+hjIcjRpRHNLVgzckkimT2lXC3f/2dPin6vNtLZwKAWn8rA
DxNsti3e1KO2rV9J/5k+XG5WxXv3Gsuqlvwo4rejQCd7wtde8O4k15/TSjmORaV/HqnMZrQpVWED
uHAcqw3JSxD6GGDH/QYGSsNvBaW4O9CyRRROxquDOThpV/A+RPfkb72UU4UbObtuws8MhiTdakg1
HbP5sgs626QcXkjCQsljLG7W7Sso1hmeRZeYGmX9fhc/CwuM9CT8WSBXCvMjfoEZ2lq23hUevilS
SIy6CUg3LZLmC5DzcBEJ/E7Ucm05n1c1XoE+rCSSOc7lkUaacy3X6ldlXhKbgK9yxO3mjYFnyFAJ
KCcGzfkGZq2j5CkToyh5uB/Cmv4LIxsUKwl9kf0tcUsidb0Ei8vqGa9S6PM4z4pmRu5boWlAt51A
izQrSmBnEQK+YEaRi4GgdQ5DEsp5IcrdOSLL7BzIfWiqxNF8zhaM5Ba1c+z830OGMrMJwtTgF096
8SGJk+VDbTYE0rc0Q45SSihBXKfjGk/1bQ03Cu4UdUU5WTiQHc3OhZ9ZXN23iZRQ+WK+QrqXUFXO
7wLY64/hMJ0HI/en7+xowAPKi7M72g03NLshqfvyad8RB8b7pq1o8rwEN2sbWnpRLO1/bWGY/dqJ
CVQB0Eyy4FOf4O2RkCFh2GYCFNmj34WblJ2p1CmrDslgICVOqGQ9dJP5YfQ6TMoVzuAGBWnAXfkW
Y1PlkNi1b+2+o7c+NHeX3YkK73Ayj0H492uHcWwK6XaZKVbvwHyFxbxm0F7k+9D9cv55AS55iq0V
TqnxwekYHFp1GqY+7G66OaOfUifH/HnqM1oOq2Jz0T7C6taWflx6i9rZG4IKl7lEx3IKErkvrdaq
hGRWDk5S+/0vAN2Ef1AY9AiB4C3IgrvPBV0mjVtVQi2lAuDga/msS0j7vM142tNcqGd/aCFxRiuP
6AQF3AQUIaaUU3A7Fpp6t0cwRFviYs2ODu/APVy0L3wFWj/o/Ba5jgFe/d5/MY7Jn8Ndb9BQRuVH
ZTK1H+wv4ayI6Tm6UK6RFQPeK8tldRiZuXqOXTMGtZ08HF2RcfmPDqQbhSG/ULftKN8r7Y6Fy8Ps
srJEJGXPgtGL0+/99O0QdJI+FpJenkNMJkWzJRNdKEjTtyOd6LVzi6MHwNmXlz/HNAJZGXdXhZ3P
FutNy5CWqJ64NBX05KI0MUOlYcfdkhTlQvNtXlw8Yjn28bOnR9DIJi5vFEmEHYhACseLdCfbJJJD
75UeHSDGrVI5SYiyp7K9DVJPEI76WprQtnKJ5WoM+mmZ6qP0exbmOT8KoHM7zOKBgNz/h4CPRybE
HOh2sDIB6uKv2g1cey2rDuYt97g0w9Y8xWTdT9jum+DWn3Rp2vO19QElno4NTnoTJ8X8AJWy83+u
Mi+e3LOOAL5A8CMdkNGhkFb9Bgb3SyXTyxe4MiPLTvFRcW2wpktM4Ye0EIWAxA97hlxau5Jo01ih
aCAndcRMMhN+m45aO0FGm++klMQUzDKYKuPWxsS4AyVj8qEDdNMsqvUyjLT6at/ZnzZQNIuCYhnd
6Ipzl17n2c04p7mOxpeNpLvZZdLMRVxxEbgeo4AVHkehRTL/DMFNSdS9dwJEl3BCQTANyGw27cUi
fRuHtCpPMktPxnK/7B4onfRSWSVKhte5N8Lx9s8Y6XYABvLVUQBH/5L7Dh751yMyQG66G5oDeu2o
/2Yp2KHpDHykvzOkvpC1MHbYa+jNYACJNG4VyERLfn9EqmLy8ZxqFT+XTjPnwnmL08Ygr0jku+zJ
45h3mVI4qgmGPZSkbsU5U2gAlvpaL4/9N8OIhiTUzklzPL6vBwcQ6O56myN2PFhl9pYvmvIlhvvO
jhWNUX37EVWa0Q2yCyHGFkOMa1FXVRSjH8xIU7kUZnRszDT70yY86nnjHx6pY3hSJKK8MxI9mig+
OIM9XSs3ISaB90R457l/JZASe2APkp8eDY7ZTeNkoIEKw1knRQiLLyOM+wV9FDFyDhO4/HkIa540
RaDNSazZMkeO1myr+KDWfP1I1slLjmhhE9W6S8kkid5JFLzvOudVlp1T0m9ie6kjiMIUb3b2Ep+h
dkQNbtssyksQsk4UGKjj0pTT7YsJAIDQaxNw3HG6pMBoZRMIyeFcluu4KLE6rBJ5Z6wqt9uOnnde
1k9m1jisdqhzn1xjbGGE9m4fsriGzqe7yX6gooPHscuIZJirjTXPlPlktolfOUKPI23SdbZoBzl7
F1i8I95yZZTESpe+jL80YsrHxDBxKalIzXYuRSgoC63i0LQgDJwjurDEbC9Iz7a9D6uhNU3ApDF/
ruhVvbzu5XmkUP0/QMiDJfWLGry5G2E+cNq+C0KYWXjxl8BrPiT3vthr0wbt6cLUeNlq+IC0HPY2
4q3TgPQlxahJOOxeKA99j/F3UvwGsDysThulfFZyKQfgpNSkHOuVCRvfz0VYAnk0E6NMPaRu00PZ
HC6Bs8JRqQfilxZzDcipmzeALLcZjXDMQ1499qLUZlJktkPfCdcJrpR9HjZWpH4D7C4f/rRfPzsq
Ywj65FRuFdiLDoJAzk6Axm+ALO4LL6xZeEJrqytPse1dWBqPje74PJk/fDVjBlYdpYWwTIVBLnQV
Ghr4IQFXry2TY2Jxs9//HNtf/Sk3yuNajCZLtTjkj4xQKRAsteu5670kV4T4Vk/zOMnaJWEZArhC
DiflQ0H5TXTt3V4pAW6Do5E+BcYq1i4ac+EqVqe+HGfMMFPT1JOrMbsdyI6f6PT7d9rDItoY/Tg+
OrYyu2lhJA2daasE7N4uKTc7gTATvP+VoriYuAUmnsYvi7eQl1niykkKJuyuSqRnhF7Sn2ySdNDh
XO7fbJkR5vYQmWLePFaFt7XoFwQ7ZCCW2NI6M9QNmd4oEjwvwegKHGLqEKXedO6+1M1rKfPWBuMM
KM1sV5tovTOBJeR9AA3iWIHOfr91NbwrNNGjNTZ0NatNyO1RPAwUNpIBdIMpj2yuYH3OSVU0ewZ+
Sn0w4aPnxCVG7EdIIw7KMC1eODvcsGIV46MdgyzL3SEj/ui8lfGJpP3l5yWWRkGaa1Im7u+Vx4qH
8M6dakQymLXDYjvbnJoA7DLb0VTktI4NjiPTTYsZJ7yCJ1Wi06PX7OyUUXYNEsO7qJ3olxldzXwl
iFWO2QuzGoebwA2Y4Tj4NRy/q2nRQBy+lTbmplmjIw8ymj71VJPm7Hm42Zx4ERZv9kRARmPsA44Q
sUwkD+pL9LxsILmZbKP/8vrlV758rDKOzyiu/YWezd5PBpoWrzKLYgwGj4CicgrJLyQcb91099DK
tip8PfS8RPTC4gx6c8D3VznL9zrnyAgBfyTYS5lFAXchzTX7jBKnkIxIJp1zVndHQ/zuvzvp3RrD
CxC2p6YDSjeOHlNKn862ANgZaG9DVZx2k/cE9y1LGYzECj7fRidNdN6SfxHw3ueT1gBWZknpIqua
gJorhHNdFR2XBbrVJpz2sC3U/7P3MQAHM08vHcqDwEAhvQRTwLMIBOHVoNAnZHUz44XrdHJCiVCw
kl8NghhNNVI3m/5FllHL5ovdRzYqX65dHefIJFvuXqlm7Y6F1Qj8GqLyDtbdW/oBpOM2iwiJwUtc
eSMFqaM5iA2Ih8ppIXzh6qBXf5ZGde8A4bzcq7aqYWrBGxcoLWAG6ni3dBuDBCO5yRCxKOiupNcu
7fS6LhGguABcEiaTE1TTW1spAOSYVUhIyZySk/mqlAT0zID7kBtACbLb8ioRPGjA/3Pzhw5oB4lI
ERcDsIBgmmzoBljqbb2g+wQhrJ8gXgJD5JPElmh82FslBlwiQH4+hx+OIYrmu88lEEaV+dzi3V2w
qLl60zcUgQ52geJZwgjBjoyf7rYrfunpAxjQNJ0rqyk9+5akkLnHPPS+g8ZkhWqeO+ynpsmHHEw/
vtxRDmuYB5YiTH905oPDkTa2PmOdrWME24ds63zK+22Nft8pQm6+cv+T9Idu0hxkecDGmWilB7WV
CCLTP2Jdu239zDRCn5cYI6GmUm41X1zQ0bMayHXbv18iy7UX5EymjAoskCwfjyRwe5Pg2BvpQVUk
Ke5lZ66UdrMRHQsGqd3g92ZWzbX1QlY11RO0YRIyyeCLKHI/6t1JRI2Hjm26peQPPmOCXCRPJ1JY
gW001fzC4extuhI61ucLIKqXMbk57SKfrwGQ+x0PryRB+spJK7ZKknu5sdVOoKjt54sAxVvkKsIc
C7x3b0H/5PU4z4hUs5RDinZPkjImq8dzFjpE43rn40Ic6WQXgIXWfeNVobrjFzbQAnOsVvaewRE9
+L3pzTif0cDko/lEDd6x5iVhjQuDssupCcgx9ayE2lAnI9CPqeYdRIusX+u/U/c7+6FqMjvd7PTg
Gja6vWu0Jdo5XWkIaPi6iSb/hW/voNyWC6UHtRYS0yw9vwmmzXkO7y7rkEu6sgxrVLr7zTwjNsSd
5B9dPL6jixwYCdC72p8xQP2AhGLzYFGphTPJDbQnyN2FzafdJ69nGfGwJG86PHyJAkih6XIsgZi9
JqU/Q0VlyqV4T34YfOfQ5nMwvxhoeohWU0FJdQTEKO5uqsO0cwzfqr0IX+Iyknp/ycZYYJMLL6qk
Ndr+uF/4y+rd+B5vxrye1WMFptRIXga8qP3ycDKBOppK97iGEAv87VC9xqsKE1RiwFfKVW9kD00G
h/YH4I8uJiblXybsdKxslips5XGKjR0Zxa/gs1FEjSmcv0ToA39AK0/XDVSDTG4Hv4yRc6IxBO+v
zIO7NLutULXmUzVpxTuAxRYwLoM3Nn5yR0RRww1oKi56RcmVCj99l2s9uz34JGXqiRN6xqHU9Y22
3trm/yYpAwEwuKZcDa4VV0MdZMonawuOlNjiJ3Tdyp6UlfEWAvsJX8agFBNQFa01aplCQE6yO+Ra
FPZIA7yZMZKDcCU7ZCBRzj9xpbFpD4O7Ts2GyLAjrR+XY1ju1olLOl0aJtBltMxk2OSTdAoXihhL
ZUTwLMkPfvyYh6Ox6ZGzF443oXZRYWBrWzglDjhFKAp/MwQDI03nISZGxUisqkaPbNIpN/i5Ztgy
MxH7TcOtwG8pCJOXYWXgRmkb9Y5hyY8PCXFb2YC0GPvtLN9s1eNDbLpFUzY4rb+H+kCkVTG+Bjdd
r4VYTmjRL+YmXi/jSrPDJ0hme4II6LPfLmwTZGArXxL6pHM+6URjMaIrx4IzKf03q76RszYTsfFb
KaJdQha7/935Uq0onKqYvaQIhOJXepoBFWVXZsMRyYX+Pqk6KNFABk5Mtejcr0ed2XKT0R+XzTbB
tUcvNtkcbj55njTZhEiCkmJKmmeYTsiD2V7CUxDFnrEP08dJfxwkTIyO/FKMHgsGI/gNEqHiIQNZ
IB6lLmuruWvX2+3b0TpSJncJle3080c5DgImYonhAUkTjrmF6d2Wl+GCDlqCyXQS1wbMGb3sUPjr
0WyKR5CqnEn4Hf5iBn0KybTNXnGV1A1BHEOKV1IBbS30vYAcZ/ZGKSFf5ZylXbPGyfT5bFNwudWr
JejjKl2akBFhrRvW/leY11Zabtf3gYqu89K57jnFcBxK6GKUN8CjZrGtGwzpIptPxltzPT0qVcye
KtD3E7NrkcoDVpUGqTXGKGPY9ArZrS4yCHXU+1hN6CFU4lLjJ3edSCWSMN6z1gCs1SW4LSSIQgg+
DslZ6KrGQyDFKChzBzvEbYs8FWqnBzrSfdwdTcr0snF29UgK9LDyo1Pk5cy+gl9nnVDYzlS169Ql
A9+BTFDcZWe/VfsbJlyMGMxCgjiu6Hqgk6R3GzCuSoPPBrcNLJ2wy0W7QWPk0n5Va6iIFZZQQn4t
tg/BcZv3OoAfOq6FryUVcGv911wddrXTIvVDVf6g3ywcgAs2Sct4HXkBdPY34JvaCBDUDokvN0c7
q1IobweQPVzMbQTl+fBOvf3JCPpwBDWDDGnA7UhPQyit5+/+Mi6hAcRQyayZEJJgu+xq99tuweyH
6zSWHwhaF8iTYWwwoEUj3WngzJtFhsjaqRxUIrGsYH1A9v+LGDIk2NoIdJFnQHrqbpq5P1THO7Hq
FuRxIR2cXwldIrLTqRSdk71SLGO2VG/VTNv7GfLGJjDWGqHGNCB3Tl6pAa4zAMLm0yJU15gxMYYg
TlmtATq6sWmlQW/YURlwviB5xejJoT0T2QQGOGGZOmMZD5SRinCVJASTdRHgBNCf55hXcmhhSKX2
83LtVIQ/+UxnTLwcX0v1+Qzp/ZCR0Jo3L6qckNVIXU/5XO967Dqigvat05m2JoTaCc0/One4eczQ
cYk3Xgjs6WNjXAqmDFrQCVBg8UEz5XlsvpT7LJRXua8s+HbGQf0nM66dxPRuF1gAqVQ+q61gRGub
snAfmoPqi1QdtlX4whsUr+IyBh3uW3y2w05V0W9qj0ijdTDufW8obWBrehxmDL/NRp5ORlAM9wlF
H/X28oTqDfLCHt3zpaTL+gNPL1qGNXykDC9WTk58EdOv+6bs4ickxmPU99ASeaEKebE0G7NIW4Ka
NfF3PYPKI/rxMYqDYqPVSeQvKbIqOXZBuOEEesPwooOAi/GPg0vMNhhMXXtihUDbF7tdstoeWh6/
tr5miE62eVGhRKLrUNCBWYcBecgOtaekhcoddOdcUIRQ4XiAu9vv82HpftKoqoQI72DQqB7zIyds
LQfBjN9DtB2AQ/sfWGQyxWGDCV5OtgwCmJz3Z4EPkFC223uvUYG6YKWTQBriVm3eg2xo4xxZAfNX
81xdodQx30UnTVy3RR/FTLvfdwdJQGZuLjM52A0HlCAnTFQBM1fcVBaw/fM6hqBMxiGWeeswqJBA
m8PsOT7ArpJy1ruddwvQDXH3fyJBnxituhEgIXRD0udzERDCVq5UtiXsJEIQiwumUA8RT3V5uDnR
68LDgAVt6rZpAhXB3IYy1JVHGmMn1FR1Y2ZtIyKeOus/Ai2jZ5ZiQmfbMKPawJ+pd+XsIHMx7jK4
CW0fRovwDVSh4JA3oeCtmfhd8wSRUJPNLeEQR1IJPpmHGuQtILdohTwuh59mw3Bsgj8KpY8mfw8u
aHTJYgFbCQQNr/H4Jb15pNYXLb1YkijrLFMCRGYEiUXA5vGWIgRLHxY2rR4wnX6x3Xi0+QCsbBc7
sYQ/CskpgeHAmd2UCoLg94qxk5AZ4iohZc77jl+x96XNxbTlVXIyd1US2rVtKLx/BtEvCQfj1aaW
sclT7J6Q2N0XEbHer8HcNMJtJHK3JVmDIgaDuQsiz2p+1uknhAU3n+BL11W/2ehY21b7OuVB3eiS
q6DGj6DiyVLBA6LDdYdcSS+PxiABYhxibV3HmaE9ZPtUab7X/nC8vaugIpwnNzBsETDWXCGUQ5a6
2qEQNN8AEr+MSGoq00rgiETrS68Q5mJdF5qbDg2cXIDfg0pnTHGEUNqphmp1HhMrbY3CJRJHkdt9
3E0kyzoH4YrupJJK7zomU2x0aewE1V6hPg6iW/RvtB1yf2zg6rgP3R/GUCsmEUor1AfSHTD2p6/d
IpOzLzYr+Ve4EHXs+RXsBB3+jvTShmo+eTagrz9sYkDl5D8lCdVNgP/32w4fwDC3wRTpucT/2fpn
YlIPP0LR2TRHhhyqAmnEFN4oBC0JBs3jE62Rxc8OcIuiQRcXc4tXaC36nSnTMzvZLlYcEF7MMf3F
lATnsSpflOMinf9Htpf8QKimQXcAsBiE9iXveC6AcgRGV9hLDilZleylXllxzBxlVdKoeYJlpNBD
0zDgK0iyn/geDlabK58byOPdIQL3ENZAODa6W0u0GHm4n/Fbz5TJyszPf1w8/FTvJP0TqxFYUWHr
7mL7Bvdt1XXNglQNgyyPizBhKD1yWSrU8qTxJwwQKfMzmE2wSoWXRb8Re8jNoBmawKI/JvRdYM5B
lmYlE2RDXeM3PYEHSEDlcnZoO5sMpVZhpRdIsSQhnbHrxlX+DqZOixbWXtHxL1RqvgwRtcPyEn0n
QTjVHIMqAZTuqoPsLMdCaZXPJJeakCV2gsixTrggcI/Uw4EwiOPanyrUtrFy3n0GBpyxN6stfFQv
3tmFimaTxfrF83kCNbzyTubJWGUjEf7gv/46+rGQAdhCD+T9HsMIGXJ2whiYQC1Rl+Y7jW/ZZHMZ
NHY7RBYHewdVjfWzHFl/3MTQKpYVniTsueEHI327gC+ZllIRYYnPzCogoJCgSudspmKZjpnzTwiw
IBkvawebOuRQQRfjIdXbNvALLmeJMoyvMsrDExbJYdYXWbmeOzaXxmpakZOPcRZLgCWi2HIZb41I
/lxu+2D5iTVD1+01GJrzMcFErbp4jMpY1HPym5OcLu98Q3+xepTp5WaYR3L9yc6ebSXq4W2JUPvw
PetQKfUJg7+WkUVGfDPO67ZMzVzUUL+hHdxGItzQBv4F5AAv42B2b4A2382wkO/j78bKQkJv6EVZ
vLRPk6NaGLh6HZAieqbGwFc42RbpprLZmoVK+cGLGWvO6KuT93dgZrPooF8Dia4bTf11QpZiIhjQ
m67bixYjt9IK49KQIpJyGO/zLd5jgqIm05bj27q8gSG5ty3E5tq6yWxYsMN4kuvo6noziGC7YnxH
rfTX2cuWJjOLYXKiO7/yLS+u6BS0KEJI8giPha6uX/K/hljF+Z6BgheGsxLJKFKm4vYWoqSBE6DY
QpasZJ0izKZkY86pdSvN8wGCyjMirbPALNmkK4FjIgIvkAuhXMiv8zUA99+FbP6cuWcH0XQqUbG2
qA1aHmxLYsBOiS1V3XJUK14I49UczVpbWb2yaOMkgZBUHb+G46ThYui+ZQMbQrPUZgF/a5GBGX9c
EE9i54x2ZOwYImESFyWIJlT8bKR2YwLBjUFejjKHbcfn4xNCtxuIXSsLUSLdf2pG/S9L2Wg+d4ZT
hsbW3h+o81tAUXrkCW7pY9CfnXCEvbbi34yAOlOP7txmmQ9SJ9aN9EJKWNUBTy6aUgC7IcMudWql
um1ilCM0wmj6F5398zx+xY8Kpu9mqAxCwssNpdIDyjpHxKY5K0ftz6UeX2wmr8stNb3yDwEo6x3n
5zJ4Opjtx9LgGvrC72HBysBVZVYe3AmTBgsoSdjOkYv96hap1Z40SlgTY09mjnfwG6ZRIEHUAifZ
B2KR1pl6UcL2DFUrZ4wAoDS2iId0NQqgq5jr+dXtDCaHXnj1t+LibsZudjJk8vC2dt97ulJl1D99
XcBW4SRcLeZT29P/QqDOWGsijHFFqkwglqBFtEkQuFf4fLkj2jmyGu/4qFsHbz9wY/bLUstHY8uq
5BWpP8dyQpwOnz1RvRFaFkpGEqv1RrADBqxrACZ3BVe2Q3BT3TLqOhZs7wp8+V7rkXA/2QPXB6UQ
PkRnVNzWZcJ8QpIHFP4pdO433LqSl6altBjAvclTW9gfR/1PN7aLrS0J4JwFpr8zdXTQ8riWle+k
3O+7iBc+BmUbm4dCNLDzMXtmbxClRYvgNH3eqUJL9RiPuiy9lulSgw4xvDTsfTaedL90jsoiefhP
IQ0mko3CuynYyNO6tFhMsCVM1QwIu9Tc9baVUmAwq2fuktaVYGVlzT5DWpnJPk5mYiYEwsOEQUhI
YC8J8Plx7wTeS4/w8v4IOoGTNxrLvqrP2W3LNORHi7hzPM0Pd+9Oh9AKIzhnuIrvtUzyGku2nB/g
XmW0/3h+q/ouMyCa6rfHAZTfPXE2yZmTz5hc3SbPmmqPfMtPaF0+P9V88w0Ukkf0Y81gXpVLsIlS
WqiduprPtcG2zL2WUcw6vIeweVD7XbykSMrk+pQk7lkV1px81Gmkt7HLnFh7AkKpWnzjX3otHzCN
hgC/UAEN8AbHkLZ8G8FyCVmaSn6dgqWvAWtKvRUtfJySy+Cx5gbFMizBiDof5m47Lh9P0tQIFkA5
TnO9w1ucQkuFpfuE5X7UATMJuzLBK4cyX5VfZjcmhBg2mWmUvPX8rGGn8+8H1e4w7VfuTfnVKYuv
r9ko/vFEmiYZm1sLAD36HJsDK8OVvSZ32YqkHVBsaKoQ1+uUCHiqIiGka+7rjHA4NUYXNaXovoRE
V+2FI8vfzbnsD4BOvtp7lLFwuS5a+/4H0tv3NKV7jfTd0yndoIR+KtD4VvAiOyDsRH8uoePzyOGH
u+yM75n0jfGZj8uiXwY/hs/3vsfa63Fk7JlF9VfoYYtPnIf7dMcHrXxEgd37iUbOOyBacPp4uJu3
9RBI3Lllx4QSznPmHYh2IYLlKEFnXgobNVNAHh+qUj8+29wGezgod4t60b2f3Eu6gLcww5Gl9WfQ
xKYDOQGyg7TD+rDbODxPAFPL6ZoxaqzHoAG+8Vbt0gsB0FkSYcypjsiRk2ey76YyhhMWhgXzVUre
5b9D5DXszTk6F9vb2bh+VlID1pEmh00Hm+7U9vH22tq69COu4FvdzZAgVzK3Lz7A9QhGnNkgyicO
ZTKRQRuc8U6FoYBPCBVq2oi6QOzbnt7/nQoQujf/uDFVJMnOBQsNkGbaGhn1hbJ4EBZ+gbDvviiR
0CTd+1NWi/cg5qSfSMEISdAqm1izaPinX4wJVgpCFvtVg+XL/umpbP0EsRHoPyEFFDuscJ6TwPRp
wV6b+joh3j/2Liy4H6gCPeTqkshnpYYMGivsyvMVFZg0i6VpTu+w2I0XaxI1yk+YyOxUb9/ZOjf1
LrlJS2DCHtZt1olSi6GtAbJ+6J1ttciZkoOY1RTEZAIUwZHMdjk5+/KA1iL2N3Wmem0XkbgRIb+S
yZz0ke46OhmBA4VZOzqQMmoTGcqXe9cSliyJKWhLBaBvvmpJ5xcGtrQkDc5/Qggxi94HxVyiLyhy
e2JTe0rJzuqAsMknyeFmyeQOqNC09iEuhNIotbodDk+ox+RQjpqz4P32sS/vNlpnphiopFe+ThE+
SlY6RYjszUXSKC9UXXdksXjTqbZl2W0HSligPbmO3BwBs/OEWPvqKIqwxUVxhxcT+kFb4C1gBfHo
CLiipSz/bN0TCH5Wh+ot7ZFt8GVJiG5RI4o+oZVTN//HLJUNF9YfOylW9N5picPhP8vmnpSZq2UZ
jCBwSsESGqA3uDkDlaNn9/uKeghNPw7CkT2Qym8MnnTyTcHL2UoyTXvrGi6GqzRnG+M7UZTc933w
M7UYuDgMi/UIvrD3lXnG/+fmTLXZu/kCubHZTedfdmPHRoEp6VovDFYFm1XHS03hkwFETMubWAQl
8M350KXLs529wZCU1WQ9WLufQpgFGnbLGESyVOo1Yu8nh/xBDLmFR6xT8EXPx4X19f9Dr1JgOnqT
tQfOCJLudPOX0+540UMJViWnWMEZVDdIbQhL1jnovKcVIriTV5QERV3iM/JurAEp0YJMP5msPMQU
i1mrnXWuaQQ/dRMeYBRBgWIIX3mjHnf1fgZ57LPMBO+UIy7tKEcaMJHFprRxouMcQch0g29hQ9eH
Z/YtZBAK5WYCRkjy5s+9S9EMka8ZIZxMgRp2c4mx0CISGgGYVL4rnjMjZXTJB0we23K43VIZI8yX
TGyMG6WIU4TmxNIObU3a5AWNYmesQcthxOdcfGlBu4VWphfKldzux91TGIx5FVoYLhO002G636Or
U0igxnd8TBRnrV+F5SOYIxY3fBiDX/Y9EZ/Xisjpgnjr5hKzibeV5IxTWdZ2VWo0qO23Rs3htuK4
y5khKWrXJQwQ/izoggXKOSbFHLn7U+9Z7AGlTug5+utfBuGihvOC86hQ3/8kteNu3RRIJ9ufGdJc
raOntRRo7YxZamWizNT75EwOjoKeuUa+ujkhGRUs6mmVS4El7evRZ0tK+7qrKdCgeY55pJP8iQly
cAjCmHC4AKjfzsDB3G67XeFeZQ49UPGi8ocD5KeTYS4ruxhBrAAXK04m7rObKweaObHiFXdpTFb0
EGj/2ct5b2nT+sHghN6mzjQ3obYQfdaMFITuyBPzL6vpX+MjJsMnpz9RdYKJapuaKvUxDEc2GJZ1
uclSp6TTDbZ9gMkiZn+kB800JXPannLBBCsTH2QfYoL2QkxFB0HsZjL05JXgMqwh9g8CCwNvch15
465Eh4bzW+PN+aR2LgyDVmYh58zXYTR68BoKbgPGEheFFHxCJ/YY1U4GbMnPsSEO8Jem1yZsj+GV
jczDT8O2QwNx8eRs6Flwphs9A+bkWoOCoafFyJ4VMCB1NENHBVxiFrl+mCLLZlErVp4giSZp8KKd
ydnRN1Vaksrk9BsCQbZrmzrcaWamfK3UYcbcy4up+2iWVv4K545uC1Uxx1qPKhHq0pVmnPaznqS0
FOwitupfLlXmhU/dnxzlRXBo1/liga09T62Y4iuykx7lllXlWb8g1SHU27xc0b+YbcwWa4Gw78+g
p2kkg/NEwWmaVOnacXz83pCK5DZyGzyDWnTTqNQm0UgzI26wpPVcKBnHtqeSCicfgoGFO28BzBRT
Iw4lr3iYMNJ0oAcckVm3Acx1rY0eeBbxT9N2+OpXRBJ2FVINOXXIsXh55AFx7jfNUhSjZUUe91YN
4cvC1N4GmQAME7B7DU632kSrTbctP40vew9FkicZalT96Dlk9TnabiWZQofqNUjYExRzHl4u+uL2
YIys2/mC35952WqxjrffTnFaAtHhO1c+aU4S8i6H7MPZyBnYIQr1IHAEnHS0txbn6J2PIaz9KIxt
cbIXBG3385ov7UF4HNcrcywG6sVWwajN67o9BqxxFrjIvZYYyX3ic32gWux5Sva7Z8EBYCWbV7rK
u9CN5x1Xsi/BGVO/uUGBO0d9oPaNohnbdKYEjtIN+b1ej9pbLUGwvQlKL3c1gPqdQjjUCpznNqkg
SlZUxDO8LdFF531WuUC5Rohw4kEDjRLGWj0FVyPSHE8j0k/PZgVRD65VIPicDCklDL0HXxU25mRz
RhaZr8oTee3aQ2leNIiyJZBMvV9+ww8lzs7Hgbt86IBaImnHN3MzgDAUbs9w/yItU/p/fsCj+okI
fjhJ8AW1nej8SISixC8cfi6dO8TkYqdd+ZaC/BI/VB+vhwkJLt1SPdS8KKJ2HGJhhLYgnKjxyaQL
VWu0e+3ZmkF59Wpc7apvnu7EgtG2JSL4cMOeOUthELhb+i5JwSxoIUM2Xz+/EEMNOfloOTCD5qSF
99NAJZRCFISmmF8Wjl4ZVRzU0LAuJ/xNH0nwh0PM8O58wSpu1Ur3JJPtR4qltwiYfvG/yCA4Yz8J
haI1uW9byg4dM0uLUZHZKAX2uksQOJLM7KPrUlikDj4HBvws2bv4YORNqA3/cdNy5iqFO7dnGWa7
9SSqGbpaLQ1X1SSrEn4Ehpfl/IqO/rmyIV89Ipu0ynagFx0ZSz6QRAxj32aRO/cR0EmXfrDFMOs0
GFregwy2ujjV28Hd9w9KHR3XBfuEG08QRwjVAbjKW9IUYwgiqL18QyiHsdKr/6eh4XHXaBk4o3aH
8CuZqRuyHp523QSwylKQ0i/1qd6XRs0q0SqNRvqs43Uw31Og+DnIZ5QHDZCCJA1eTP9WaB60vwwt
UNKziXC/h8g8DT6GomONspto3jSx0Y0ifYg3ynrTue86CMzcPndVBf1TYH/8TBW9A3MaTPUTzXbR
G+/ndghHzz86IIlgtXG6LoQCTQhd+OMJaoYu5sLNQi9Du+se+iQsx2BkqWcH8uNLidu2Exse76t5
uCv1WTCJI1dGmGCYK778zZ8lfuco2d0jYbOqbZElueXve5Cm06PW0NSvMCChjt8g6rABjFPghzzl
6cJjS5nO4xbI2ecNUCYUcO3tZFDG5CB94zcUeKg0TAt2sJf4DqV5EfT8lmxjIYs3jXuwpkfUZrcK
VLolcE04mtVeDSaeeN8vrBlUCxZ2/MTrohdFCFd33ACYrrJxEcjhFOhhaO/nT9soDe56CPC0HV7i
RgRYoOdGhh17gp3SwI26Az1OTau8HmP5eUvtoJM5htDM1+QAdkFsrm9XZJWLUaQKt8xPM4+GCnNA
Pq73Jb1xzpHtcr4RYa0f9tdKHcWZkoUA0F7sKGws7f9VG0JrJkKrcw6gU3byDpfGfzpQDTjEP9ou
iKxpZ0mNmAQLJ2vSISKmmG8VIwMU2U39EcXUUR8ZClDUw/ggqNu3yLKHOrSE/w4aesboKk/dW8Br
PQnRCErh9Ff6ffWKi5oAq7PGAVIPbAJJll/NuRCWBVQqQUZNgS0L0P/PMhMXFTLLmqj56xWhLKoi
r3wFD3CVHz3JfeEYH/KzMQ3MafsKQ96hUeoeOnb60YF+sLN7GzWDqgv81nSLc6A5r6LxCQdxms9U
Rp4YyUtHXU87ioE79NOGqRJmC1AaAU2mW+Ck/v8jXs23jhijTQ0QytXiJon3Or1xluXciSsW9XdF
EgW8FE3Ny5sw4tm/JBTa5Sd8fxGL/ONTFjlEDtnJXYw5DifIS68bxeGQPq7DzjQ5G3OJuaONAeix
1ya7bNYfyd+iDLx6AMe+GmwpxQfqVKYKYDesgs3UpnPH+XYioE4trsfoB0qE+HUqTK7bp38Xng/Q
tLBf62qjXO6Tm3D2ZVWMvV4Lx2y8z/ltOHDzrurKB0N6ulWiJ1IXsT1Nhirhjes9SYXH5i5NjscP
0jwvUf/TsQq+NBztVd2CzY4D02OD3wzlD/9ImyolcWWQtPE+MpuRtHwEcberllqKaFZGkTNKe1mI
psErYa00v1UjkrxZ5OuQuQdO1StY5zhCKEzRGieZath4VArRuDZXhMEYPAiHuv/MmTAq1/fz/7Cz
4wNRqHekMcjF61+XGwZP6fgmCJmQHU+WuMRsGqdQvIIwnpJyT5JCGIbkNOzIDabDuUvXXe0GxTe/
txp64o3PcOe0FHRz3+BIf42nUFr9X0ox3iOM6sudTv+cYYRBEG4L082ioBMp326G+YnuzQVTJY4C
szQxr1yY4f7z65rcZL8sQhaGXHbLZGncY4/siZEFmpLo5C9THZEI3PM0nVpnsBrmanszrJabiXHs
B6YYSdnhEc2LGUFDAM23XyI+FV2Y1i88FFz6fAhA5xtRfFQga59+/6d+2geYVTxrgP8DV6w2/Re3
YPPinvCVy3YXt/HsofOZR77Fg6NGejUowudpPZpyOeHUWye7DsLS3W63EgL4Nrv1DwKM8aWn9WXY
Oea3oPmbHtRvubQgEQHXH6EkEwGfJ134xFHgbsUXdnwvhafq9BjvX1cSO1ki/sw1g5TlA4ai8oSs
RXKGA9KIF2qMdoYdnbGLHkfulkWxyRxxT0CH5ke8K6/MZP/WCnbi2t6sVCVpv9DRVcoAYazQ9J8h
dKeJXGjomBd53GHOc8NhkWId/8IAnFp3GlItm4+GGT8sFtRilDVj21wUoEtKU+ndpVHKFn7tErlT
7P5zItlMq9MxWtahlYIX99i8hiOXiVaF681oSy5wNCv02APgApDG+jXOrxUESmWea1JXnGP37Z5l
lefQ7wi9ptmYasbkZgZI+EzOfPYiTLQ+Hf2sEcDyhjo3lP/FGobml8zw55Rnu+y4Sow7f+NO0Ejm
hJjHEJ8HEHPHAx7B/feNkPY251/mB1vIobt1jzz15dHuMqRH4y7oFdBT+1Oy3LelqaSbR1m/PpDt
r77X0YkRHIJrDyD0WuFtL5T7Hy9Vk/IHEMNY+VefzYK/QHXALMDjdvO0x9JXCby6ovQG1Z+JqBtS
zn73a1fSwtG1YFuQkirmuZOsS0nzfrLyYdutrvQZv3wV1iGtTBM3dVjvIZinfEa5VPMB5zjuKiLA
HitAfgEAbgcA4vulk1FuSA+yL1nINiAALFc6K6TbRHI0TzPGTBPwomoGBI9Mfm3iZZV8Z46W7gP2
BTSb/cHbCPsQIzyw6x1fC8XCoWGTPSly6MKib3o/KsmI69iWUxXJoi3RmkoiWy92b5136FXKLMaa
ZPh0TZWclRDGAJqU9z6GD7kRxr7hZySyK5B9nf/tm2yvFk9/jKk2IWlVtu4Seecx5rCI10bEiRO4
0F6aDydtadgYb8cgb2K5mRyoc9SwMCkqa8ogw2WU+6/Sv79rqGTC93pI0iSzYJIrHuWKMni05n1l
MP+VrdadmAxgaGrNOElqmYYMLNfVCGiaIHsxgaL4fq2nReH4hl44xZiulbIO8CyttIyKEIY2hL6L
o13vW9JnCtjCLeTXnKo5G40LrNGzpq21I31HmAqgUFnITIszSTxLVPw3pESn/Xx+xya0FCaJwnK7
hrZP01ll9RNJhLvtoe8iE3Th516hPVr0XmJcuZYF9L/5jeGlta9hC/Rl1xywWsJNcJ7COYrRsJrm
Z6lx4lLZrjbXkvwChbzh+wIwyIlYLZTxvgpfneLW4gU+owuJkEhRL/90m7e7Ye1WeoWHm59JZDxq
SPXUS44lxGn9pZ2b40ynG1w5iFOKSTEx3Rp4fdVErMMfPgXQX+M7GKBVZu14ynPOqUUoU2cI1eUr
XhuUhATLUJBjHBI6yLu6iC55pA2bVFLSNxCv3Onty9hpMJyd6ReXqLuMfYoxlHrDDv5BZUWX9O0V
Pn5DrWW5Buz/P68JgwGlunoMph1vswmujfQcV8XyBGShbLZtHOiucpD8zkij6rT3TUHwtRDfdl7w
YDQBdoryp5HXAwffbprn9sAIMblKvyW9bHQ+C1NdAF15NQzeijs7CT31uUZTk7/JGHHGMEXB2S5E
yrbPpoZhDxtc8BCQS7Y5IcAVKffE0Ztlt1PJqnxAEND/C3omWtoZZooo+U93mEJRdkuhipQtbs5n
TFF++QU82A+hn0u23bUFf886zYTU+Rmktd2mTcI/DUbOHEQDU28KKIHinevkx9aFy8yU0LH7yccI
MB05KCv54wAShVs+qjlA1wSus2hKIK7xSVzwRMGT3EBGpse4nMxhfsl+2xMuNhsLmaecSsKvPbFg
MGBJWjQLwXDSjW7rmL4UrLVmxWDna0rZ5B56RKqwCZHgzy7SUu3E4Qks1SbE15LAw/f46ljO2TZ1
xlWYAu/Nk/rpddRZ4nNfLZY8f7Nr9Y7W0Ft76V0cpoRpdPgVg6bpwGeNX3f04t1pOV+OcdeV3zHG
DJ2+tSWWhuytqfgdt2PCky+x8l5lCjzJNuywgydHn3KNoHs0xFmi30xm4uPMwkNO3dK1am39I4GB
EXDPxGk+WkP9e8UM84TjAjjmKhJ3j4LOxBkiBXMyOsYpKt5Vhi8B1onmEm74Pd89bTrNRn1j4Kqj
u2/bU6VMTEJyI+kogQexlTL+86FlIzT8ZT+K21znbslLyRTMO5d8kV0TKk8RnVK3UHCnMmyOe1pN
g2SQBOjTIjb5zb+F8iIeSsEr8ecpw7Rm604aqi4MhvMspOsNKz/VVQIDquQ5j4Tm9P6DMxftoPLV
XfUwnH1SxaKsf+tQsSNINkjpnK673WXgIMNvuTbUsXMNFFTqPGKHWOin9/Oe8YpSMYnAnWOupSW5
IhZ7OxCwCRjA4ODhKKmu9esQP2JbZxtbWP3wMAJ8luA7RYB9qNh/M1/7T4R0GYRiJ0zm5xZx7tkU
+yLXPF6/ixwV/DMYNKFJ1VpVZgfRiKG0hVZ6Cxk/5feq8RAaF5+FCim6s3kPX/VWM/HbE0YYUuAO
U49rZekO4VuKEzZuSfXTbNIMTe0M+Z4nfpLn5WDLcnq28XXlsnGGb+y0BGuooC18ktHd3b5DNqrX
1wVuYQcHrOUTtBA35TnA9uHF70dvP+CkipNxH0eEkSKORPoKg2wlqKjnxKRyQUxoUL9wVE1RGH8u
OwkglBwbWDyGhgV3UEApQWJ4Zru0td7Njxd6+zJveAr5PicqSJHY3hwp0K/TT7V+qawJ2ZUWO5te
pmIIRmI5CHc0nTQ3DfEZ8qTi4IRLslXNhDBPgsw8tEUhcmisdMSmuXhIcsS+WSspRNACZZWT4HcZ
fk/vFnAeac8GIosgT6w9gB/fY7oVJAcV2gI04VrQOhfKloma3O3H08vEfK46QYYGvxZ9BmYClGVC
PXbhgWThJGNwN07mDVmqgzEcyurNuUVq1lrOmqIUq8HrxtMIOR7tQNFgKuCJOJHVmksRnhWPMTUL
GqopOn3tEUIrRf2KKYZTNq9pwkMrGAAQwmvG9Qpm5UEqp2SGKqPEy9Wwnbeqx3GYB6cxBDeopmES
SNLFVnrw3cGSOt5+iVezl7k905v8JPEvL+JWrYGHCsA6oQFrm27Obw8q84xhiLm1tD793IfCOw3X
mi0OYu4f8Kuae2NiBEh6LQpIENXd5aino67p8azlFcMgtsjiBfBeQFMo9F6ygK8cVIKOhc7Tf09q
mtpT60PRi3AzX23j+OrUID+ALQAifCx7rUno+iJaIOiy/x6HZTRgyN6hSI9BL80pTIFy1bRoNtzt
B7baQ0ofbYGjiEzbWEcwBggeae8qmkWMTJdSxXlGF7bpSOaMCmQXe4WnBCo6nO26rs/It5A9HJ1x
6Dk8zjkij0fsDswslD4V4sesB97qrh9lP1tl1Tgl8xh8om2MSaWwog00PYenbPF1FxGc4rNR1Uyh
Jj6dAqgk7WbxsIfUHjAdi7ANuLgW32g2BSEanAzjUw0t3cnGLAL4TL9mTK+kRUhGdyvW7GUfXnKS
7kFLfYpzqLS1tVhx/GblQkENig/AmzWHEyqdRnLrWp0j89dq0LuHi5H9jtXsqDFwIBXXOCqnm+LA
0mR4J+/pbXYohk6gIPiJySVS1uHGObjNOYoM184+SB18BteaByi27lkC4N0bdTIEHTAgiJbqfndx
8prd9jRUijodTYn4ymVyMscAot85QiOeVGEWEl2MYeQLdcSm6wmjzdFntcBjFCRT4oNX317VFVX5
RrgQ6EsqWM12J0jJ4mAJ3DzG5ai5UrKUvLRdqW5T9/ageaN+Dek0lWmnyhqNqnUTZjIaHu5Jq4JI
n+WGbKU0WYfsS9/3sbhhB2UxcMScY+wegmlCMD+cDzBa5ZZsgCS7DYbQYhDeKjbilEdDsRM+zl38
Avsoui+vskYqlTouotWAU60AlgDKA5TqTg5mVlpgJ0sjVHeZhapBxgA3Ky8h6pl1irXjripGX09V
15K8avpUEpQNlDq3ipMm4OCWOEWskgdApYg2BRnzlVboidekCNh3Mu9urfNnCDwzBPBvYMAm2UOH
uWCtc9oRwMxLuPZNRJxU7pXJy2xq2YxvxhJA29eah1VYoVhnYyu2Kn5GsGnoQr3rnBdJOBdmsByh
/thkmgb8Y5z5PB7qpVCmViHgbr0uVMSzdekF/rJ6vDxwvOmtEXYGSMR2yV6/8z9FNJptxDs5diuz
UwvxfXxeSPbtHbwvzeWhObTfufNPm6qhznYhR96zwaE5r1Mhu0cJr0USKAp3Hu6FLqy3+nI2FEJC
/sUPavF/eXCc3KOqrCMfJhlqK7+xStuRWVoNr26girR+ZuSz1SpqfNmIBTSvB4FjNVBCgP8CEB6a
P8wNic7HOvx2XuYc819t+Vq54eShn/fU/zVqm29geb5AVCBkvV07F9WbCEX8xLEVlcqwLnbgwh8P
4atDtqRD4ir9aGYQN/FUnArPGlPuIXVQ9XMvgbX47bSdm3tUgxK64IHmhiBlNrMBjER6QJMt0sUH
Ybr+Lu/tAzlx7FPgVMdJgwLFpSA3qp1awrRjCMoBdONGuVjM78+h/pg5etoAPqexQYjoU43rzkfJ
Id+3mecVb6L1x8Wt0F68cxFETVRspYAqXq/N/fODHLP/T5TrU8ya4Uo0nUQ752kkUgtrBeSl/XAo
DoWIPra3pQB0gDOXYzfSQ4tX01ID06A/gqYX4QMWEjgWwMhqsBHQQOJWohMfNDocoRUbwzILSsY/
oa3WQkfb58p/gU68U7YcLfEq+Tq7Kj6pVKIP1jRB1ZSn+NJrv4gXI7XtEgTpxNMtrE7YQUa24TGp
rJTfrohv2hnMLd6SUeJirBphdmZKBYxlE+sVqwRTfbHEpuOuLwg5tCzqgi0lgnvwlkwsFctkOfns
UUjIZxjb3GSVWjKmGGLmxXOlwepSyawL3GycM3Lji2Yrgkg2gCAIgykn74OvgR8zD4YuW6DZiv2F
+DkAmdYmmRYFzMsi0WGV06FLBOAMVtrvG4NPj0PUnD7J+RP7Ey4AUCdg1cexCcC9FTbWOofcfBl9
GKMEPd0fmLzY/xtMO519+N1Ld3tdQSsucopa+wlQOXEBhIcM6nKWoLRN/KXyuhWXYgzJuXl5KJ8Z
KhYCNUG2TMn+oJDWUk1bV2J7BjWcuA69nSk9DVQ8ORDCMCaac09LTy4r04Hu8vume788dCXlzIYD
bfmOhBKzgt+5vKJkSoPT2WvelUvSbtXz+KItncLh6EKEZFTblVurVcYynIu56i76T1mBG0u6Qs3R
LDrwebRzuBv1BmjMBp0JHsyVyra97DQgoJ82RVg/zHLFowVjK2iMuadi84BxZZPr/tl6aJ/tVyCQ
fZ5/3Kq7jIEbeDKrvF1ilYgZpCQIhkYi5XHNE/GtiRNCPONVKRLJGVP3zPBiMjbRlwqegCS0w6Zx
Fn1vkZKiJwT5LZNNy26fkCxvtubeCVkeDjyLpY47C64OiRNTsZ/z5ugt8vNJr3Ks6rufmUy0KjvK
HSKy6j9adlAlCQSGMG3/Xq6g9qfuRBsPT1mIidoRpsl12dyHnELJeDTNUUGnqYvBX536BrbK13UK
1LpZlqV8WSpC7ttmmi6dfbMxA04yRl7Y5H2qQWrNVX7yH0N+aNal0tbfbrMRLvBMaFa9BJevn+cC
Mu8A17f5oNVozLRzBnXrg99lp5YfNaooPSYnpTCBRqLp+//clsNeqWekVLsyQQ+zyF78uWI/qrIZ
/bgUXnToOKZRtc0HhkQmcxCipmijzTAm39/xYNVzzqXQzb4IoTUIXSvHwkHINLSBzS7mVkFbVlLv
WkkFHvCBdXc4fihm0u6Ri6jtp1RFMHuVBvWJd/eVfSiOQmr0TWHPUnu6bACg5XRWhrtmI1S2IspD
PalY5sKyOTiECSnjACUntWBQwvSRbOtIwvdr9kRjnskOTVvfkYhoi+VojLDRlC9+uFWfqDNJLvnr
t0aiwJJXAnSrKnf8sqQ++JrZ/wwwP2XqKavUL/yTK121SKWDWkKsfL4pn7fgNnnAsOOW8ZSIHQf9
1qKj/RgHKLw7lJUPgU6MK3TUw+XcD8wqjATrWdH/vpb5KTDwntWl1CLP4uQdvUvZd7gm+IvuFsnP
hqOsVtDFpsV+x7raEALCLirRcEhNWGv09tgGUtT6OWBPhm6s/Y3G2KIPQz++IXVqZu07Q0cTJkFi
HwQGTtnY3Qe19Iup7FgASFLwxXg20+1Z8XE3KCHPlk2G5h1ASE1cNMjmJ5QKRl2ExazqUdBKXZRH
AnWtN+FNGNehFiPVw7tKSbLmQ0uClUZfT4aDzONfThN6rfoCheQOyKjFFGOCDB/XMt4M+o04gOFj
UTVEXtKlArXJnnGztvAoh4r3cgKJrN79aQs4yWraRfjDZNmorZXmwbGtU9uTzq3rDsnpMGz/ZFYR
6pBvh4T0Gyf8Z6rtw4UdAYPYF/3H5s28bvMsYlkbT3WM/zHiSvEeOOoLqp0lBg2G3QTVoMJV8ptJ
of8/NWeAlLpT7uEPmYFL9MNUcnUqFM/EP6P2X2HBGxQqJaeq9lfo/ZGjyuONrQwylCZOUFC6TtJU
zNKZUeG4v49XZwhvDor+xdAkFio+/uhlSXLCws6AKdxj66xSTT6qCUiUtCl3QpEvjkZbMoS8LmmU
0cxBzT/2CdqJU639DMwglyFqbS0T9eMhdJHexyKGXqkDpIuR9quUBRpV3L8KZHuAuZQXVqQKHHUf
AulKmQZ+bFJ/gK297iGBhNpZf/BkafjxxsdfSYGEiyQDByQJOqKQw0gVYSqehVsfdKViHt5oAKiB
QHwN9xAPqcwt2Scc7Ruzbc9ONPx8SaQfmLCGUMjz53w9803Prkgef/AOIetjfScVUfqDo41v2MYt
4Q2s6TRyPLDBKE213QLtyXLoiAG3Mrxg2mhCL1ykmU7szGgK1kXitgCfwugNvtBJKAefv9MhEe9m
sfBmYUT/90rIBQIAeTTs2OBKusELEqOgFm8UzQV65hGRaqlyP4GYLwiuHOeFR6roj3HnwxBMlktB
tEy8sqtdoDIhlnF8t0GCI0Z/tcOqZ6RuYHeP7T2yzf0AgjJ+iO6R9cj7ic2QCwLjZJ83fDi7WpEJ
n09M+qABA7hD4DDtIXUKkUmRNMp/tjymPBIrDX2H5FvSQNmM2YmubgXGcmXVd35SEzHv4C3D50l2
JkDRwmgPC4jJTfbhFVjO830RpkDjl8+8d+psGYPXIb09YX8MTL0UCZznQo/bJdCjKF/eoWPEWVFI
HQODxqdZ8UTbLEDF74fUoycCvPVSe+6OFIVde1G8QSqrEcxxjcjkHvoU+v+tcWCKR5tQkFqubSSx
uksDf4Z09tSsJbPCJxdrW29VEhNURgLbU2CnzZvfuktP4WH+s6BluSczgbvI7FFHjZ8+eL8He9b5
aHvVVPZDAE/pfOjaAXLF04Kpj3ZgfSp8W9JGucEjMV5n2m98AD3Sn4dH1ytT7ZfI8OWWkgpFzYOy
M1CWWMWXVmoFl+hy1hJ8HV4wKzEr7u29uVMdDoKQvRC2EBVStfMRKaLQf/dUR19n68F7fgfUuzPo
EJ/67nUleioKHkIFDxHUHxafIJBJG8Kw1lrT8EfRNQm5DwKSc+2kstoWah7Op9fIVhJrZMPcf6zc
XcUCjQJfGlq5Nbvdf9pCS2zQU39gI/tfoTJVK7eEvRwSaqPyIx4eRGzpX9aMfErvHjsGT4Z6ssoa
NzQTROZA9kO45OPk8F3dEdJtB+B1QzvaIXywJ4bp0qtXbiB5cxP0iFtee+bM0RANqJc6CVeEkGkd
tK674txkFUy1lWezFsHVoQlm9mXTWM3jE9R3KQnDDflhnXupAGVpChAj0IcgDRqThDoK+l6RjzRP
sm1+WfEPdXUsDRlC/gEmdnkf59ICd656OnYJNXlNO7ce7SGkJiowsvYm/Kjl4+nTeidkgcI/ZnEf
H18oEVpc+2gfCeR9PNNk9ce16+BOTZixFKbBQzNQ5dqgq4qxfwZPMq7rglrP7g6Cz2UTI9izKkW4
1mdgGAtV7WlJ503AV0MQvZFuavkWOMwhWdFFDhcJHWfoCrpAk9G2gTQBSLU414HGOqlRhcQ63uWw
b7hbOM/zd1zUM7HU0CQADiwb5YGsxeR6I66AyB8qPA1Zeb2Zd/vnt/wqGlRWWrVsh5rDKpaNHhe6
kBxODr11sQj5jMsQYLjclqs38hA8CLQFBqVjvwD3gw77e5tosTKEPtP1vYcU/PK/3Gw8ih2Iav9G
6Yh5MCkL/mwc//cT7SDVFegLAosmrpNkp0rwv+LobamULFrNiNJ9rHnWFSk5TtuCWVYNm+1pbEDW
i8QobslvvzdG7CYdwaKiEIo7z1/KcUM8kLLZ3ZPYbx/XA9JfEef05kQMg8JW+9EczR+WkWvUswBU
EZuZiMEwTfOzL0Xesbhozi7oJw4QLT5eSn/Ynp/tz6He8IR89ck/GV7IBuQKFSWrJR0xQ+QKZ07h
r+IxMIuq6FsmHvSV+IwRjFtQ98ZxDf5CR8WKrfDgrWxRPK7cN3EwUxK/NnkI9I27DgmGzSWrRnBY
lKdqHCcGiS0FEbzdAnY8xoAZv82wz886CvU1sqg5YWat29MKs9oEQ2cysBrOTij0USfeMMHzrBYw
/elRGdjjjLUlOB7Bj8YjFrlXQJvGNB+U+iJBb31V2NvV1K+i7d2Q0mrM9Cgcjqcc4phbVmf2H9DJ
hsTe+rz2Kc2Ju0URAUK5gUk27B6K+Gs8j5LOVA5QRGrVs1SjACcRKfK8IHnUjPMj/4o/Bo+0RABI
L8VIJrc3GV0tvLz71AamkOnGGAohbaFGTB8iUzszDZTW8/HlcLdmrhX0WB4kzIEv82C4CqJaNvCj
BulBnLmJCn6Q959dReQiQXu0GIxFhgi5UejYfc1f3T/tYmhPqmdbRkqjX7inCCSIfGcLFbijb+uj
t57sKyOiTPREV18GpAGvBHzWfAeGIkZNNXCqlTF+7qPECZQc6mo4OdljmmFmqZzV84hPNyzYrJM1
ocT0TaHIeTTmxXro7+c0hOby1micSTmfOsRJpsFaPl7ACAr4EMu4yXIATD0+RjpmbIVNQanK73Bk
IiDotg9o2DiQeQs4LG3+59JoIHDaaLB2/vFdVyTkMFIbGlreMe/WR6BTsJPYC8blVgm4oDrAhekH
CiRTvtcu6xaoyrwKuI83GK7XVE+FDNZtiyX/+JfmjOaUdnSWWrQQYV174x2ajXscbPYZI9k6x7/C
CVypI2cGYHAxYRYKtxfWhD+2mxbXp66Rtnegov3/aVirau4YAQNjmJZd2E2N8C7Rsb0ZlG4hp+Zt
XwwID+yF8dRqgINsUW+GBi8l2sMHiIGd2V1vBZghmAiX/DbYEAXa1fTxjJFn8X3pGNx3o5aZpUwz
7JUk8a1xob1af+TMbYX4RUTixqsCwLc7bF6a+wU+n52slLBQhWWvGSO0Km0ddomqUSUrA5mpqhwG
DDj+LSXPSgAJIwogAwQ3VHeIHUt77c0YchHGFxl4RJdFPT6vKkIgFkHPVN01FnvxTFnANtZbAIvy
wUOfq6C3RPrs0cdRmJ/aWj6BlBAoTm/ck0AQoW230+21m1HCzFR2zvLxn+UaL0SOToLtPW5YProk
hPoMtHbwc6KiW3GzD4KqacpH0HH1pmR52HO9yIK/7aTubAlZJp7UP1gqJg76AcVaLfkS4bJ3fdOz
NZR5+CltPQv/5Urw+ozQMb8GV0z+fk9AoUWGdVLWUTI71TGT3c7lOOn91D/eZwoKtQhgTXOO0eAg
uVHcAK2JrHBSAHaBzyB/GgdJL0QBLf6oex5CA07yuszcx+WZtymOGllglhiMSjmu9x4tU4fBspJd
dkQyGyFVolRSS4FdyCZlVw3j4xzPnw02RvUpKvgfAx8NaLWxhNRhjmOX8XxAFYX+fCsgT5nVCDfV
TQd8E7hA5Y/F1rR1CnrOlcujn9PJWpMtVDhCzOuoYlHtpUlBgeLnQzHSwD0qUEmncOV8BKwr/6Xq
QEl609uRgMQ//lgs3mh/vMFKj8L9AA/uEQwNa1S/B9O0/qgkGsGcwNWoBV0Cjb4V3L132Lo6WnA2
Q3KCljSv1bPf3FMEz4XgS0Fk2tsld2IPJMI6R12zWK6n8KE+eECFCSvleCMcTSYoxjNXj6l4vKF6
Qo08+uHCdtWx3ro43uyoThw67LN3tsPQm7Q7Wbf4ptKcAv2AgOW4EvdVa2TMGZ1LrSOEtCpuXblk
Tjvu2AlzaIhn4pQtMGLKACjpod273iQFbR/9d5ZGNgB7NODRrw40L05mPA2fDEPYsbGJHnjCzlDD
mHawev2LDEbAu/tDURIWp40RZs4UYe6TBvnMzF8P5WqH1/17Iw++CJx6NQEqmWZ2TxnSs4QjCPoN
5C8T0Fl5BCxusaReVQaZs/V/YeTP9XVv77Y2CvtZ8VhqHG4CIUa4lsNFhf35W4llE1fmsoC5xJpt
LGNXgZrHgkMgoUCWFtcAIli4Qb0QEWcZEgtT7Q6CQpzhV+h/E9VwKsl6/ud6uYiwUM7tJNxYa1V5
NRH1k9LexPta/v86i6tbC/08cco3Thss7Ecc+jBpGpOaXslHHq0UVwBQIUqbE1E9kBrUxfQ9C83+
xZEPNtWapLKvjrdy4X15uumI/sXGiZFEQnSfjC+D30ZZJWZJHhjKdjp+vn3xe3mrCb5/QCMsqxny
+4DliYX2c6iCQZ0tKRDwr57fe+L72Wf4Slv2QK7bW6+hSdN9Y3ikDFs0/iniFEAjOb52BceKmB8T
jWqk6fcK23qVYZaqihATTqxndHvDDukR58mhGWTpDhDaCr8NqJP34lYoq3Umc3LEL7LV+ooLB/lY
JYLRO3nvsNErbFD1JQodZZebCCgWxNS/ws1a8ZHAc5PuXK2ohjvF4gCprOU3EU5p9SoKszr36ZiZ
1BTs2B8iQYPnMxWE3Yo+QdvYFFgODKdG8lYxBZVQXOtPbkzTfEtz1BBf/XXqOGJVXX5H4IH9OlS3
DhkJGkEC+B7jqvxHnZjGM+S90wde6HkmO3mXOctq7ET9iGIzSDpyy+StnMW4i12s7HEA34WpR/7U
wAF3mCWY+NYRytW3qqpaD/Ms2rlTBnE9LZ72u58DtXSgutvwY68aCJ1KhKcGQ84PEpNfCchwKIjl
wMsJr+/2pBOziVPvykaAtuz37AsK24sYey8eqGh1OgWCaf/0MoWp+xxGkkc3VPkDiUuT9vtkuS3o
rGX0nACH1vZqYpJB9ZSuAfVtuRHpaco0cElyRg8BPpixCaU6PK3M6Qiw6MguaMoI1FE6yCbASJIK
paSiAJ86RuhvESCOBuG6rcuQ1Cn7Nq9lqwsKpi80WPLr482qD0daz0j4qduKyTZAZ/3byksD7QBp
+TDmlil6B0NlEOLpbhEIhA+ymBH7QHonJ4rfCCedKfeVZBblsg3ADYIYGUoROYgFxH+YanqVd+3l
fq1ln7h1VlRJPcNJN2o8tg9mlJtCjVgnP8lxS7nTdAZTLSLDgmOlEssxSmiYSlnAD67w2FvKni6p
SDj+S3SQvY9OrCPB0XDyw9pI4cVE7SvDMaGBAzUgOjxvPCtqsVao936qxvwoJ6js8LyDyfI7yEcy
UN2TtgbgJG+70L9JZY3EOPyH7fahkDGg/9XsIuCuESkkG5RVTqd2rafQ661Vzlo1S3b250xsT6Qs
v6FgM+ymIBzHSACpRchjPLhYenj4l09lGEVV9hSHdstBxQa9s6T7+GUNEvup0pzEDUm2ezRJMXFk
WAA29S4afvgLBDFVKfV5UxOkFlxosWRdOfWTh4SwSaq9kqRZ66PcNKkgaUpe9zXz6YdadgepwjEe
0JNvZNtFKduyAxVjqijSesB8RdhWeb3tRikbu5XWZ4qGcefl6hzXQaI8S36bEpRAudK4dnDlcDyp
c0iFkVZCWzUkfpgnrD2E8KRLXgmgqpQ4qiZZCzq0Il+8u68B+cOiYqlxPQ1hlh22QsLvzi3avUNV
wa0tn7WwXZm0vX+uFMMQ/AzWEKtnTHpSUZPGMslM/03DWY80ejdwbaVNsVJ4ycuIZ9h/Q8GGa9oI
z/oBuMCM6OlA+1gTZVqcJPP2QSI/vGYg922QRMKXCcL3WwVPF65CSM699Pzb/FXkWNa1T1BqmbV2
hzHapdqKVl3lCDtuxqyiOPimj9ZlkXnyDLiuxX+PpBbtxbVZwcMGhf1pZD37Yud79+IZ4ndmIRx1
OGs8uFN7ypSr2C88kddie1gB/z+1Qx1UZVVZUxIFRLeysxKmuarXWFe2IjA71DmvLHJK+L84bmDS
EOnseYiyYwVjczoe4WxzShrzFmJiuf+GqXvoWqvmD267QPLucl5ENVDZYxN/EG4z1lFM3XzgUllZ
mMkv1RnLk/d+hEKCNdaQ8A294fIuxzCq1bFSM27dcwObEt59tL7z8hZDQU+PiIMxSHqJvGqBELCL
jAApEMfDKUbGQZ9rCC+IAuyXZosMz/hQpvTZtSJKLvUrGilg0uDoTXaaVf+e0FkWFjSZRweBwdp2
2AOMkH0w//goQBNnoiXb0J45iNOhGD0H0msJXQJOdlRW4KUC3SD3AD/Jjf7YXwTtyoHF6Ua489zd
XTZC4vgDLO9NU+PEdtzAX9WVXIgkUFvNnphbf4FGAxAC5z8IlH/eo8t8ZquaiFUWlvdQlLU0YOmt
uSYcogcGjZWh3veSjIuyWyVcc9E8iy6W64Qck0TyFxc3HiGB21YD7p9fXNz8Z+rR+8H/ItTpKOqQ
qIvmWUoUYFN6Az5cPYUDPfCUmip5+TG2Rliyy2BAHHFCEisM4UG6YNj6L7o4+DiqBtdlLh1H5RDZ
f8GGHBOIdGEbx+/lv2fn0cS0wJ9X4rHYl/SXcPvYD1zvlgGUUxizO72VSIFEFx3EscLzRrLVci/+
I1MEFUOB0NZ6pYSnR4v5OlcKp9umr41vBk2ZfDoN7mCmB3WqXh+U7KFP9IqU3ON/UcCZtnfkjPA6
GxdUFdN+YAiIWUACDv1iqyP+YQqA7jAduMvJi1SIGnWkGozgPmQdWisDEmWj90Bn2anY31QXdSdU
LDvtxjLFyeTQhROE0TvxwrQRcnYN3i/p/lXLmfBkS2qoqzO+TgTUlYCktGXXWqtKz67niwCytXEs
05P++TStb8CCsd+yaf3shNBofB7ZqKFhOmSPS1LnGWZ2xVkK8+Pl3sqQ0gBF6dW26FBvmI54bp12
zMW0Slx1D57Kl9xoOeGJEGDsWZVKzzp0G02IaXjRG6shWmc0MK5MSRtNJ+Iqo5dvzMG8pz9TNaU+
DyqyasMfevthr9+/gxCRmerx/ASFNC2ZAuH16u2Zr1gh5A/q8LXtHg1+kOo1OrkLcBj3hMwoeHKX
0wDbHX8kqELfQ8xkRoDRWOfkVAOx0sB9onANT0Zux76JgSlyjqXaf9i3iP8IXUd/12pDUbtoVNDe
CUB23k3gr0Yvnq6Pq5g/9UxJDBgQR9lhCmiR69p2MWKbgrYjj7+6vxwSnoNCF+ZiUEWxKbxhmfyW
vkfvxjZYn5G7Xb1BXJ4tkOxziLC39WTcPTh8P0oyiFK7qIOhpUQtaaDnCX1sAfDueBrAcpd0BC2d
fK6zUMIp7PO3fFwdY3pOeY9tD0wtwe1gMHIsgZCxIyZuA8YedZBBfISs4zx8PR5L2kyu2Dh3hNpT
Wcy1DGCWL5ILIcse9+GMpqqsEkgWxZUZLC2L46LDtdeX5wt7/CmwYjo9QaHaaMvI2A/GWndr1J40
MIAbuXWkXTEMVmKkvhFuPZGLTwH+UyaWFw90nCrrAI7wHir5jYD/pv29HxO6ZPey2xHUuiLZ6A0E
Wy2diH4XnU7hSCmJz4Mhbz/8YQA9uYAiOJxduwyPTVMxsaqnxJetRloGT2SC61It/jGY4WpqddLJ
VMkeVF708am3mTM8uWKz4/PhzQschL9mb/W7Z0YsDuIAJE+vCPEDgy15fuINCl97WIrgO2g3PAEB
Ul7VUW2DX0ytstUyYYv6nLfdAWNF08DlwyWxLOShM6KmauqsY/9EjRuD5OgexFhkiW1IvbsgOyOU
xXLC15CqfIzO5olro24gtr93NBwi6koD0KBBKLsE4xgQsMAJJdGdD6t0Kz6Ff36yhsxMAO1enEaN
Q4aPKDPDpCU2EpUSkXmKRQL0eSzipA496cCe/HtcNz9riNftEPl/2dYGQVhA/jD3gFqSt7wt9iIq
I5pVQKpU80jlNuCqXg/yJ+BBbuePgqdlts49jg39NhsGopSal1Sv4iHtCpUS4EScJ4peysQ0pbKm
vZf9LshmE/1rasKaTr9t2hW14EjYHxkdRYH1viP2oavMl65Sd9rE+plCbQ92tbtZP3vA0zHBfnuU
0rkn6DRpihjqlXiSxOLhJFDQYH4fIeTY+kXtlnj7skrZM+hoLh/2JclJxXuZ3Pwn9paUHluYJ4kO
XSZnFDw8RFItmo3vihqANb+sDfxXlkB/8v83MjF4LQs1Qsz3g3LStHTtNLXvkYd2h8KGlauTcsn9
2Re+OS0IVQhlIlm7migpAyARgsaarMizONjPYiwSKlH0u2ZaCLctsm9GWsXbfhch6qlbrJWJULAj
bcb9/1RX+MxuamhpYWQBKMEOy5LOC2kciNR755LRYVpXn6bdQyaWtUEyqywRNX9oWu3fnbiapis2
FZnTPFSLBQzGG8ziJ1lHQSQ0tLz2/jaLzIf7Pl/KeSR50LGjClNkg4wk86PWNtNn+e3X+D0N6uZA
YguIcsKI7unewkAU9jWRYsbS921TPZGMJPP4JYWczjSOlhqjghon4izenmaCo5mmFWQHKCUKZRZr
ByejTU9DzcVR6qi0E7ZOnsRWE3AGHeBDZc9lqB2p5L6E47mwmjdQCCDdS9/pa7EQ23sM4DaNbd9L
gcfrvVXOVRBLa1SBRLxdfVNIzIVvybr0v6stGm/se16hho+eNtCUKtscP/EFqO70VzoaC+JZOiZz
/zUhWxr0TddMEnxGYM7gPkJLtMofDQT5/ZH/mxDhsO7xGKwfJy3n5RkTROY4qUq/Hwicpb5UqE+g
sqkYNEnocd9A6Sc4kBCj7ak6KKXNOl4aPeGsRs8qFoPxbHMDhDAXGT9XtW+xk+QDmXTNfCNgOc5Y
irOOizsMxl82kXdWy6QrxyTAu/hI0O5VGofFF9esMZdEef+klociMeyrx2OXfvbU5DmFlUMkEZ4d
wiev/3T1IJfnmydMilSwxT+YpCRJUlYqAKzizPEgvpaHP/ttzp6XZIzAe+HQMU7WIYKLrTo0r1UX
xu+ZqFnT7eDi+8TCUjRp/ox1F5XSnN433M6tQ0y3HWbUlEycr9qqBVp5MQeTq6nwH397qyz7PwUq
fdMQ97TEXpVGFY1iStWQlj1Egb35U2HeJ3FU7PogpwSJK5VZAef8rnGFy6E9p5QIIqCzbBUXMdnT
EFklcvA2/Oq5qeAFn+ETuxyqHDVUVcyVj107YJj8i9wOSDxiHZJsT/G50BiNExLmJUxa00JNX8yg
qlD5wbCe40fcD6zQaPoEeDDj9Z9fZiD2RMBBpiERXdsMESJ8xLRGbZqYHrcnVTUXpW4ogzjQsj36
ZYgXR2rSV0rysk1t7fUiNcYKLKe2xNUZV8KBACr+H9Nes40+oWCXrPLEVGEgsJXfafGs0LyTLfzb
I3EjGF3dM5BdbpG+xqiOOcHOuYRxKo2R/fZjGkrnjrsv0suVeKofSzztMs4DReCaLg8E/5+Iv9Qc
K4IwNBwTx4SGW2rlbc+d9KTW9cju1f8Faa/fNWhjdER5S1zcQwXl00YjS3XhVXIR9Ayn50kFVjjh
+K0cV0eYZZelCGdt7V/lZnoq1urQwAotouLueurewhj1BfFZ79MykFUh58ebb3Yf0D3aks4TxpRM
f66k6Gnnhw2hxWAm46KPJ2Cj/GqFYnkrbyRw4NWUZ2Y49OK2vnExJpRnK9vPe3Bq0oEifjeDXgXN
6ykrNWuG0ns400d7tp5WbOuDM+Xs4AS1wRg5T2SsjIBBL7sP/RmSpd81Iis4DbOddEI3NZamx9XF
iCzpOZtJ4xWhUTpau3OX34CL/EZvdFrK1qiLmVKRbY1lyoOdhvUyAbanQu6c/T+5uZ3qz/56IL40
KGr3tDFS6afR5+wgwLGCjkQA6rS90Qs3bsQHBQid7pTy9OWj6+sGoMDu00SBkUjISwN17WIvozSZ
jdGuJgzpwS54GSW1W6MHU3mh9yw4jexNViB+/izlcSEI7qr6Xcj5yYCwWPGBytZDEAH0zqPI2uxc
AZ9OAt9MT+mjgqZWdm4xSpfgH8MGcXuvXqz+lDF/RHZ9BSdL5PICozeFzY7DkpQZR2zSebLF8h6y
Iw24VuiNlH1Gwl9oMa2KouvKCaeQMc8kdQ+kGLqoYoAti+Ry36Vi8P9gUtnEOGed0VWO+DWJ88RI
//Ct4XxbD9kk//YLYIc8lBuDjJQRC6Q51B08jC7NuKuepRw/Db5bXgtxr/Eg0yDBLZLnGQwTXl/P
i2T2B29LXaqFlHIAOLFrGwRBrfc+8Omrul7lvNwArHRtlTsdYvbY376r7hvVvvl+ltMREVyksHS5
TO62ovXFppUl52LEODN0bznuw5TjCmF1uBbvntVioQTQC0S+VSV5sKa/YwbYzuJwdKX0Ri7jDVn8
gFxPgbyD6Lahh2MUjzWj1sAS9gRlX/HaUkwt1bdP2koH3I7uRNghE/vgANbsgAIuYFrxNqecgPDv
h27Vu9tMYXPx0l218fE9WEt282fS3mNZ69jREY6aFBagnOp3Lg0k5U9hksVMGbpNS0n/fX0+f60b
lMvRH2irB5ftK8St0ESGcoNoZ+idBz0gp7h5LJkLKHnTqKjAwR19BGxUPwb2SDBozaoUHfjzYkk4
+bjDsxiAy+WyffALL87NM8Uu/OoL7N/tNUcbaJZKlFZnNXDaC6kavRd45XLyAp5hlnT3niXtVF5p
ZIli0wROorGHA0pvc4F0JoFBBhN0xWFTbcFynn6UK3GIwYFY8gurj6gWgabxCE0QRtfeHzpswqMA
n9WbgAEzFg7dQUhNhtT/xafDueFh7LToYu1YxLVC5CK19fZo04OP+C85Xu9FZ41RWX8AyrVOMBH0
Rfgp9YykQWL9IusO3iLyJfDPktDrYmErOzCcBbeeRYp9RxGLIjtOVpCftXjNgqXxJUh9aXVyHEms
LZb7w88vH8nVVhnwOCsLJ57/39nSKTHHBYh0M9TqJbrszi6OO12GdT4khwX6mh/rmbQUJHJ5olKR
SAShDMqS0tdWViBiJph2fp/7uSA7xtA7fwALqJPFDaU8IieZLiKuQNmBTtperRvMbHm34L20Ybsr
g/pPMlLZaV6C1312INFTZgzWZKFkUKKpHabMDKD6Lo/AleVZVx6GBN4iYF0Y1sufsTWVlGLP5rQv
thKbSnWSTbhm/i+GIfAFZ6tuyo8+7v9euwg0ZRCMv92EjpkzcNrzrOBFuECarjykrDJifIZ4de5x
6RUyR7Sf0mgsVvY3FtQ7yTDh2SgLf2NHv0AS5HRmWBSOwuQTGzduCU7DCiRnc5Or1abk8uwBgImh
YbhRqR1LtzZwemf/81pu2qeZmZFs2KFQd3T2nBdls+7rsXBgPRiwD3vmV4fELRMPntDmby26eeR9
DuGkj2PQjnRUVn6nE4Jjp3pXfnp0v/xQ8VhoASI+Gv82r7UQq3aeAI9mbr6x4gz3J1n7iu6cEY4z
nNmqw9bqEknw6H1kZHnbr3IKsGu/rc9/PPKu7mKvo+FrmT3m6sSZzpPgOF1ELvdW0yfxbNm/j/Bz
j/pQyEXKwtU7r8PDxc5DYGiS3xH0+eZ00u5kknPo9+jb2eJWCksGRUSxZkxbIlN23HrgggNtUgDy
yAFfuwRQma39ke9yZE/tIgpUV3lu2eq//+uGQLGFtvt8b5BjlyLU30ZaKFeqQ08gLsDymeGE6wPX
06/H5IVe/0fisv7y6nSTifMhCr82BDyrT+9Nni7tB+9UYTT0J5eeeZrvSzRZRmiXpP2RdnUxOt6d
YrLxyg1XMQhlH5FWQZmRe/0RpkX01C9ytypN6yTDQ/an4QFQSE1ntpWlcO0ItBk9YWUmmeQVlTih
B2yGNkXozmduTxq6515Jm37KmLwPSnOfOc+BDRy7k6GE0o8gcCunR6rKLKQnxQhAVq5PZltZDbMq
UC8T4kow08+aO3PqzuhVz3mCE/JcBvUnIcm0/sf9+i1XDkL5AHLOjsejEytM7mrNQLS/cL/U5NPR
s7qWwe1d03v1lzd4UbLM/SAZn7QUwa0Zd4rvbnBlwICxFOT/W2VoTDoH7rNFAF+LNaopuQIL4XUh
TWRPBkcIqA/jVrFBL3QCwOt4Zq6+6iGHPWNM+PPG6kVvTg1holMeGK1Nl2837ndDr4hdeA4jrNth
uBj434z+jbLC7XSa4IA9mkkRixSqw8q5LiJ5ujAHVsoiS141nl2UcsAWJ/2IyIq9xKveA54IrRrx
bS6+7hTlc8M+HASVou6vliKp7BJ7YAIg+TRZaYfVrWeBEgbCtpckAxlayW0vEfFyqyIFaE5uqh4Q
Xs3Tts+bc0K6illl9eG/iQDkKI/AIFgK888FaVjYRaupMSroOFPscNc3NkOLrC1h/Bz1YkMCbJeC
qC64LpjZz4tyAB/6U5cdhX3CWbv57dMP4YAI9DS4BfT7BnsLZO5pFx5wpZN/u3OAu9fXFkmzYHVR
FA6Sz5LMQRCVClgaVCf83Z0AphNxbeVrz3t24/V4CqNoXZLOdVJa91GYsdx/i0IuIGu0HipGLlS8
4iWDXGFbyTBoFLHBX1b0qhgxWXfOAXhB6tJNY+Yqo/K/pGwueWMVYllV/FaO9lOmAaN5zXa4anMW
EjSsGxo6PuxDFLN6x0iMp0FVLgcjB0UYt2WEDxgJtKNsI5wEcVd5/pjjq1VOgoN275Z/TyFAfuCe
jFq1bnmS5Q4jWNk3aqPLaSyBS9oPJXZwgueAW6Gxw2gOFBK8X/lCmlTmDwoLB6H6m/xUy0v2DbbP
f1gLNPXXOKWdixKIKgKTbLAi5lGpwJUMg4zHsb72drlhBuiJQCMANyt3TfqCaTriZFqxPmx3H8Mf
qkswBvtWxtbgMr+1xMzLr4kSdLl57EMly+p71ZdupGbzbKZjfcpaVXn7NcG7310encw/MuIYWfA9
eWfNA7sxg88YZp7JfvsaeEkp+T7kyGbdA5va7Ze61zDz3GzPW9shXUIb8pf3gz0Ro9kFWRyVxLKK
gkqYLJdDLzN+TYaZRLAU4zohm61YovDu7jg2IUj3xLXOvkEGuzMNjgdyEuyD2MMj7k8Ejc+FMJWb
7ammKr4k4T9BhWB9sbLqc1No0kyc3SD+sZ0NpPIETDKkQbHZF21kicvPEQ2608idddzCsVAZrq9M
Msm5i4tDyBeSs9C/51UKbe+tlX+B5ArWMGxtZUHRS05t3El12UF0U0jXJl54F9rk0yMj1Fgkz+1D
SaC+5NLWj9E72bOJCngoNnCCsRS/5jZS/UuFLF3TVA+dQsvjEegaxp/Qg5ZhaP4pGWKDDLgwAbJB
GEfx0YWhbysy5/FiXIh7QUd4JiOBMakXwpiY7vqDIznRrRaMFUAW8UVUYuVMGQpXMTXS+0vQYdXe
+KgZJvfSVncMaKLQCghDwCIbcEbL9qwV7dJdEORCTJz/OV0rhD0ZBov/pOYXlRr3Re2wh/EPsgNu
iDpg9VCaEtCjfkaAHfovn21hukEAoGgRf+SI+T+ysdRbE80twLtzrwz625UOH+xulq1d9PdSgNnh
8zGp77HUsr+GruRMUyyjk7119vJ0GwsaZJNwQ6h1pDTG9d5XHpJkVtaZkyHvtrt3sF9UyOXm1HgO
2DN7C0WW37Gw35rPGaL2ZDphtt3Hb0BRT1FC5qUMVnieNlNZejcGOhCqJTnI1afRYlrDwbL0yKli
JTKYRCGPcPbtijXBVNplu/FEHWLf7feORi8ngKee9VrrqKQXAbjdm9LEeM9u2HCADVDmZWS1kLv6
X4XByOESMdZtjGyI1q5fsbs6uz4PDOPrdZ968jxvX2rWJEhjeUw8QGNh2UDsCzStTJXlPp5Ghn7b
EVmxJ8YXz8tfHwpoc4jmxkPupKAcydB97aaKBVcQORgwG4s2kqLOHkY57bCbJbjf2mXbbiH7ExhS
EX0vS1wH+Ot589AUgQBmNEFjOnOElQgM6EpggZESanHqXbsLI0BIfjkNtbKgu+lGmmRFjeMoxQAJ
XK9O9Kjocnhdl3XRptFDI6yiWESTbNTZM8SNyPTokP3cV5HYDu7NupKK3BuJA93GeegUk76fbAHF
yD7D1YTfiJppPMxHrk6Lhc01uUdeUO+XsGgLEJMC29DQnXKVYerpDBguBVQrvf6P8ihIbjXjb+8J
Na8FawTq8UWHKJcGAUvTueFf/eDx909ZRYXbTW+CpIuKMwjiW58dzHXF65LMvKogojKOuDuEaZwP
EA+Eo7QzEh+Ob2DQ0YZYJcW+maRL0fWpO9zIoUWqpjAZfx43P5BfCzLgeh1PASNWPer+5CCEwsoB
H3uinwloJfbYQSEMB4/Nei6JN4JfqnuF45wh3hE94mDlOo2ndbFjhevA9GbuviPbuhWyI/OwbEBq
9O7Sd9heIetuRTDCeYKVx+WWPMiN4nrwBaY/TuaCpe4+JsqEXzEPHTdS6oD8KMDa9kP5UH5/stXW
mXYE+4tE3x/IoSgMM3W10qiMfMDoEZSyePRPewRUUIVp7+BObJiUEllGEqn8nlMrLjYaNGAEFcPf
/hNf0vnhweBLcXTnkfzjYNS9haKJOLo1P2fz9FZimiCgRubzG65bWniGcvbLcJNb1dcDAO8Zh1m1
6voaBreHpx4ockva5vtvfEG6vvOERFm2MyV/ue+5pWnDsMTGQrGyv/SM5dxikFfrOo8bj+TRVBJ4
InGVR281imwNmM0V8oFnHsLW9vyCuz5XlQPz/09/KeniZIx0+0zQS3QBSS7V0waGLm3aKMADZJlk
FJBAetqiuI4Avnb+HCZdlxUnhBm3IfItj11Z9HtUr5TzokjYGM8/rAKa7S0w16hr9dk8pPca0gt8
1ftOAb7i8cNPgKh8M76ijJ6pVMyoW8GDglJMv8zEFcDORexXpHChohf78oQpA5Y3qW5xgOzOBU00
MK2rd8MCPgAeggABiM70CIcyU+avuofBUgntF6fNmhFvRW4lniN/K/rok3SP65b6hdm6YvCXRdzg
dR79RUcjvPMqmlwT3PVTKD9/f43i8grgqlpjb//OKhVG6cXiYqa7b9HbUEuX8Wx+YH2r3TuDapVp
NtimIaVp3Zss7qmg3M+4S0lHERIZ563lFVZb05qP2CSakG4MBpYGkA7BZFWUlkTmi1UwOh2ShbmU
3cqjWFF2eVw8gbsrrAlvCIa3sQu2B8LbmYRebsK096PMh7g0CIiCPAChUBUR4oI5/V/O+TIYuzVj
OP4fAzx1wlDuGGkonzNhW3EHscVXn48ZmCNZYKZxfWnc+tzJMBzBRqsCBuxHSrUsgX9lexYTek1q
7JAV8NXeLzN+xTxF2uws1l+vIXo88Y50TQTdB2nN4tY/cqCdB9ac9IKm0m037kmifzC5CerIkWEA
wzEw2VNixkLT+OpZwykoWq5FFuEccpZKRHMBgrA4qXGUbozC1RaLrdubWztc0yA4D3WG6BhOYJif
xpjeS56geahyaALA1BLmXcNuTLl8UkMB/n4tESTmv/Ia4u3q3pggTAQz5m4pUfYdeGPQlhcm4ozK
PthRyBpbZJutDd3+AGZTl3abkPsUdF2xGH71U/Oc1oalK9Zb7oyYvpW0f6bqucqcPJ9odITUEigq
pSB1dyM++Ma08LLuw9IO54rwHtqYMBaSF+0ZElj/bhnN6Nu534wI7XxqKw5GgV6U7LXqxSDzo8q7
mSJx0EynjYjkF+3njGxatVeIvysAyUPDN87UMsn9c4RSeD2KSE5kMoRpkuzvqST1uQpcDrLOOtba
/PDauIC5ELigq40Q7dSe6shxULniYTfqfarQRVzMMVjYBk0UHdSt7uAX3vPfIKok3h8qNONVaevx
0lxBeT/VKlQrHazpyqAkKbWJD415UumtsYTwNUf6Ec38mL/PBZ9GvWyUglIhLsp4Q03vVQ82FWT4
B592xrmzWMZLgk6wJw39s74HvzHxx+LFrrcKOPG3x091yp3Z5PYdzexnkGRlqIf9Q3ctVIPVUfQp
BHMvOp3zsBhDWGlZ2h6rNQBDV+W6VdK5JnPFGTMOcI8uFi9j478wJZYWVl21adqPVJBonkOyZKj8
K1rn420LBju6tAM2rtTVKX2RmMTNEzLGHDZ5+qF/m5818iCvHA4xEfJb6tpKZEywrLLxnue7n8fU
efefvCrKrdEw/3iXLk6NER7jNPEPcpLGJYHI0WY7FkLbPO0W2gx8h75opyDjLP803EIJ4oFPxtXH
IQYPGwoOjhXT4Y9OstNMUzendOrFSgleC7aETuQpzQg788Ay4WV38pm1fBZAjFZGZYSiliM5t9wn
wQT0FHAqoNYcoKDZ0gF7uYHPjO8pAMaSmFeCDKsc2pOaKJWty6DvMvf7ts8Zhxw8xyRYYBuquCJy
O6zdvHBShS4qHobCagIHr0yq4BTJRef2FTdwU8Mw2kOb9MBFjScUhlwsz+Bcvfom5CwFG8c5DPMy
EAwxOgxCXx6ElVqCWZd0dGXPCSKmGoVwUUsmGCanMjFuPlnDSwShf5ltLny370PqlzueuIMeTSVj
rVuKZb7MFHoXsf/q96tiDe9I737MHLOHWHVGf2CU1fa3YNvL63rCxeTbURUHDg4vZhZwKcrbHZ0D
OZvj4u8/Pkn5qHV+vmBdJpsz5sSfMyl/JuM00EmBicw+hCVtRl2CYI7+Eq55DJgXuWXyozsI6sZs
s3e5MFhqiTErPfHmZkI7LbFW0hlJuNV/fNIxxqWRMca7gQpMUXHSGT1+RLAVoVX75zrw7Peltr7P
Lj5O9f8TsOM/nhoX8AOTIKc3B9vnN8mu6DEzSWZIdtIfr1V6beNHPCztMQS59NbPoIGCfq/aEaJN
aCgcWM335bOoqKFbXGqZB/+4EnwNdaBfaz3onPf+ZuxG9uIcMKClRnbcDFcRlTTtRrdyXxARTSDT
7EsQOoN0wsWvCG+4cbpwJpd7/zGxHZPm9vqyj9T03BhzSBO0+PXMBxJamM2+0/wnusEkcbMvvMsS
AayDrO4xTE59qY7hl9xREpj3SPXChCnkROF3jv0SO/uLds24knPNob4FWsxhiRjLqce2hFmLraOk
x55gEEeooRej1f9ZKq1Lx4xIlnAaEtUBHIwwqa1o6p2bY9kxEYza4B9i7fa7XbeZxKwnegRY1jS3
KseItfH2JXN3FoJ8ELcOP0IqaNqoUZFzGq6/OTZ4Dnrs2LVrkxaNdRkmmTbyn5Wkj01meylack7t
+Zo4xtsaeig5q/G/z3Z7m0QUIiU02xYr4vY/sAF13YmO/QdA6Poy+GgpeKhzydoh7RZFdisVKfyw
pSHs4yiW1dL6ACyY33cEkBKAgCwePaLHarb4ucMy8URqtQCeWNlfiKB5Y4GZfBEbh9bFmLw2cU/J
FvtA7a0r2ua074j/rMeBCqe1aUd1khoEIVvX0sXLxYE0VZFx2ZFGVNTzSCTYosPIr1ma3MR+0fA0
E+xN43exgFqWKb2TPgoktBLd/JVAxI3Z4bHQqpuEUlLK9L4FmprXJ+9b+4DwLy/kJI5eELwzZYRb
L+ioMqgGPfmpB/SJvCXD24ely06BvuJaJMEYNm0XE+PlQCcslJl9OY4TbXz6QCjySsNWbk4zXhHU
gNACWHOQJU59TJ4rWXzV14A+a1jt7C3PYh5H04Bx1kUVLKOO2xsuOzXb9qQj6LdkBKHrVtEHa4qr
nav7cLMaFa9OY+a/pOe56cBSnnF3dYgLkkScFISNxfhCxCiNiA/QhaGOjyIqjoeG9SI+CWGsbLs4
/BNon7HO00qAk76nbstRp1xksFG+Vjx26U5T7jerLFz3tReK8/9zyORhqlKS1R9fYcaeCGekSfk6
L9eFHOGvgLU2DCv03zeDNylCpUQqYK+1qUGgK5kx9kerHXuqONBlz6mHqzG0exBD1v+46L+aVM1y
PakS9+IUivMdqJBSkkCyA18CDHAsP8WHpLjt//OfIMC38uFxbfgpx3G42SgwXfMZZVR/3tpWbq2V
B0eQXAaEkkrM2BsYJ0P161aBCZTOyEUCykfuYjYoj3Zdqe25YmdPHaI0S8Qx4Jw+a6eCezwcP28l
Lsxi7OLqEzikSZE5CI6A9Vz81Nsk7fMpj1kBjZxH7+5wJxO7qtKs77d5q2+S51AzAAa3PsTDV2Hf
QaskYLHYPSs6sBlSAHeV+LkcX9xzSGGh+7QyKK6PEPKsarGI8EHFLGQln+hVM0FlCLiXfWEm7qib
0LZ89xxqjvbtApC1MWkxHiFm2Oydhm+ULilD/p00+Lj74gYZOQDLXarDpu13Vnc/BplzTE3i3VFY
Obu7pwk9JyhxkkBo7toY6P9I/iDc9W1kDuwCm6LqGYP4ZeaVm+T2PnwDLres4yZHoYuEeX1SN4/n
p3fNc08tJPevHGMUfOx4g4bXNIU1m7WQhwGhB+EANWR/5MgCmozciuDrGojPpGU+YvXD8mod8mOl
rrWUQ1M2ZmvRNJv005TcjJcIkQPP31qW1Ph2NVw9xuVCHRIJyp75t019sgV4Jn7qX7cAm+BOYgBb
kSTTPLvEc6tvODuoMuc+mYagLy1n07WvFGpVFiJL5KQbt8y5jmCsbfF99pgXvcJYau+Sw8GJEaU9
MokpTDBC4P2nvffYXr+swnUi4djj0F6dOrOYV4vD7mwYn3RWRutZ5Dl+rweuGqbPnchOF3s3BZnH
Dioz+s3J19uUj+FHRzIQGgGBHj4RrWM0fwnw8jbnEcxCU5quaApPJBv/kC3rAg8ETTESXp3gBpuo
brhydJTPFPIpIL3ajim49gMlQZ0pQbMJ3PXB9lKHd3aJEzwxnos54AQSNIdofu/XRPg5BEUl/mow
W1kmuLbu6lP1ufssvCG5EY/yrXMrY5oC5M9ze8iB+Rb9blzxSS5/E1WfwJQhwtYJF/z/lOEPB5+X
c+Ewx2YcltirkImCQQB1L28kp9XJwBjMWzJVBXiYDpXpv8a3PUJtI4vlZBWTyFiG8+sTz2/qa20W
ETRZmJLRWCdidC9zB0oWu5PX9FgyHxbc70hprvcS2sZxg518YLebULwDA0tMXv3FTnvSjaP5OxrS
MiGGyrdwYQvya4YB9fEMnmPjcVmYD+MODRZKGebv1bEurvAdL7Wn/hm5DV+iymTj+OLdlb1WVOuY
ee9uglgVwOSLAdNYzo3xNv1ixGEiO2V4m50tniVNKY5TsENicUYPdqSpQsHQ+9wFksHRlgdlInQU
UPqliYqTB9uZg3oVoqIfIoDR78MpvBh9KwcQwsNAQdjbi3sC1zhmMkBylOIDq8MIm6k3TtLrssmB
fgvqiLoXllB4ibW6yCf9khC1dxDbO9xPflyo7cEpVXS8LiOgm+4aQGPJFff6x6jak5Qr21svNNyg
8zkag1QSqS2zFZfE4C2o54uQX3s13Nl6sjZmubnxySSBKhnu/KBySRUi20kJScKnFyr5Se3tX+B8
Z9ZTaUgbgEsnVMuczXj2boGhSfuvqECUB1L3d8+I/t4Vnw54omRzfEqacca49Wpyns0Qq84cfYy4
NWo9RRy3wQZ2o9xzQXz+y80qN2dNanWuPBv+q6873KwXbXgkO5tR0MyJ+k3ohb+tIzkt09qnyLJm
caFP8oMSAzfSeUQZc//iS49D+KBwoZ+HiMV0ZXGh4s4zZzJCZWPFDvyZnkjJmTt+M1x+we8K1RpA
lIwVH11EUbV5JgEg8w8MHKA5v76qlKtASGc4zCVuMsf1169uTEUCKfvR4iGKVsi6QVc5BEzwbHyx
O3VetC7DpqL6bCkI2qxLlvas0E8FS2H12lHf4exFUe4f+/Z7FfNjfGGVYx+Y6jl9SMp4KKFI6HiA
JzQvuaRqDr8CEMXForVLPRpgJsBvvb0A1iyaETdSRpxH6X7bx5WAWZ7LUUo2X9eRt4wdx9IUN9B8
Wy3qzugX3zWl4G1YiSnRtzTBHXWKB0az5u65g2pUaQ6IQ4BFq5aZFbtusXOcNd10HRmQNAaC1lo7
GPLjvnjgnrMhPh86TAoxmOaEXF+RIVT7HpOI6lx5j/BAgeP2ehINpca/Q9k/2boMhC/rCVIrApju
tnqpe+U+fSGwPk9ypwliUAMJgcxWUvF0JgY5C0YzfzXmbH63i9vk+g8vFhi3gHtz4zLB0/Z8x31z
P3H8GwiJE7Re49xme+YOJrmWCEhw2xMPocdnWfUtzkuQnkvZ25dziWfQSDwwv+XFVmHPkLO/5w/O
iyd0I5kBHZX2VKU5B76EFG8z9soU1gTRWZUxtEUg746qDElOji4h9PxkkpFG7/QqaRcjxYFOAxr/
O/tIaCT0KvCx2Ul7oMh4IjJgJaZYKddfGfI2764TqSJOkt1RYwGlWvzGuJTj1KlBjZ9kmJibAwDD
OXDHN+p1Xf61Lrl89DEiV+UTxwxbXF4eSX2sFtFZeLUWwfcks/a3CfkY9Nc2sBQx0CCDkx81+amN
uYJrfPMQ1Ir+IGDA1glvVhiA4LL3SyfnzjF1TdrWz0YlX3qg9woaHyiWugP/93BCWU2G437xCEV/
NLwK/XUU8f8WvVv8LYJCPKx/lx1W4p8rlywBjN3rEXMGpQV2nGmqaZVgKr1drsmI5jZGdJbGsbc+
cgPtpm2ovI37WKvtEp2U6+CcysdwNJJav55nwrRlQPbQwhDooxUYhmBfgmmFTtqHkaKbquWAK5te
pBNuoetT7qhePbPec8XHH6wqNjdPJT1+Qg/4o0OuuZY5nx2bCM2YLoBNfycs/QX8+VhAeFOm5tr5
l4Yoh02XpVBk8F36qleOnwlACE4CLJMTgNhfCt3V55HzGAea9T+JbiOYjXQ/oe5WDew4Qtb+Ml70
v2eg37Hm+iRad9pVStq6+IOCcpf5/6oIH92SxstVQDZY6mLtrMJKZ3fFhTXyZCNQAx6wpd6lmGON
3UOsWS9Sgn1Yu7bvymRkO4mbLvTZbLjgxsVDeXyICZrxsoW/i0p/LGms5meNQGjgofxoqUTkrpwv
hZgA1w15YYYk9TsyZr5U/qqTkPS7Q4Zj9yXgIvMY9vejMYebA2ox0psvTATSkOha/jTyP8CkP8u2
WCfxBs6yC+YCjfrzojRzyXYFUZeoi8xnIYNwaq51mAhMA2xSIQpI8QZjx5pU8zj2ybY9c+ns1zDH
swY/6FU7T3jVirtFvrWCUr1WAZsV76Pd2Ufn1cwtFjVpza631rblJgC34d1Fw6AAxMMWlx9YXQxO
GghZI1nIQPobCXdWcJbr6TqtP+gJZkfIkaDha1g3/Y74yDrB4d+QILVcKX/wQ2yLdgHs8J3LCic5
ehcPSIzSv2ayTrTowOYqYHhi8xT3WRN7FpMoC1ed78e8RGwd66lo1QzwoZKTnu25DLgAutc6mJh4
W+yLDFtoneA3PYee6AKnhtvf20uzxQ9LF7ibZa1+e5PJWC5pX3bZXENnP/rn6S3ottk7v2zd2NGr
7OBjNYp+TMvIAZmhT4kty0GgQ1DY/HGUI6ufFsXFmM9GMyWURK03HaUV/Q6o6oxkkQB1X8+qIsfX
UJBs55fMRMZfGcb1YKm2hnDiR+cp6xUn31J9wBqUAidd/UAhjeXAE3yUDJWep7qCJpI1A2JZCe7s
84rlygl/79TONzD82QHiy39jqsRQlwQNvYFWxuEoTnvt0e91alMTtxld1dDkt8jfZeOc4sp3LSqJ
FEj3KiTOs2pMCQjgNUX8NP1TcDrsf9mBtrxjSKLfnKRnGj9L3PFo3CM9KpwPhyJAv20otZShRZjN
0WUhpuU+AUXo6nvkqC+kNtFHo94JOmVE/Nkt9G/n9VRubu8UePebCGnZ9J+1fg/xQygs3xXAXXet
q87KdTdBuBkWdBaabZ6G+Fh5Vyy0ejaTC2T6RabM8lhWEgXVVT6/c/+PopDt9UX6LY7knByNlPft
3AABPlYykz04zW7yMU9YUyfz389QYKICOm7CgvhYbzm4a6IoQkZVe1VKoYIi8uPA3R0uMVKRuNs/
TGRIrMmelTUytDJPja2ljdRg3fxqgJ0ugluWz+egI+AzlWS0lFXbCdaeYfZrkO4U1dqBSBsb++hT
Xtc1gag8/mjABtLiQ9FnGrxMUZUnpC+UE4nPqc8oZb6Fp2QvLTPbcpZwOJNWawgoYSKsr9dbJy0q
sA2lNKi4Q6X0hw3r9BT+D3Tia6QNuoRrU18ryqHzTSl75JnCPpyWakM15vWI7y+elFyOl5dyZTQV
iJj6E44wZQaem8JPsxrzUKDPwXBxy9/OBzAC7Z4MciyA6rpjDCOZ8VkH3MZxntzDxI9VjBB+9UNd
YXuOCmuAfcPSDS7YEAPUrzdLKcCv0Cbx2KCwCA4ncxbAaNYAjHQoIwIl3KVG0f7t6yTVURBhDZez
9F/nqAdtM1SHQpQPqQcu0tYbbgzfgpC2qJCJ6IVA59w/ouVJApOwzryV+2lwEnE/iugM24+80xtI
9zznqSLrAPAT8rJAKeXPTwntUCtlJ8gw8ym4bDxT+Cxu62+v1r56NhWnRwlrpkiUs/xnMDNvYGM0
FErap8wwOy6J3+Kcev43JswkqnNTL305S5qAjM58X51D4biJytldTv3tLqGx5F8NESNL/DHAEiJa
fUAj/y7/Y8KfOTAYor/ZmBNpe0ICxfDp8c/0DAN/IYm0eECAmqf6b4RlDI+1bU8hRvdIPykTE1Tl
tAY0+KRIRVbZJvtTHahtX06uS/R3FSRYE9X0J68r42EVmYK5hlseUXdJ/Cb/HzwlepHod9V/ol5u
PUH5+26x5iJ1I6r2+S2Ehce1VqkrONv03wbi+sDN08sX8hzFCjyAMH4menbSbW6IrIpKY3wi3UQt
6faGqkYjo86wxP34/YUQBdHPmWl1gZnOMrVJYnNSs930YE/FS7ClZBvyRI5GcNHw1m/r6gxp8SzA
yJmnRwiH0qzKaRkAbchfL4w3cE+CgtvkAPrBnA+I7TM+jym6XNqcj4aG2Cqr2y1AonFw63Uwxd0W
H0q3pTwRUUmLvr8PHvvy+E4jpe4SixkqOFBd2erruOzppJbialQhYzp/i2XSdkTzUcyGpgLz6p8Z
p6HLWHjo5Px8smVgqrGsmOZXBPDeUDR8M0AApbMS6ahUXppRfQxXkeORj+7dK6PUpl7lLHPG+kzQ
eXdd7quXpZxuU2DD2aBaKVbFAcBN4Fs9PSMFwwxO4pMvcpnVVU+31B+e4AxNFVY8Glwru0X59pMi
+CMEYdhrKHGHK5TEKM07rvtTnb8Au3seidY3yNSSu+A/wEYavmmp9ZzrZUQqX50Jwl/NrBf8HT3a
/2SXKdSwfl3NEWKDFhKV/k44bp6i3fx6uUd1twtmzZlDjeydGJZienQGS73QKGZ9nR2W16td3iEP
TYZHvBZxpTJZWb8A1Jjr9hKl/BeTH+k1ubgaipHW7M7EdjvswaslOEZS8e+vCUVy1PP/zu9O4RDm
cSjbI5ODfBNtUMkjRk8LAtZHZC9zXHPtiqyLjiVy/cNrlTwfbHFSJbQZ87vM0RD2Zo8+WJoDSLCp
OZ5xMIMTPfHym2HrM5QgwXMlw/BSoxK/CDXVa5j3RfTsot5Cm7Zw5+ZIT03YI8PM2wfAB/XM9l/+
6cEhovmqwR0keFOXaqPs+/0FMpYPm4o60EI//iFim65osMy3U/F+nt0X3HWlodnrkGY8wi0dPWvy
i0MqboTScB1K2HRohtbBEO1hvXwsWF2Ix0XEi74oxxU+3t/4w9wDbE1R8tuSMcAW1pvgoGpjTkvQ
Zc89DqNI5Z9o+jtFWrYzn7p0pNKAxzN1+cQPicfSKV9EH07Ac81q5ery7yWQazEgt6NAjh9CBzQv
3zVl6uXtk73NnaJPkstEd7y18sMNkDh2c8Nij67iST1ElXVl+rQY7qknMv6EAxyzbPA2ME/Baloh
txGS/6Lem0K+I27206oQAeDmwTiIFe7/91S8Pt1YHJ8vZ2OVGuxeydLHf48gOlScdnbegUVPJSK4
ZoERbqHs2gsgHVbV9AKzhD+8bYYhpKwV6v4rDwSJVu7M0obyffmjbIZrvTaYalLG68tJN0zWlV26
1qTbaESeblBSpP1j0KKBPT7TNpG3XPADTxsNHQk5Z6oQLdbFZTiNq/7/Elo8aIcruTpnDfoRwTJY
Z95ElcSDOMSlua96cj5oxhzgPtDf/VwbVPV4vkhEXGr/6oE9Mv2CUjyb1SPIrAuI9sbU0iTSn9uQ
KgNRvdnovwfs6+FtVbR+1fbBN3n54ovNqfkOf2w4KNyWhh8nNGye3oZuewoO6+csiKTu4jqJsmju
h6SNHNIvuVRH3l9+8tp6RUQGxENt7HBS6An7d5smQWUKGUQDQ0zWtxOhJZsuG9Qd+h6Lv4hOLShw
JYMibP0+UUs+6PG/DSfpbqZ4Gy5/FzfAlj450F0pLy+WAha6IH6BQZJ0D1+XLHjbEq9myoULcP9f
n9UIyXf8WOdnVd6QoOSMCisKmkrGakZJUo0nBH2DqhMPseDyALxmxMjLjToZ3zuYZaydPvEkFG29
QtTzLs3eoF/zYusaU5Pgep8fKtzbQ/4g2yV+3zDpJT9o22W8R021xw2jdW09Ubb9s77k6ChKwm5w
aafq5CDSTFHJketMvx9HFzB7NkGZAeFho9WzKj+EP0qNGaqFjPOTuVJL9VhiXz2q1ToHrYn8w5FG
mUzt6APCFXulx6x1KkKxYj8nYVnFaXxEB9YFynVeMdGHaK8h/wcgUgI7uUA8Nb+t1D4vgHY1Wp/N
mzAIkJWzkOr5qV87bK3rFnz0WCGspx+HcQwwibimkY/xSp4lfjZ8e6nWQxLNF8YL7bWFw69ov/hp
0C8Un7LKZfbq2jPTovO2rQHv3VDuFYE6IaFFj2ZWe13YFxL28E6Bhq3EycZd3OnHdlgeqOzz5w2e
EcZ9hMnfZAR0iu4yYMmfqL8iScMTseSDcjEd7Ge17ztlkdMjnV2RZuLUoJWnbx5XHMo5/ebRZ6GC
vanZV0nki03v7azE2vmHh7A+KbnxIxpWByy30DUJQkzTgILmiL4BiHGmQ6EegoaI+6r7jmp/+23Z
rnRLd0jJVNKveey7bz9zj+mhf7gTMTP6jYkqXhlcG1YJvcQB/yvsBkGwUbtDzDfFWPBCm9rb5u0j
NnoxjxAgZY+4e02sw/hszH6pLHKcAH4iYWEBUyXUZrQtSXUtadU2tukA+uATgVseADHznFoayH5j
vmyMjzf17tDqkg4U5P+Tw8bJ3Y3RNwjRUfZ0k0c5iC0rGU/MTMRkmWt6QA470dirmGLdgbyrMAVf
vzoDBto/SMHVQUzkz6ggc0lfqMV/P9yxDTPEk+Dee1iyQPfhoc4ZlWPXS5DdZaw6/OL9FDauVavI
NIhMFIwM7/W8xVEBEqeOP4QTWWU6jpmqi0bTZbrE9js8dM1RDTeiQW8gzbKNbPgUucQy8uKqaIHO
L04a+cNkj3pMmYGulK67s5uXu5qXkSyIy3et/xcfabAOLNahim0k7r9Om5PCbm8DrbP9W/SX3L1X
OvT+75BLZT4EFFoDFn1s7VZMdmzaXjTt5kSAYMoKsWFPEfxOUCA3wyJFjlUkjQRrGtqD38aBfMnk
3QXZLW5F5AFw1Eag0RSoPTojGUvlHaGHV47c/c2D616kM0bYtamcuQEo0BIkVb1PJXhCerxLAPxn
6ZeLMZkRak/ejOXQwWXDgIPQzs7SptyUt1wXNRYJyxJ0CtnQH9RAll1bXgOQtWZEp7o+stlaXPQp
nIB3mhcNvfZMCaEYXyMXIaI/E5RUufzcJrZ0aasskW9Dv5dc1KqdAYA1tHk6Cym3s3GDVND5kloX
5PmgSa5UyYB4mgjvypB+g5MqdBJ8fA/WNIEpd1lRw8o0fPahXB+0cbLyjroKL4WQBJbBDeWDES69
rKBQrz3txCUMCXEdHAo6lGG3dMqLJcqk5wyL/jton6czYQsUlMpSi2Jlnczs+of6lrLOyQgrOXrf
rusi0g80A1GP2zjiaS1xwvhZjvu6OkHVy4OWOQwotiANaU+zL96ONacZqtmLorBt5qfXSjW5PyBR
ILxZ6iW6eOt29ZgrVj1w4vT7cgck2NFmG8y8oXXUKf0xtOeOtGSduG45LtwkCQWOGK9LIr1bH3tE
H3ieNbdTn0tBbVm2vdPneHZFytS9wVAxDzUNl4/Y/nH+T8LEe4WJYcmbgpqNIuMCXLAh+LvDP/Gs
wyMO3ZTVMX/D35s/XtclaR883WnIbrflKlh6B2ySIqjM54/534+xYxboQkMq6SoKelc6ahHtc8oC
9JpS4wngmzSmFXEyj6njufCnbEqdXuAQE1SL05Y5Kwl4W10Uzc5EBDJ0+fXecB0HxRF5jGahuLeJ
GucG+L7btrBgS6Or09mvs6FBAYn7Ofmdr7EAerB5MrIi3NUXX9n6Ump5ayv9C1scnHARa2Gey2bu
rD4fOyvkSfFr77ZvLmVDCgyDNB9ITqn+HKRHQqCZh4ymm9ctMxkWO32EszVKbdS7hDGIiRuerlNK
S/D/ojFIJQDdxnzOqy7DVgos5fJqRE+mNSl7I8U+kC5pCWrqEbzZ2XfQFGuxyzYsBE2h9iH++vZG
uspb2qy7unoVqcYbe8nAQa3UZRuOdOqAbVYwlAYV/iAVlY6PJi6YktGIEhiacLh44trCX1lLlCiJ
OFFkdQr0maEvf2R9mb8f22d3N2HxknMW65ofq2tUgX8eyM8b1ZIwvBYpQe7kdo2LrMR9PgEoKIEC
ydafIF8vzuk8UVPFuI/ycQqTTuz/FMZKlD87djHLOAaK2vA4MkMWxrvMRJrEeRHZKZraE6fDaZha
PPnrqrwE2bzMmgwybCB6MXk9mv+oPfbRuRg2eBjo04mtUpTaqt0URR45ddk2+z/tUS3Ng/YfdrDy
TNkYLxXPYkaV8+/TJww5ixNY8gRElR2MXDmL1m/snfE2pzFtkb+VdQsreUNszjyik1mI5BQDH5lz
9fZAT4SaKT92qveZu9xWpVYubNMALRik0J8qb2TiQBvlIe2HCsqqBhttdR3ifNrbxDToDUKo943r
ikUBWcxlfa+iJyHMaV8JY7nxT+WKL05BySnBrc4JsbptcmJC9QCnz4WZpBWo3T5/0Pv5yc1PBbQq
UGC5WvCtCjlTJersVTnCObwLf4o4UsE6nXRo8FJNcj/qUDGpNxFjlTCHyPpDaVgHLKJcL3bzGigx
GTDIQZFAe72RLWYSbKQNTlbzDkH7Dvcx2QQDFYk2L3Fw/yjaeUuL1jJ0dYnSSCECqh5gHqEIZlMa
3I9R4g+X16yaf2GnbUyloVms6aGSftNS9YncpY+lRdvvW3t9Yq42l/hSLNksXqGflm9E1SYjrlHz
bRm+CiMqbkZLk2iaYB21oBoMQFFzj3cAg9Z7oDwglbOckEOri97jMQMQ8quBNrykl4d+XGojjUQm
PS8U/sdSp9Dx2dqdTIaWA03m3AGZ9SlUOQLqOAERTrmHzH7bK2oBfbtaEZqJ4+zSkvdNTHHYc+3O
2Sco85mwlAjv9f2Y0EgRY0xu7v7tjdHd4KujSThEanhMQppymB7/CNnmu56WzKNvnqS29lE/GTqN
9oKoYdXclue4A+gn2MstrJOEyXL3sFb39EDg6EHQEQPwvKTTBZWE+NHIhkwqSD3rIbxNErENY4rk
2js/WGaW47Kd8BQFELj1xeqcll1ZRIXvN9R5YkEhgYoZsz2vEZwlXep0NB1jsEfWUu2WkWATJ5jq
vD04R9CcrzZBQT5aPKEZbxztdkV0/cy4xWKklzTL39GQpjDgdSNxQ8fzQX5+uKoqqLWbzy/ZLRyg
fo0Incy+1+1s03BUUA9mwpJVkUidN+sFBAGCKT55dJvK2ygpV6zGqBrg1XX92SQJ3F1a0CgzEPNk
aUiBLsd8AtcLIdJIfP+xi6eda8h01ThP38GVLhFiz4PD0wdksYTHkC3Sgu/6WakM8DibhkTo6pT9
FzHORJ4ssYo5U8a38fghUe95EapMocdR3eVM6L3SKj6sAUfmdMdjlBMXSdVBzjnTC7leZQjBH0Pp
/IOCKtUvZFD3G2tpjIWxvY87bcfOPbN9V+PXUDXGad624Oi/GB2P1RS2zdM5gSlDHfFTliW706NB
LRl1Rf8NiWlQfKLRGk9lpFvYaADyXwv1Bh6JE2BaGdApjvumxm5tzX2UwzQGsgcOTm9C/Lm1Jxz0
kGILiFpNP67a/oKpnZbGWvSUfSQ6bvRBNEjk8TnBst3+JiyTYWAhdAVAXRCIMXJm7Cj69alrESw/
W4COygeG/YMOr3NxbnvPbt49s8slXpqOo0bGQir8SIPdtVngOwCKaxsr2KkUvfH9DZ/VKKrk4b65
WRYbqM8wMUMlTc+ePEstLgeMahE1XyMlNmh5VO22N9EeY66T1Ks+3AtdDhdONWM2Dw32ZG+MrdVw
bY+GwkBBRmMWto/MTDS1XdONsylgZPbkKqQCTlo/axtN2yINEr4KgNESHN4hQCpl2rxpXuw8M8BY
tY6J+M6yW9M7YojYWs2UMtQGUUmg9ghbcdHx6Tg3x/3Q87rzlEs3G6IGbTnUoUZvNeIFmbDdPc/+
i+BzhrrgimUYiJQMNPeBxqa8Ay20J6GIHSXdCS0NG7BTx2Gm5xIGrHWI0FkLfGyHgWTjkJ7EqkjA
eH1AK6Ejzj3l3nE9kW/Q+/iFfUaVtmPJO5Mh66msMytD3WwUHAmVnM6GKjN7YAZL8PS3dQTn3ZPl
DihggTke5oCLiovtDK1fTSBt8q9VGQGdvIfnjfhvKmRvQjIcpRSH7jx9w0DuD9/Ttzcu308ofzUz
i+68ThRdlzVhSyeuYf+s8oNmn66UBIS8nFNRZAsQ9HxNfpqNrYBj2t5MefIac9Qli9zL2P3ywiuh
cwh5RBf/4zCz+GvfJXuMh89lfUwmVIyScdjdECCut3KnP6F90CoW93XtaGOTIHD+Jqw3Nk5+1SUo
bMo/X3uz4dpyg/Zbbfiuwyl1qGjGw3duM7fZ/+XJmQkk2NxjSFhN6ezNzdeAiF7eitoYap4q7qNo
pCDKQQj6/qwvsrS1xXBq157ihzeF56X0jCoXO8I3DPziAcvmFUAV3UFavfMOH1nb7QdRS62i3uDY
hZE42ihQuxGJhl10NoxXGUhUl8m3dGuxLWfeJyegURdjN1pQCAuHRe5zBRcwEKIIkYpnrdr9PeMv
UzzxEuPw5wpx0DesAqiLGvMYWTxnfB0uVAYm4vsbKQiHtXZtYbsJ1GjprmO8tdDsGeb1YUiQWTZ0
CAryeE+W2lvDFiMx7XD/qmx14pcQeviHVHZ26vyMkOv48fW4DHHtgc1yFMhBttHVsDbDivWnkAV7
liwAkqLdzuEsDIG/adKYvyjVZPP64pKJEcmY8AvAGRfvBlCIU5Phcu7eQmAneEwXI6yoQ3o63sjs
rvVVPSk55wAhBx4zJ/2rQk6PCz1D7bh6oVjRWAVn+Zw3ZVRw2IZ5DEZweGBQZl/3cGtlOx0mZmJh
K6eHZGJZ0D0ddbNcl8DI602l3y4+w5F7UNb6doREXDAQp0DMxkWCttB3xC8AqNUxbmktqbX3Rnsh
fIEYTxRKceriSauwr61GVgML74VU2JPk4POim0frN+3v0Diu6bweQUPj4JPKSqNa+cjtGuiyTo2U
iB0fzBhJAsuZvyuuih0W+REGywJGqDjkvh/+/+7Z9y5lyAelPe/ogoN7ktbXB/WAjmwPAMnzLlbJ
RknJPnpevAamTcib8PtqUABvLhrFW2gaz1dJyATIGje+EhqCglpFU2M03kUzFv+g5VAN8F4J8wJm
zhMn0rKXyb77t+AcE2Ra+yUbv3vIxD+s/EzurpeA7wmBjR9zqF7HMEkkBElQXpjKTNIHzMcMmGXY
WD0C7qf5e7tOj+XZwwxVz654sd3gFOy0a9uDxZFwwz3XfV02qUFyZ7gnRf0Vu9onttjanHr5eVdX
7eTfVMSKSEq8RD2l++f+vM68VxHCfg6eKjhR4u2kU9wLgGSIPBM7os5gB6BsZNqFlprD/+1VYyXC
jP72FyWdH+VaYjDKwBo0tCKotCl0Cp7PABylZybqIjXB5xzshS6ltzG+FqaXUfcTeXOgFdWNFI0m
rz7X6UQ/xmL0/yHMUETcdCgBxxLPubwcbtkMvpE4VKS0vEWPPwn+A5CH//IeX60KieA5tCoYg/Vy
dgPsa/EM3iclfcPsGmB4JKIRr546GTjAY7ZRHmBiEBdOqkFstbkEVbVN/bCjnntlnr6OIZixgNWE
c37V6bzaaymtDxF4tT71xximENSLPpn9qEHTbUX5lQAW3IWw30QMcK5aw9Z4VvrqejXgtzD0rbxK
XV5M6BO8peImDEQmUvt2j2I0zAYkdOkaedTsc4mRYuZqeVcvR7hZHR3B98PQHu4m9SPu3JROr7mN
mjuCK4jGY+kZxrvHRrlTHrOa6grH6NVj7ojvk4Xa0R2EY4Q7rWu/k3ixfPmbvlkua629YhJdg+yQ
6lF5JRvpXUHxQQkeJtWL/8vjliLaUlYODl6z/AGVOhzUcz/fhULFmjG+QYwD1q1BwhRglaEPdSAS
/1AJi5+5qtv60rX9JfWqCQb4u0REa+981XExKhoTbdzWfjQ5LsJ5hwkKHxTqAQtsVwXxXq1YenM+
IwoSgok74EYFWAjVsqE/F4/LKiI27/Ti3/xmmclbqcYB0r55uP3Am4kqc5wECoRSME4WW3Cz4b9g
v2RG52goibL8ATSaBZebla1FdK9TJc/BoH3Wr0cvdUyvM/0wrZNLYZXAJFuEkQM+TWUBgy3UDQ+X
RE7CG2TzDDG+U7OJLPHHeLSNkKyreBl0fVM9yCFQ7iKOE/5AOEVQrV1+yHf4/uckxYrPNxJE30PZ
wCjjrAZzXaPWN5DO8TWPXaq9efJ4fL4s8TM+MCA1emQ31+OKPwso7N9tcEU5kkmevuA+RWa+lkHo
ZGIKWHqnckPOTpRWh6Due7Yqyq6kqHuOhlBnUtL3cxIWrMm2w1EFmoB2xpmKATT5yANlPKQbsjLU
kOLhgs7IExGb4uYXWD193gBRLQKapAdBIjfEy/wjAzMxhvIkONSTlpfqB8yI69gzjv8tbJlgsufp
RrdgmtcyI56mdOY0hfPwEhCpC8vWrvmccDrlc2dabCSUK7tBaMGMhPkAmbS8GRxKwnrEivQDn+kS
Ojd08u0Z6adaruYymQxmEeeQsOw/5qwidvNjHwqJ2I8v+749MRbyLG5o+72w/JPDrsoJvMu+wknV
8hQ3Gn9WD/bfAmkHAeI0J1al2hJ4u8aJ1Ats+4QJgNbf8UcXgKzH7jm++6vKUphe1PchCP1qtfkv
1yzaY91loW9yeg51Zv6OWV1Bo7leXlFNN4L6+6aHAyIhp0u7IIcTnuCNAuGoReEPVv6m6xgsIGXR
wF0Gf91EgRIQLyiUFnIM7CXXjaiNJ30l8+gLGCTuNMnGHHxKB/f3JJX61qIWaxM3Z8Gcwu6oT+0i
N/Rmwt2zqoUfXYtpVmWjCj3SP+wxjRRD8ZIkI3Lr9qHWqou2oFIwM4z6wkZet5kN9lDVecsSOD7T
wLsDIHWvnCiYsBO1KktCF203CiWQZs1uRC/fgLQ5okpDlI6TCD21rp9KSkWULYyALHmSQlAXGZlf
y99UPryuTrtegzkvrAFRypkwsfOIH0+oNcZQnx2lZqGUwbatq0sDhFz93zXKr6/Qa79Z1mGlDFGE
ym1PFv0qAJceriHDzM3iokTHTbwD5zy0YEN+hPfUVIRSzd0mhsvqCSTZ7DBRKFE/Yn6Ewxhr8o4d
wIO6pvCvs4ygJZ2sP6qfTVNGvYrJGr75OCkGA+1EzxsomRP2d8VjAiNE1Bvx06l8ZDeae/bw6jhb
h24l91EZnOtaxOpM8HWHELVH7pVGkhyRb9tGMo26lhPcC+p0vygtbQfUZ/BQmgYRvNGTCuqGFQ/K
y6MglXFpfS+6s1suhh+CoSrROYmhqCeFeo819UwYmovQhhuqlrO19mx6hWgbpYz05gY0cEraZBPR
RlJDRB0/3FRbr7Go6Ww1vUWtZxeGSlJ7WMZms4GLCgzp1aHRrtahT8uEr9OaFGF+ASohx5LRy6YL
fmoH9tNibrdnWtFIxywuur7v6jKrhGEhPdb/kek+pe1WZ2azxVgRBn2JyKgA+WEflpkIAKZfRY0v
o1slsfdJ2mUA8mM7pB4cyO2+fMiH7FNTVFtk8xaINLw+poDpc4SOoZYxowsbvfzFX+7XfDfZNZtc
JV81sOTDjWjszydNP0mT3biqX6GoeV+OAxAVaTeBDR7PP5Ac5S4QiHTPDpsMhMuGfJiUxGdse+jl
ol34u6WqaLo4vSLcDYO3QvUTWnI/FTmS7aIdZ7XelBIqalaoljoLJvk/hMIZqk/ta+zljj7LCYo+
oEe9qLB4VU+UogUSIRKSeJJHtdSzl+o0L55RWkimrBTLSBYdeYyfrxo/N+T5p5nb/Ch431oxpT2o
s+G0HaE4iV7IwP+ir0J5ceOx6gdu6CWPVED90NtYhSwJkaZYEOqOnUosC3NdqeL+2z0y43HscpVn
OUbh4Bt5JG5bK+9hu08fN9NVWrbX+b7kArQI2HsXXCCTtndkCsEOszbWwteT2ul7EMfhs24FHcbX
pn78+TfUygUMjHRqviZwczJB99MUfIStGkgNJVpZOYGh72MVzf75scfBFhYuHBuamw8qFYuo6opn
fbzCzGH69dmLxpc6DONPFy9aitVXUGlWRKPdIqQ9m2U725NsmJPugRtxZAAtKeCwXHL/yKfIY0y+
L90riEZxLxFLXMRKvUCaAB4TRb/6S2ytra+2qZQAgXPMrZbtlNGHrkprj1yfupD0119HdrCjlLo1
NEWpa+aKQXtKu1StvflkaOTc0EzufJXpCtePQZSs13p3cvJs5OH0jefvxFa7zuuSRZg10Tid4yRW
MCyBqZ4xt1+cmzWb4syuaU0byyPDEtQ/ESwZL/ipO1yBvWMBmgjXfqooxft9KcV8nM32crkG4bbM
o9IpBeX2kGSGvhDsE+kVF4JqeymE/q+v+OcNfojhr+UNYiRxsKjhLVH59ii/ROhbhYEdR48OU3gd
AMJ2Jd7PE0a/EeYLt/UbsrCnj/Ojm+KtmCVPpLCAPVCPM5tAn/6Z1Ck3+EXeU3RHAcuQk7B9Byi+
hxCrAENUs5JA47iijAvsZ4j3ikEGG8HI+klTHMhuvaRPodu/LG4PFESNm0CJM0q9hmvDkqbNJt5Y
M8bLLsufD6p5iGClzPc3qsqv2Z7vObuT41foYwMf44FYtSeEbWDEN4vA0bvdZG/+L2CsTVyi5WbJ
P/1Ggk6etkotK54HGWlPnc+fzzPmJTgDCpWetY5RuKxAoIrAbdEWh4XfAgyov83MhmCVnU4+Cj3u
yNBvuMmrdQ287lS4aYOqwn8ru7MkEUIcf9wZNur+ILgBSExK8n0pMwI728KXf9ZyhVnxZ+uZFX5S
rkS457YCNjpLWwoiMYTwI5bhpTPH1M5XVCLvpf0ICPzBMxCvgFaTR0Iazc7sVYtAUFIoEXL+KV8I
sju6Gu0Bdyv/TJAy80mnDslXUH+RbsYR44BGuEmaEdgwzxT9+bX/+tRKaV2o82CRcFf4fmD0JVPK
F2IjbRY+6eUuTnV5d8ftbr3wuqR/LNn/q/zDgIPgxmLR1b1b+uxyOfphGeeKq000crF3hinVy6LE
Bp5nRpnYYDsIdZBUzswhqLoHD2VIRh4npDOXLdWqLMMS8e6BrO8tVc8dnSTBZ9EQ0emKSbNVhwDF
BNrwEqtBscOsnKuwa3zTjhMdnRPthnyfR8W+BVkHbeZBiGDdssFCzNdHXGzVb0KBnP2evoC/ZRNf
o84QoDg/Fk1T9OHitFEdn53V9kzdrShksUcfGnLcD5lVaMCM2aGnppfRTz1rtOqR+4pBf9N+ulZE
jryX+rGL9N59ElrSpBOoeN2hFERuCMuyqNjrMRVTgUPXzNd1JN05XFeEDoTWVSwQCsWR69o0nBoa
r0Z8FMlEuQa2IrJtjcGBRybqO0eOIvJPRdnpm/G09DNAxQ9TOlGbZLoYZJeheE+/hpwEkP/15l1f
boojuPV1AYG2VqgfT8gCC2oYu+o3lF2oYZht2B0C3PwkmuRowHVf7sPppQgnU+je7jjLDOqfETof
Xa99xOFXYg85X2bNhXgiEYC2N1hEkxlzZd3QJ4rEMA86kmVtKMcAiux5s4Dc2F+qaM2mPg14FL9P
JkhsIhpfJqIW05HYUy6duDLEvgHLYaLuSEIi4kiL24GrHcE56vlh06lhW4pALoTDx1TPayvb5DU9
RUIxoQ+JTwPnEBl9HVzUJtvokGcPzMxwF8B/reb32maQMnfGcGPsmqKmEYBnv7E5TfDJx2VKm4BB
j6HGZsJOtDqSJFmSisk4Z39q2n+sWx46azuTk5xvOdt4Wb0CceaC4TndcTHhz9q0zb9Jjy//dWvQ
O231SQidKtSxKM+hpfJ2qjkrhbJpPkpz+nnkysCZBHF0T6zzt7yvOYBztir28ah/xkSUIdxFrKJT
RdqQ8yIOMvpYoaKO+OcAMrTP1hAGa475HeqbP+5hC6V3GRFvbIcjdaGng97hp6mz339pr490g5Z+
7JUvrE6HZ97qKuBP6b+e3o6cYHHw5GRHOgsm7ffdKilKCCNJxiG5lDrNV8DFRMTevFo+rfp0ofVc
GYXExM0vfiLyTVMuQWy7mWlSI46uEV0sO2Vk3GjD6XKuIAmVwq8sm7VhIAo8XKbafeSesvEoRoWV
iPj/Sn+KnACjYfIiGYvJNfY/IWli+IBUBrX2OIb+DPGaDj6GkXryWzf9ODMmvOlukwddQW72bytQ
DskrN/0uLJGPq6M5PvlKH9EXfXiymUqKvKfKl1o/87w1p+7AlpHzEGwZCR/nEAAPNDnOFxIJY9Zf
x8SJSNnWAHOfiLsl9WS7x2hBqmvuvSywo2s/GCxfAuRyNzyIszdWgoPKJ9ip0qrk/voitbVAvD4h
uKyaPuTMe3ABsUb6inbIfj9bw1R8Jl1Bgnj5Q169k3arhf6K4BRlj/9c+CTwpJg3QDyKe5oxGMXi
XagFGUZ0xcVp9MAAxWtdAppkSVA1fMKhfZ8nRf5/baeUeNOaXsgPAto+BnZsYWiWNts3b4SlaAqT
9VD9vBJ/MANH8vQBMWSA8nEDAF5YUO1Y1KvlZR0CdJPRJR2bl/byx1H9b0ZxlFn2FjxkTMaYvj2v
kUkFNZpWkow6kNOJYFq9JnBDCTMNxkd+yIprszcVVBc8/ZsUYKHlUM1zmovMtXOzds/bTFdyOaqS
H9+Yu/yVjXZBzeZzY7z0cZ58N94tj6m2IaovnfEysK8W9Cc9of4CgKAWdhGIZs8zyJZ0yyrt5iyv
V5STQvZJmDVPUnogrhMoBU/3LYbbuNkz2dArRVUY8QuDMjHMa5CTGc5bJBehj0TEQIci5NsWGR1N
km6i5XprxngarTDsy4nm5sp4XmTUJQUyhZ/OqqH+AOUQ4BxhmDthOka7ftGwBH2z9OvAPIxBSPU6
j1rHwQU+YciFyqtzY54lFT017l9lb5qtRafKo8j5UbyDaL4u8y0ik3fcYZdtbBbNbMY9qjWCxfAi
o2QCfxwhPh5rYZkigty0NAXAfje8fQCuVvkmi4nyK8n6Mr8LQicbdnlzIumUhac6jGzM3sBq+gyu
PZYsjHJOgxZS1gpqStJnJx2D4TqOioyQFAJvaw5iQcLQThs0bZaQIejZBDzDQ10jW1iaZv6PW1Le
kbNlGKUV6Cu5Rd9cJG1xwtBpEMHCPshTAtRwtVk4dkYq6qtQ9tVojF+JSIMM+ohMtGcRPCnlKaLi
1GLmTQUoDj6Rn/tmJ0tY8hI1nXPigbMMhuiQxxMK/nVTQN5F5hsPqCZThBgbRo6LyuAbkREWnSgT
3QWmU2O7/6OAKoCqQifpJlpwLV33/AxqUcMGE+1SD/+laPaCMy0m9RDHNEoqptAG4K6DfBubOeTG
B3HSQACT9DL3IRJ0gq2FH2E/HvSWNjkn9sRl/GOr0+xXyd0HVbj0ywDwWvO3QHttOiFj2WRMid5r
aOc4fqenG6XDYBtQpclZs6mC/J7JMHGGA5kBA/Udf4bi1MIpwf10JaqwNSr34JAUeDaiyAo9rPXJ
TERzBvT1m03U5FE+MJ+atDFR/reeliiMxGtfmnHVZQhfgKfBWQjB4ILTcC0rwBKyCBD0/BI+Ge83
pxVIFNZWvbDGVfLZ6vTsm3bJwI+/t9/o2xSHVprx1nPXH2bMtr2YYt+2wSW/j4A1lbzvaoqjGNMy
Z2GlbWXHFhWiJEoxrT4VUZQjCc/Yiq25Fn5RDnE7tjii34rY9XXWhTjxtXaQtqcQz2HZ3BmEeOzS
BtMQsHW7PJgwbLup6gr0H5Q/QW9cUMRTFdL/IRLhaXTnhWUb0889gsTawSndrVfgyWzrjclGobl4
IMF9BFGU5J3r1lgHX0rPqmxmbeUUGihAocNlrhvviMZsPCJDBAK5csXFZBrKBWTdBY8ERrOFiSJ5
bd2pSdBB4iSMWy/ELXFkmfjpow5O14OkYLUbL/eIIokAMhHhucfHM+bQZqNvAj6GWhmv9oqKsCYZ
sG6HgUPcpb5GxjzXZQ0I53H/eKMDX5yKqKs5KCCYatpKEU3c/JOHN0eXMKkIUE5FRUnBsXS95AAc
Cd+HpRzCGayFwvtTC3ZIbKxxi7fDGYAT48Tvru4xiRnYApZ4z1WSlRdEe35GRP9MNcfETBBsu1cn
Bk2wMeyg9TsCt2w0EBI2do+E1tf1WyA/3/Lk4ewaXl2D277r0m4Hn7hOZGr/H+g11qNjPUlK9crc
r5izg9wYtSWuVJ6FkBQiYlXjDAm8zTq5a6/TMo9tYEZ2G2XcY8lT9jq3GqGAR7+G9HUk/8y9OxeB
lzYGnCtmyyojz+w6Heb/dI+yxBkp90I49i8fHcKfVCybn/XB+2zLJbonOQTfw86Ye8V195tjvpkD
1769YBq6NPzmXn2qqVtd9fMZVPsSdd3XHuc9k64EcxjTQFrYWlHibYNVNCdNJ1+SyaqnZ4EZV4bH
6M2o2I7ao17dFETkeViTbV3ARrpUQa3zLj7kjaeDgxYD4fHtHh89+vjQzAOUBS5bm+I9D+c71MU1
yYcDPG4ouXYg1a8Xe7D9If13MHHq6ZcA9FBwzGHnG1K/RYhKgwqv0ecL3auT1lFoKlFNT6Hia5vd
KDDo/W601bJoGdhRH0y3+c0dI7CKPG+XP4LSGxDFOCWAvnt5nzTXnAObcJ8oVOZyoU38fB9Mpk7W
Y+2V1T7Xa2brmx2FdqhCnQUCb6hQRd93e5QjKEnHcgbemZ9jitE/AjMeoOokBNsSII+sVCfEFuG4
L0mwnlZg1eL0y9RAQpEkEfYSiro0rqfhTdG1tRc5RrCi353GvYibVyrIOdElwdiJx3BK6EZ9i0I/
PXQImzB5tgqK48FdPN0SFPW1ABS37NLFhE7VctE7DWUIeyG5Zj5qXTgTvabm5vH7XLSEki/Ao/+4
weJmowgTEiCmR4s6DQM8UwcqkRgKIgwcc3Dd4sbAdmu6HNQ+Q4cPBYX1Z4ao0dc0XRpPzJslsblh
JBZn782fXEApXWCiZEXxyy9edtDLOCwLyfW8E8437KLqthWStYiH9MdWbBDtq3B7sLChJO7fQseK
cFSQYX/BrdQ/7sDZTZuFSXieFcTn9HC0KFTaOWSoj6XJAO2z852XPHYh7SX+zGwWBD52HAXhCbie
hWPeYl8zD0sOro4yNc60EZ/neGEoUVmrXsnbjG1HW0Iux23S9CygvtKQ/ydL5UmORMy1wOXNFle8
zfB4eUtKRfs9UJH1FK6iG5XGvR5+k2k/gALefZUCFZV1TnIdldvuxxXUS2gpW2O1yPpPM3jBFpxe
+aqNiFIBEtWPvMn/dv+rdpIZZz6J6bHFkPJwPLhs2/Jau4hWVWDU0oNg/68gvWmsxT8NUS6PBmPl
MMLGFV81gT3WcX1ZhjKy5ujMXQRiRreWryopnO95LPETPS6pCUfnLuvdrPY1DlV0J7j8/TjVRLaH
r8zi1DasJLf1aM7NA8NTKxz3SjMCOiZMNV68B1VbT9o7SrIooXihJU0CFNXW77twOvEPHVeCYe91
J4jkL6m17sdsqzfEcPJAukBtv9Os5PIzoNLZogGFvNMfAx3YFxToWmPhWUrR3PwKOMT2fgJkjgYR
zr+jssQNUfNps3Tm8I00J9/eYmxHne07rmF9FjwfJjuT7nbVV13DMONvAEV67bFED4hT/ZDOt/tw
oQvDOrWrk9giv4lOLUhUZVU6v7FBPf+LQCsH4l8JNuUNomth6AlA4U28WuW+02JsB4JUKyiCo0mG
zOunIQZYaRl/DCPKbfbkZxCjJx6StPUDoKblZqqyM0jQ4BAsABpwb7YodOtk57MqDAC2zqM0BIDh
c6MqM/cn9OGnQPQNzATlisLwP8y32oTociOzmSksTwUfDq+Q2JSifCQ1oTZIW21Xvl6Srg9xo+Aj
r08hEqjudQzW2Mpe6RSbXdsaYhr7usZzW4rqC6N2uyGOiCDEAYYTjcS2mPbh4EfG5lm4wO0RlsjJ
WCrVB6CXHIur1Idg6PAGfSU649mH/Fk5LM3tg87++BpJ6mtwvVtStvbDeVBhzsWiQNZOFGATVUh4
xpb0imA6pTWmos437FELsB2moOkKGQC9wZZKsOHhBLuSrOvSTwswyA9lPf7JfILD0KqEK0rILwqQ
6WaVz7nCInFyoXaH9Vz1KF161R+zKxK7ID9QnUsAtedUh/zviiR0CCTFHtFAS+lxA61ll33BwC9+
wvbydvpsKP1R2ahx1UiG28OdDKErtzbxOcTyBmncOFcgPmmbUdP5vYwoS5ehktW024M6p8KNFjbV
Df6oGJVKPXJ9YIajCTiiMqOjDDwXpTbPsh2vO0qlN1qPt5USPfG9UWLjWVGEO7FyvHLmdfok6tTv
cp0zGBK6EdVZoxoYPHCppneas9iu9Ssuk9uSAMosvaBsJyVOnJVMlKeXyfjJecqWCSnyA8YDW8xQ
aylzK4oWswNo4K41AHn/BpdZVmzSNQgchy81BYaQ68YE2VmclHzhROx51+2W2QlLTWdJuTq00cUC
t3TrlObNj4id8rb0OY0BZ974KhnnVXCcAdOr6+LetgRQbOHVJOkSwcGkRzf/HKViV96+EP20Ez23
3NcFFGmdoo2e86GCCBf3rtBZlyqbHDvLVII/4Eph1aWQRBzT6cvVYjf0Fx7S4yL74p8dBH9X2b4d
yaJQPN3yhAfDJCpMyZc8UcXFfw5KtWACfU16UN/OyKuzce8m96/kYuNA9z0MXDqHC6zEDzkhLyTP
VATSbEdTWFWXmmUq7XPMSDT3jowg3MzukeMwEeTJXJWhcQ108UMYKfsJ3fxnlf/jfZW8yKYJaKww
9nc8bZ/Q4fXFGS2Vx14psLyytCPQGGyaOoV9WUHtF4mAt9BNXAshofsuBZ2dLOeyn/mnTjcddNsQ
GZkPDO9quGNXNPViY02DQl9/3EGXkkxwm2Lr49gzDSbHDq/J8dV334WoLLEjDa8crxzTrYkLBVWY
bNm7uAwAoEVP957yq5VcS1iVNmRZ5jaF5CbHGsFe8VsllRSzLr6/ySlm7OvXIbG2/q8wI5BYBRDg
Ag79CK7/g5aVvQub0Pcc7GU7hY4PB2bIj06qXcoYRR10wf43bNrksHGqacfGuDHmnnQwF7veR1+V
DHzmkuMFEsB0V+ZUnVU96t6hSHjZR2TI5Y6pD3aQHUBuzCiulNxz4i2yBifGPzrb0oJRnxbTCmmJ
yNgtEOciiFlZISck7AcO0omF8gh5GLon1OYHBtpFKfpTckN14bHZrvgGqlUef935y8WCXibmQ8OM
u5jJUnpC5GWhWQSNdsOJ6NP43rI4paodw0BsBCp/1hS8ISpCWIJppR3TaxYtNFa9UQg+D81I9Bgw
wo6sueiKQ/zAc5QC8bnhtzVHNBAwq2axJX352AYmVfNPCzZdmnQ43avwPFWutSlG5mioiCKBZeNy
IKQ4wPsR0dhWagrj1Qd4K+QK2j5dXz6sGwRNWKtqXpf6e1Sk5Iakn3iW5uNW+SfvYGCitQy+9Jnk
yaYLvswiRm8qtVLMY3kUuFrlBMIa/tY7uGlHCZbmQP/S2U6eRj3VRbHkaZNQu6hMIZgwbTt+SjiQ
nmPoex1CeV32ONZuuEQDcatTRyqysoGJqGtmC/r2a3XhT1S2ufu8zNzBmfH0rK8X1DCKviuk7Uqn
YRisEb1FSj9MpXY33bQn965kNeYcYoSV71UKi0xIdv6VuZJ6lm+arkKe38hYasic42Y7OJe6LVJa
nxu3z75OwU0ND7jOdGWfs9ewSAst4k77FTJXTiPzXTGfHxA/VUL3+7T8lYY9TMKCIIxrJ3cLHYkP
5WW1qcov1/cN9t22FM9pkV0GqcNk18UIiM+v3lfr2k1ld49LLMZLfZZF/I4b4Revl6c4LhetJyjk
U4IO225Ch69OZyFRihqRjhj0sfzeV4v0Ik5NPTEaQcdyE1L7umAZY3TJ2LP8ytxULntvbt7btbtv
IQr3FMcOR9Sj5GZbX8PXbWAHTuEoN+E6idxoMu9J18Mz11RljmNvMm5BwnKzeKjStknGE1DPU2qP
QneSkNn8kTqT8Ra9fSoyeWqXzne97dNxX26SJE5vDR78DJDvhYaqBWgsitXL6wYSLKG5U2pTrQ1O
ZV7loPpkf9ZKaLg3yh8npQcpnC6iPoq7LC4W19Qy3qpnwRCtGN2EtHXJA7TFBleo3jeVSwU4o34+
/Wah/v4YCzQ5hcA3LNwcm6BJ7h+SGCwa/TXP4onghOIxucnaPN5G3fxlP/6ArMoQSzDUsXV1D8yK
8VS31h9rSEWUfAiznNFBJ4apvfBKST4YH3vUhXS1um/ErY2+4T/qxq42Mma+OcplByi9VlbZhl+Q
w0DdVSVYGfLDx2DiFfmkBLsIdIikzeOd+2ae2+WrYu+gykCmethAfkyzjWY+lZaWLhmXf0J3LstM
XNcf9jzBZCEI6CSpbURuqeazuQ6tz/5mwCkZnTOHFPws+ZTAwBaRmdvNgIPo4ZuA0PHwyT1LKX+X
YhVZ9QQl6uK6oFKFGmmc7f+v0MfuwkhEmZsHj3IgAzFrYcRfiPuGkHBicegovSNWSvyYBiCQ2iZE
gK1Nh/8Nu3HOEqutGyRQKaMI0M9J9eQ1Yu9GKhnN3Fg/VvItRG2MyyyPJV1qtPF9pKZEPpV/DRzT
4v93UOgwyy41ox69rNyKqhx+bYo2Hw1pehhpHBQKhlmFvNPRak3PtkgHP/a8+7OQOI2aGdaLGlsp
Yalo4yOryWDYSDYBl+SzOCypbMi98LXsIRRhX0PItZrrV7uFrqAVmlBoCPW1ESWGanwkA+56MO2J
hOP/pkCPH+1euVzcP2Potg4JNuAY1Cx+wVBK7TLlbtV9lXh8WhwIOgah41e8IcIBq7MnAeBDXiAZ
lGvbXtedII9O3YCx07UKix5h1dpUXoI6bjOd6usOAMgluOM9yxPgxIdOhY53r2onNLJVUkxgQ360
7IX2dgYnq3t7Z/RC1hgzox4h7N81+6DWO6z2w9NBkEkUL+uovRH8ux1oAFafuoZzUXzNnHOe0Klf
Mq+Mp53S9JmpEgtPGXeNy0vGSRw4vMMIfT3mkhLGC3gYysYT9UxNklZwqYlJL3vycYWzJthEWIgf
/mgdZaUnfJ8ySU9oz8kiFMwi8RB2rI1GTuItVo4O0Sn2YgmRUFjfTyHl9PvD3nELD33kTS4YunNk
DM9Fln+1DvGT9DIHoi37wy9+kJQcPUKOBf3uvb3RCMwR9mY9xarImenjev3louuxwPRoMFTxBGk+
sXh2cBKRnuh7ZDp9lHdfUM7BB6idJybUpWQo2V5Q+l1XL8sYoj0GWSD2gST+K5EJWPWPWVv/6THY
5YlLTN0DpC63UqNPo1uHHRlL1H8eanMTjdJwAbqmwzeDhnP9eu+azbEYRMcp/pS8R/IfczdjKcMB
oXnnmuhvp9btCzgAJvh9e7R/5LneaaFILbSmXt5skNETNu8DbX4O8OxHlxPltKSjFyBPNL501Yph
OAncxujZsux1QiMz3+I7KILXhFxrnBTyi4k56VIr5KpcaRcJTF8l6Q7Jp3NRIWEEWzSLXHfeKvzE
sx0DTFic+oxNLtbihy7MuAtJV0HK0TQrubxZWraZMd844/7Lhc2FJI7o14qmw7krmOZJLz5g+F7H
H0RdbGNJlh5meh8liLGcVd0g3OCI+ZAQ6TUX/Eu8dex3LhbxLCt1+ojJ6WdWLV0KJd/P7+0GK447
eeu/uKqJFbNcZAzltpZS4e/SiTVdi4tb5nSz02G/IhYtt7OoC4OMSGvcjfTY1t18sK6kLUYNGzYC
N6IVVrQtrpBioLclHvFTOiyctmN6tucPR6azdD3YuPbwVwtmis0Jd5Pu4nRKuR3M63mgf6wrOiub
AJyKTeFJXnDHSWrLlTB0OJMoTRC/QYrW3/JmgWqNxf8fwGnWN+Gamm5N0luuITKHv9ZFvGsHOd1k
50IRLf4HiHV221pq+6SaIjvGUA0cWUv0Ep07M/f7Qy/mLiTV3Fr3yTVfj3aFWVlD3whZQTmowmti
8DtNyUl31bowfNshFptFuF0GB5K9SkRbl2HFDG+lPZuTI79/x75+qySX7mLi31wCipU3go8zfykF
7jQDJOh+LlYXjGRGlFG9vrHDOAsHoZv+vPqavZtwo+rhQlxucpvqE/2AhBbbrJkpKCHX2TTwbQ8x
p8Pqso4y4C/7vJvzj1c5gGWe5dEJGTVUBz3AXo8HAXXKo8lylhB8aHeob/D2eqrSBlww8lnW9MeZ
WQPJq8qstOuDBlBC/jqrVTKuuxH1wVm9QMYMqM7QZovNG4iXUOqPOXFL+nvTUDi19IDq6DRIYAk7
CqNRL2pFJYoxagP8UEAc+6sdtHeolg7JBiR9aN34Mvo+PkGIBBZM9uFLgN0EXdHzCnqaNV53Yp0l
HL8Px3Wd1VzepnnnSC1wNRG8Mwv4v/cpbGBcHJnhQc+rXrkC8HT4ILyntzMCCCc2qD+EBK8Iwynv
P9jgAA8k79hnheLRFYKAq2kHjMvj9kR5FE2abIOwAFLzxiVk+HN8L05sKigRxHjV8KmHAZARtqM7
ejw7w4TI33ILUwR0rvdQqHT8RN931Zt2fuRdC11eVF+JVoQx4NyEPi335SxKdctHLPYMcFZ3RNb6
cY8+k+Pf0GUWRCjR+q/jqd/GFBgkxVNS4nepfwiYt90rR5rgDnxlWbQN/zg1/ff2yOPB6TFl9A3R
tBLB75AO6WA42gawH8URxGqYe56XI6sHM93dUelpCINOuLfgtoH7dB28P27IkVQJsexpW0GL1Maz
enDzGp+LfKBLSCU9MTgGJKql4WsS6VZfpw6cowQCZ82EQvMUeR97r9NrGhvvMpkvpUej4vzUqhhq
fSnINkmh1v7+VIwXSkZZ2rulTURNT/QLfogLj/ng0pKeoiJ0/MEfcM4aPaipTswxzwWMqB5jmsMN
XQ7/iJrLegld8s8BUWBUoXJ35bRFI71V51crm87UKQNVgA5l4/PXiKQAXvzp9QXtjyD3VvsWWbjV
GEe/hvo/FmFs/6w8uBb4avxM2Vqlayo3+fHHObR90ABBa5e/lK025hVORKoUxzcAM71jVJHdhLpA
vVWLRG7rsDNFLcvRpYp8hzHtD5HNuVd7BS/Vh/UnLjj3blqjgaXOYh6zR3/JkhbA/G0d37YLbVfc
dWYKEC+x+nshm7ZtbKvVXu6uX5xL4C02BwZoGgphYmS4J2kbMZuf91ERNxfsXQN1AM9ozZa420ty
iqfwbuGGmAhdqWtAMDxg1UHffv65wiNgh3oLFCEfOfYo7eDc1faDpa9HTutq/wvztLIXj7azbq67
Ch9xU8mvXPZ0gzUpCJ8XjmuL1HrrO29brxaYZ5/A2zM6subb84zvKpZOnAYpXmWjxIjGMZyV0ub/
50UD38vZFU+ddZ35S61g0a+hFSOQI8SA+vWpkYXaDpt29w8B9lKiUYFz6p73HWEegVZg8gXHqcRr
qtVIV8EUbisn3wYQhN43dbVjMUkaNXG7IIxkqfDKNHaKQdgFHVnmKMy5kXtlvXINUlxzYzFrebVE
YLX0apYJl7ab954OiS1w6gC1T3pKrzY96to1EtO/aq9JVH1vr66dqG3Xd3x8eGbN9M6NpM5EM1HY
9mijx2RSIWBjZtihsgiWj/LGV40azUwmT21BM/zZ14QUha3HujOHuXnOcnjrbUCnLyGbcmJQSyPj
n+vOUt/f/rYQKjgS6g6rpg509UZosCQFJ+bzrUDeTc74i03/FUSly/UTpZyjYd63npLIqcsNB3FT
YuYd+XnG+ZzhKlRvctGCnpa/YqStNGEha9N4MU3a9KZUvKAh1D18OirsjqSmFG39j7aSQIasj53P
I583M4+q1YBmrSXuDYvXo8nxQttEs7csJF+8eiWis/pxAIdam7mW/finvS6ZPzT7m3+kGpAivXef
5gsjenkCfNDDBVAz+o8/yxxXw2Ib0jaP8c9LEGLDnWnj1fTdEgm5sQKwI1kZ8Z6yOTrGm+PZmX6G
cEf9RiO/H0XOwMdRyy2OdE170WMtWVJeRze3cUJyTeRENsYAvbLSZ254f9XJcQ5pBORB+HYNRMZF
WO2KcP5PIWdxCd6KhtIX+DBx+iVcwVcTfXzyZx6PJKGB5GQQY4nmJvpGc+92ZL6gQikeRoXn29lv
y2WZMHI1bWcLVoj2BD4QOAQ2gtnZAilbJtLZqdY9GrMGI7xFvAKFeoq2uVBsGYTOC4jL2hyYaCOP
H9Jhh8BbRsGwLscDiorlG9Te/2/UGlppnsan9XbcqYL70OwOpdT3P0u4e1Jn8g2mJxA6OtvfkNEA
GkCD9sDtkOOgg9iXkrgX4Pi32ycPTtniFNt84pW+iVUbJ51vIvZBhO2vS98VJMF6bwZfnVoy/ZdS
fUsH/sHLkXb/QGfIxpkMaHoSHleUwv9Mrx5TJf6TmcLT5Rhk+kWS/Dxp9QzKhfDbTi8Kz2b5z88k
tTIk0gXrpLP24KYocSVhqGuu37/KgA7D8xilTk2ROoCG9yWjYRXj3g0rRE7B8NgoaRW/aHQYH0X5
lxKSbVbBVv68uZWqu6StRkw9bD3poTnT0EwegZeFpTQegJZIx+zhSe/tPBQ8QMy2dqChrTlekWcZ
WgoffOu+atqWLzUWzOWzLk1M2FSslCHbYIlzi1sNKXwDYWyu+xI4xlISs6aG4ifRxD3HQamH+ocB
8s7JbhQhslrsBrpFg+36TExeMJg0/TWu3hpDSkLc2C6SWZIotQpf5vY79iRhrf+y98u15XMYzlG1
U/COkwRiMQjmAhIcDPEktrGviu1pa1cwdx68hvlwMEqxjSkyhl6WgTuJq2nvEJHPMcHCfH0lyBMe
t+SRNoV/PspeN1cjVE+tIP8tO2NNxPiYJebxQ0kvq6urkXgTPCKq8LEEbXbLzk5vNAdMUGbrkbXy
V1pmgd6AbV3hdaH+63EsfQXGZ0T/WSBVcJaSa3D44aCANh5wvaD/hBRt7kWVBKpqS6sFuaTLFnpE
LsbNViBRB1cfDMkjau3jbQxlSozVzS8pArxTroQGItK7Fb/WRkYC5+6EgkMuhiJSsXhyAb+OqX7n
GMFAf4WzMS6gMbmW0RNvMDmmQ1Zw+ktKC42xBK9wIxT62tRpBsY2jTtWP7mePOAprLNdgeUhy5CP
0c617byG+tkW6dTRUR3mHVJYFZScpT27oofec6aSGgVriotw37PJbP1KwvNFeDJSw+VC+gN0ghdM
tQ2vCdVvvACXGRp/GQppS4N0++qVOMCSZ7WIG8g4nzGrlt6uN/zrYcyB9mUK0MS2l0Ayv1Aicjah
wt7qqyPJ6QQBiRWUYCuCIobiEZeUvLIvy3Xoz10XopPGx3vw85kkktJCYuLD0iwC9TMuvaIjy3Nd
GFJnoGq6R5JwvJfHfyQ946q8m9jmwOKW0A6SywL9kTPUViNLpNqfXOwtAelk9r3tbllkUAldqON+
d84PZyTaFIQho20Xyn+p/YMDNteDmDSGWSYxWWsxMcdV1T25xog1Nmx6qpLdeUGg8VG6Leg5bROw
Sjg2cJkfrGDuTTiAUkON2NBDevkXGz9CDNX/HelSZnnRtpUG3yRdKQVwLRRUvQ7tjym+NODt/xoi
Z5hf7+5CbDarLa/+78cBKDjEOutu61dzqus2/GZP+tO4s4c8q4AuOxer7r/LNWKw4TybMljkZD78
LNLeAAq1iNtDjt1+lOABB59A59VH78PIQx009H39uYcx7HHGKA4PyZV4ueuSp5rhZCyKlxzZ+3po
xDd5VCtkaN/7U4oxEP/Lf5GLbfxUbO7yebAZo5Oef+1vNHw+NoecxJAN6BwyQhXkjoJJ/G0QJvgS
82jxU6YpGle9TX1XaIYEmiIjR7PNnWMPfeoyq9F5+4KrURnFWh7JYykJffiSTFRa11+Q6c+H4c03
0qZQzeSfCNn8OI0RcEdZPcEFr4mxWxvxK/97UrPvSnTyC2QkRmNj5lVS5AphK0uSrnwY18bPTBif
CUTvDOWwy23pETr55EDA4JFhidwIgc/uccQiPG9vCwcHWf0swiM9up1Gv67dfI3BQSkJalf0jbog
P3186x5BoY23M2MOwyvrEyECw5elFilIkPPr97fQbXiMCRfR0ZEmV3xAVt8ep1w9uYTRQMPMaS1F
spORT3MT91z9HFhOb2l1LnGkfgVnp1mmkMWuCd7vMDxNuAMR4YPaNc0w75O/10Z5Ey93WAffHJqK
SE560jMPErDMj+MAzgLt/j313XVZQAzTCG1cdeewBu8YzxHyvUUfXap4Tujo4oUAlmCgYYBOQGyB
DIM+IzHUEWCBdpZe64S7TBQNmOkiDTSbPsPnc+pg1BCWXKtEjlRdv2i68Mxre8xb/vwLGJ5vrQoY
f4g3qZ5I92KnMcYBxmMWG0OrmTIf+r32AiW9OzzD7BtZX6ZseR2205VT2Jq/pTTSOeB6m0X1DJHU
DhSa3K+ZFtDOKZzQaacrMDQ23HuWl/Ad12MQMh+Dt4JSmc6uUo8Jsh/P7ujAyf82UCu/i7waCBN+
FXZDVBL/q7djWwSZO2TDab1M97UcL77wi4gHQPFJY5X4kRT9zCesh/v4/rpTHwUsNNV1lZAHz92K
OTVmsxlSNox8ckizQf8w2QRLi7R88f+t/xAAi6XbJYlmU5bCW1fkXgauBhQDOAp+BPWzYi4w9C48
cRGc3RsA4GcdcVNHZazfWQ0bAR1z3mjJWj1mbt8X73o7scQ/6NsgLErXw8sn/MiAFPDExy95FAVu
nnqbqmv/4nXAAHxWCYWrMI14gfRoKhEnuB02BPIDqK3nCsLfPCb83GAgBUuORhwLyf9Vz2sSX98L
6uqo7Hq7pnLepbyl5FmQ2BDhSFWSLsYPx6Y0XRU4lbK5FIqkwu1qnyCpAxP2oh9uaqGQGvSv1ntS
0ssVt25bbiau55Bp8bTOU3rDjNmfWpeNNZFw+6iYK6uanyZ3xbYBMQ5wTsfE5Fy3UpiZyPZSwEkX
tFBKRmDvxoNm886BDMOizdUFinPTYtB1oF/4zvT21ayNpx0wR488AUuMSSxvgi/z9KadP2EPsFnX
DONQNS33H0rdg0nHL8bSoOZR3V7joBTa728h4yxajM8UR1KZ8qte6jbr2C2ZHPHxh0MjfN4Qajgu
xIkVXIs8HAdVS1gYxmu3d3j9d2/ndoYwicdNSG59faerJ++lXhXn8OyI7mBL+83FKqYwvV5z8pRH
IzYQvEhjtIHqcAOD+7S/xe6TjeDxi5krb4bpzJHApB5d69jR8cRNM2mR+/vV8YKYr6IpPlP1/EpO
Lz/Wg57no/1IkwdirjAzXYUTqUSnvqkmEt7fHuEk0OKEy7VHhWgTGpfIsoPtdK900Wzaj44WL/Dx
cynCiZU3RIdZv9My0sMVYp/pHhx9ihHRu15K1qOMxSYvluzMjZi+jqKic6++Jvw+a8UC2S5HZohN
/tf/UNoVRjnF3yJr1qjSiTYkFIYJXiwOh/8x4pALLW3Aya+tcXR1xXkla3xCQ3CJbihtF1WRxn6R
oofv9EAPWcKlUyiAo7AQi+M5k9MGHDTyTZsgo4hjw65gG2czgr3tb5NuMBuizWc9CR0LtHPo7JOv
JyFHroKeH5fmTunPxrY8PwXUOqndZk7Ng0sdDg9eBDrhCswLZAlrHHxbhAgawsUYtkf8IEEXUpqo
hOjf5zWSaLZHMtzewIK3CgTOf8VPzXfGvoITlyJPt5VpIAn5NngUmpcZmQEm8qKD62d/pj8nF8y4
rxnfHAFZygGqbfiUWZwfp63uyfgMtSjXK4ATt1G8CNKTXxd9zeT0b8ffTRo4cf8ONT3hRSzrplN2
wpeSOavsAdfe95usoaOQihOnRiDD96KRPACjptvqSGOhIf4gz55I7skzxppX+ZS+rfob860085fr
61MQa5+03N1gU6QjkYA+wPgRgc6Bfg1GKuqzv/h6ILZpCbnQP6l2cn2tk99S+v/eket4T0+sLTbG
h1+tj63aDSL1or8bBCnuljzAWhMIIc8YadU5J9bIXGmLwuvi1DFIyf2jFauoK+pqQrw/M4WkJ8tW
0F4G2A2vZwG/unPiJdmlO23D/SvnsGvRbPWhTtz6d7j2BoV0hZzCKHGygvuXlc03CIxi1FbzTuym
DFfO1YV8Cr5HQVNUrE/ku3ezUa6OwclRsdoHSGeYJXZdQ/qTjwxOB+gGXqZX3M0qf68hszHcYAPO
2gpLbr3WD2iUjvFu3+0Nn97lxNSeQKD8vq0oh1w5TNuJdgIh5v8allq7QQO4vNUOP8vfV4cS1fHw
OXD4rE3s1UZStjAr6B9qGxdWnsuLIoi9gfp6niwk/j3jfnAUwuOJ/V6DjlXKGr9894uZPBHmjRzm
qRBHJswvZs1yykYhVTnkgE/l6VCvmRPqeBcLYHS5cWr0M00d7hzrKCT9FkwakEhhXgusMPK44B+u
NBDQQDhzc+rLNVUKeXKCK536DDQa2yJwu6LJBqf1YeTQ4cNTqOqUUXGo5J1C5Xvdc8PwUlLASEvM
k4BuqLYZvNGa/WIN4vE5WE8sgXPYhTH6gbjLaw0wVNyY/BZ1ZS96snjN4HXuvRVsW4oUoXVt/OEl
1erXlOj5nOdFehSTL61fPqxrJ3l/eEWhTicaTD672MHDyadqCpSkg9qsU59bdxqjljSHEDgyCGTm
h0wPdWEIzouq/Buq/ILrxI/p6rsCg+6z+kFjW64EMLLrpK8wWBKOfUGxUowJlJvTVJDZnpYndbEB
E31Yat5Xrci7FXpfmPoloLCK6CIpyhkXT3OFCMdvENrp8IDRhnOdcWr8PBi/E5IcbujZUiyvFKm1
3SuMZsPHKk9BP5fg3nXiQE3AlaqARjnuJt2F1WYZOti2yPerRpf5enOUtGfRwTmt1em26JZtah0n
HzaJzJAXLjxTK/nxJ1j6OmPOnBwaSOdPUzpM/YXyAwpEhgjFM3O12YZPxAP0cFvuFj6cTFL12r7d
ffv4E5h8VjcVFKUbLudwxiwmxX19VJdNEQtChouJU4CYuR3Z+HJK6RDefOkAdgZrt57sLFauxvNE
0MAlA00sk0GLJNBEZZP3QYjGo/ZqrjutgUVYmpOQt71QzLoOBT/nihUagR0jn054tjOxh6/ekUg0
+jgs7zrkAAMDn89UknIdgKNO6lCgJr73aFJqBpyxHtKDgZ3yYnW15RdG5mYh3CEyPC/K08l2B3zk
kZFygtKXJ6zcRvr9wul7LyJVb+gIhZVz3Uv3Ld5r8533FporjBRlX62cDK3/l0VngvMSIXoqSEMO
NGZDhC3wBhGRDmiw3n4vH0PpZ31QYCeC66Y2JhtmnTeMxnDbErwbc4lu0BbVyx/0z6/jRIswt5eD
OcAW8qDLQ3Np+qdhepRWjxGfVyQIfHvhG69OaLE4BPlOr7V67ENvqKqIE4+JEtyvMV4VhIobYDxf
eHkqQHveG/oetHeUmgFeUvGI6DBCp2NJMW+sEOso2Rb8t1EmgFhB/5e9qEUrJYPSQ7m7fUlCdx7o
QXdbc+Rc60j636xlGm6DqlhT+B6oIRSe73DVFWLQ2W1pEFd7zfYOUAIzNx3c3O5Nmw4ejnLMpB9W
m88eFssCfydZsLJ8lFbfRwU4kEC4HMbvU+zFAsdQBfrvDsG64vtu++ueWV/z+S3zvMPs8Ov+M121
gja1saQAvbl05DeJN2sdSWXxDkbZgYZaRHgqR+4gVR2JJXU+qcJ/9VsK9400hUMulQrhUKsax5JL
FC4mLha9eGlzsnqN/2IIcTaCpg0Lu4AE40eVdyVcR5yCHQMh0ixT+cot5vjfaarzQ9uBmA4snvdj
/PrWDdaYZ25S46lupvoQmcZsE+2NCKR3IDsU1RQwPNGFZIejzrdD34Z0HGLY+9+iwJffIg1WLung
0LtGotSES+fAVHTLyG9EnIe5ZmbUoTpYCBply6C7XY+xRa5F+D793pxR7ICA+CTZpBpwfUTllOD4
i2bJhNO3FaQhNgrvQXqbIfSb29NP5aZBBB/jz9YhNVxwOmW+oEGnde+td5uFoy7Ik5aJnfzA4Pq6
fcHDL9Xn01HKoICzYnvu0wWHcfTQUdo/RSz0KZZb7BGhzrDKAkuWrzSi6L2Nq78lzo0UwXJBaeSV
4XedTrvkypHep0USYSXSTVegA1LTFlwR3LFf4OzCZALAunYVfoVArFf298wQKJtZlt7rtixS7FqL
0G4OpGfqS4FUcIVPk7NM5d4KTSEje5w3vdKPoRCexEEcxK/gMVTR90+12OztfhQJnCpuq1N/FBda
n1GbFqHhHZ75Z6hFPr6hqGRdiMxe9LoOjbbuwvqeQfHL+dRjL5mb7dME3B6x2kh22u064WlJI6FV
a80uSrSxlp0KcNCwI/gcI6Kf4fMkAHdDXJ6GTBbdtswsN+qrg3zoje769HEq452VESSBfdqvvSHB
aIL138y7DRFtzFqS4taCkOUtz+S3lXzaW2HEh2D+uyEjafOdERhhECSKG/gn3z6bRrF7L/BdaNMY
G6BrR9/uIYQHsSXN7h0TiRT8HCFkW8cppDzEp+KjKXDn048hZT0/oIBOJOPEw29gNCI0w7e1DqwA
ess8yGMmJ/gpAAPYj2h2woe16KCPAqIjvxWJ+hV05W1MhbmbnvO+54Jwm8LLuRmsf7K71EAnc6U8
vkeNvCGgsLi1R68eY25FMglm7d3tJ4dOo4DYRJMxdMd3Q2FIZdsTvNOrAVPEFI5sQfisGyEX/wTg
Ml2F85sFazGxgCEyC85+n5GToyIWq1d4i3scE+IYgL9ADtB+mp7xIzSst2SClmwPS+sZqi3UX+3v
e3kFG/9Qg39Dbhgh3N14VVaEWTnq2IGuT195ryovWiR7ZNhwEP+S/ADBufbUCt8XrRz02TEWfkY/
pwin4aAr/gVW0yRP/62eqtItfbKmMMatGmKMsrBNEhlM98LvJ9PMddadT+J/MUn1b7ld1h7Gqv9B
Cfvg/AyCQ+eqT+VLtPxpubp/6R5Dl/DDj/t5i+r49W4NWUhXHiSWZPO4PTxEMGd7NHfk7slTkaZQ
1CP4Eq4YubzcQ0ojCf4bFhp2CJIvz8ZCl9AdPHWRa+ovmOlrdOSNdsl/iDoke1I9ymIfAWl6yPbI
07omubZvORFTOFSW0Z2MPyIPufWXvMS6WXrnUTGGVRTMTBq2HXopm0SGK/c+rVdppg4cM1ukvzfm
EP1bl1RWePOG5V4Lzv0PQXmohH5D0hml51+2uiwVUFtklKgqAz3SO8i87IFeQ9ofaW0lqszEa/4V
iAAoYZ5j+OLg9wqVo6JHP0Bycc+Sl8WosAXZfJ623dShu1VR7cwh9+NLVW4vQmPGkADBkORP8fUA
BwuXCWP9u8+epEyNGsB9IMF+vLaka1XLoJRcnuK3CA8Xa0K4NCQajzE7yTPqkJW5SWM5+mAGNSW/
JyiZTdkvDCL2ANT+t99qxTXf1EiYMPgQz4hzrGe7KxdCJfxcQOLd36xDMPkzSKzTzlua0FqB++Lb
WrIDTWFpVqiJaUNhVhIim0d3UaSC6DWALQfRjATQ0axLsAvYaPn11AEyXtxAEkKv+nvmd2+4BIti
KQmfQAMpem42UR5+eLCQVTMtuWtXAaHaTrYFgUPJvtF/V48eoWmRfhzBKGZwMIFpSL0xvmw0iurE
OA+fjb746AhjbCOoSt3gdfsmhOfVc20Ev6Zthq+sUQgN8UikRG6auJuvqiimDsv1K/NPNx7quIbB
7znlp42gGM/JuxlI+C5MOgn5wy7wYYRS568a+/aJlHZ7MvvfnPTNLMeVhSuy1nv4QU+0poOtsNiP
dShRQbFiNkIIm4ICwifOFR0JY2B8sTLgaqZDj5uPYTAXieEDvuueb5z6cZ4ZyKrmBM9gJggbFmFF
8df/NPDCF3qjeQ+ZGz79+/7lDLuOcCzX9eW20ZP7PklBUppPv1aHDy7UrjPR45LN42BPe12ZmQsT
A3GDiauCm+8/6zeSA18VUCNFit+epoTLHIu3JipyalBfsNlltuKkUVNOy4Jj00AGGSmfLRArMwWD
hZWEp6jNCqcf4tE9fNTpTUIxuKWpCDtKxyqMhxRDQ5cNd3yJ83/pHP/r81RnjWqYeHjO6K9QxVi9
wIRU+Xcum0UNFvBj0bUUUBNO0IgFX+qIWEoBpGX+K2feo/IRMzXfJqQD8MPsHA9v4OAjqAgZ0K2G
fP3eK4x/y3JzpapIu1Ei+Vbbrmox2w4Lao2n3+YjIdM8C8IGDbbd822ngSTWlEZed44MaZO0nfU+
WUnAvnjyfj0QD7z7Jeb//aYWB6ADnl7ofkLzwqso4j/w6BaOAgN3KkNct2tSY/FclGVgnT8H2Uv1
XHl0pI8MiBLzF3GZCtCR3OmyO4n0iwS6epb6tkmEyCcQ7YI1C+8HzfwdlN6G+N9LGdtlVmhiBjqE
dqxsFnNBQqUG9Tj8ekJFIJItL1Kc3seVTGHIwWrNEzArwNy4mjYlycRewxWrTqY2owHHUBhQE7cg
AF72006fiL+XacFvjzvi66vMsTdUNjOatnylbtzXnHEaIhWKJ8KeSkyWUJ631rdzgWI4Dxd5XeYs
cTZAGObQ5pd+S0+WuuqF/t9TBHEGDn+42mJrPtZIilmMaMgLJHz2f8hG6nrVaYgZwxYwGxcii6QY
hqcDecbgfg2JraGb04B9WJGnz7Gx7c9Vy3IHSbpU2kLHojhe4ICIUPYdjv5INrg3UVpFsDPfWuvD
8QJje7myzNk6LI9IdIkcqurxNE1svGzayp7eAWbJcOV1q/jL2LamJ3Vocfk+YrWidPgbyrb+Eaxr
qg3Q12/OQ5UaI0Kw1qJxRxb2IuxmxwHCBh1Sz4naNmSgBqGdC87V9J63L26yjb/rQ8p2HZoJB8z6
JrA3w/uFD19eqIgEaOuOLxGRulvtMHNrzMDEgiBmmj1Umh63w8VGdcVlntt3NPlRMOtVf4FR7sZa
JC+NE2bTGPQAHW2HwRIdU0eS1aexUHbQdTPixhWOi5dk4EeOhwDrsaGsiS3pOyB0UbwC70Y+lmWW
Bu6EtkO0SS8tJPKc/Rgmyr0MxMti5iMeByIIjOWy8BLaVL+Sf2+Cp9yv7k7oeP6LI4jCVo5DkCYe
5GMQb/eEj/fwADEWqvwIfKoJXksUvqLCkGfIYrrlGsIPieaRHqwKsgDJBgzZcM+bI1uon/D6N8LP
jQzC3LWd51pJIx5siuPFjJLaTa+NtOnMDqx0772hOVLBrOwF7pdXOkjI6jlGQO16xfuXJfLZSoC+
tFPzHhNBl3NZd8Sb6FFq+krs4fKUhzUEu98lU+IoO3p5QO0MfrwOxVCgRqf1z1XD/VREdzVEyKWe
QlyDutbvLblDfxZ8dbm+pRLYuWPbixtys3yibbUjZdKyVjt0TDXe9+lbnWigBl7AH5jt32RP8EGw
FcwqZ4u8MLbKEdFGJOFdjLVR4sn3rjmNVIHDF4o7cS67b3W3gpncQfJNYwCA2lmQD7kjOucavDox
GLLfGqRiHMHfEbCYgvabztQF27ZBMCmsJ+UX2RtXhTtoLbtZzw9FkiYDI8HZA+B/ZZ1AHcCire9c
ViYUSzuxPRQSe2wtG8NLdt+pt6L/wL8VE+2GqiA3zrwrZ06XXc5SAZVA4RzgxapugTliT+/UtOS7
Abqq1QE1FRoqy4rCi1laF1M0Y8Me5nl5yWJblB8ntVUA0M+U36T9uY1zQkXCXZoXbqhNYAYxRlqv
ilf6Te5/Bol4Ua/ab4ypxaNWzr4mtiUMttos3pjaW/RS95T+d7+zVwxjJDrySAMdXrF5gw36vvj8
ONuHuIMLvrl9UGdAiesw4xGcZ4dKDhh9yWY+TYbpidM+Ptw+0MawpLMaBxX7LJHeum5T538kGH9A
A0uoHDgDfh8d+LJMBVoAyaJ5+oq926quRSdJxzDgfH4IYa1mHusnfGAFC79urm+ZPg9rQWyqvj7a
yMou8+3rvBS56xyjOtEakyPT0HuZz++BMLcY40vr8vIV4o4yO3jJZ+OgvQ4XSBgqdljFa+6qmHoH
MI87ItO11anIad2wI6xKyjq0OkhO0ChDR92ktiG2Ywu1N7Jt6z/AOUEK3I5asg6Jj+stZtoDcnqR
iYAk6twq+V2SiZG01ogCJ5JFgLmDki2DK3zKA9W/VIfAidML33+QA7fQThgkyjSSxpv1HQx4uIna
L4q515pJMW6yeg9Xi87kxSoVecJoraTamA9ZGi7g+saymThtfPvT+Kx2QOjzmwA6noK+ia6nw9mp
NbbcgBi89IQoY+5xTOYkA0NQ//E9PEiuCVoEDgvjsmtAer1ybC+Tgw4DM/Uz3eATQMFqfbsrRpsM
4HKOOeY+wjKQ8lR/TLJ4mzzZICo//2fz9zxv9u0ucI0g66F6b9DSiwvyxeUNu+3miYAQU5mHRnUC
mpUJoqNJok73knmwLCBPRgWK8oBXi8c/RcmZCT3lrQxq6WQVqrgoWzWtaP9iUbDEPlZ54RiQ6wT6
z/eJ2mMnE/sZW8c9cCftYJwAWA1EOni/TWKbdNHbh8W/tBekFEQLtlErrjAtfIFiYH0gIDpKIwoN
GCaR1Ew/Jal6EzOo6eJpI1HbsJpiAUmH7CyT/rNyiigl7fUi3IIuINqZPOGKX5rUryNVROJGbKjl
5p6S1VHja6DiZmEwY0FW+v4uqTSknRsyKdOZQCwB4vqTtcamVkbYvu9SSnmEYpYzub5ldC8rGDWb
njdpGS3GUbPWAvKDs+q7aW4Qbl1z4CzZNQSeX5bd+o555d4fU3Z9HImQXqHweu/7LfLCl9sWaZ8k
k//dZuLhrE912pJoOw6zOzt55QXEikwLF4KfaDxBHuSGJEFS+NeSTaetSA08mkahKiZXFZtmMfL5
xyLJ3rGu3QFI3JhiQacH81zQA5qf7h7EtVEEuHhyPdA3I+SaFPzJ48m2r83l8QIHOgmj31buwV+7
/+sHluBPekYDWm/t531AD9MZPrmzEUNZ7DFdWET1VKhAXBKm17Z0Ik0aSzG4nzBtetHf6sBhaauF
D9cd4DFVj6Whl7ptEHkeDbiA5bzPrnmYlbQSI7MD9lFlbiPrAmsDbNoUULfxGOhoouFio2/rk5AD
ecFP8ANvrH8NmpP1TuJDSS7hbYTy5Qwt4PVmojm/lHLHwCftjzipjaPBh73ukA01FJbUh/ki/RHm
nXcvHYqOtH1H15yitWHteeRgxvtFFC1JZ8zl7xB8pS2uZyNhPqIp0wRjgPKUWitY58YLyHkPbd3V
krr//QtmjAtoKsVDY10PYXImL4n7GG+y1qr6BlmyNuGQKX+ZjH6mTINrAfphQ6Wr0L9ufTeRYpEq
jtAuHWaIeCPyEHJ+sLIbLWYTm19lPvBdNdly8AOyhtc9S2ryHFXbo+LgFcmg4iMG28FXUbsxUOW2
LNFmHg/LOLm+55hpKwnfEd+bN4PCLOAJlmazCClprj6xUrYNLSKAs9cLQUWJBJYpXpOfAuyYs+ma
ptTlMJfOrvDbeTFemE2zuw1RKQ+5LnAx9dN9xTJp7LZzBP7vLGe7VSKql2OJxhtsEmI6DCSYi6AA
7fFhONs0VcrpLO9tv+uo0l6m3PBpyZSDxp12otaxLKH8rTA8a+DPVAXxP4dwzTjOgDW6B39o1mzG
flG7zYXmzVZ3mBFdPa2VMj2HlVRPhT6smHinRYkgHrqLXQ2EL+/lt+vStOE4arZySR/maADNpsYB
UQtg+M3YLTq3R0DGj6PHjuz56JAHVdQyA8oGwuJlfm41CGTtc8JZDkHppTOCMMZFvjkWX72+ZW1F
meHqTQcTHJG+eOnnZvSWBfYPNHsW2rGthmlWRYXFy54oqkr9pW1eS7gUXSkzHonf2koOV1aIySkN
2kbgrXx889MR21eC/5k8+MkJTsV9Kk78Y+KktcTQYoTDhYvM0pGr3uG+UPQ8wNhThD2iAsofUHdy
mtfiQR155JqoqH8v1I+fTTSRlRC4dZqe95ZfKuH9lkuRgTdVrtf3HCY/Zpzib4c7HrzaHPWzWYOK
6DZtiEqHOlxTgwpCDH2CdVNvk7KntG8Yy095xlcSRgTKsKEkFIxnX+NSewzol4FbbNTLbY8NvDNf
H1VwQpG96KgBBx3wGZHDax4G9OPOR4GfdUs9A9oXfavNqw1vtwT2B0Jb6hcelPIdZmFJPHF40pnx
6WAZWj+gRtiXN160NPaRs3ko+FB8/xTa26iziO+qwHOhm5gppw2LVa1WwvbbdNkuAwcbdcDYuxPb
uDcIJ9ocX2keoqs9k+UFOVj40OiyiTrYDlpWjmbzOnJC7kr8U6fxDBn0zvnTQ2ELTv1N/kcyZPFs
aD7tZP89ts6vu0XVNgyCtk/d1Z8ovRmyaW/AOGXcCKGIupqhZqN1CLKdPMGs9QQBRRo5/ufToMdb
3Yd2LQQG9Tzrgci/QJXy4eLEMUOWUB9cMknJVn1W5JQP9Wdn6K4DzmzikwBZ6/XXOSVXbPtJdTEV
0K7MrcFUdCz9GdQlUUmTHqw96Au87dvKfoYM/jxoKA8FCc+/WkEGl/vaLcUyTtg9xuW6r+RVcApO
IZbEyi9wOjWGwOLcH2kN6pWzl8IJJvAxFvPJ3aYM8k9MxgUVaTFPYIr+ErmWs96xRjFC+OoRAlkS
etIYD77GSqsaGWk7JOAzQJIbRJKAb6FXFz8T/+ZoiikBHeN87p+Ed5WRoJF6Y5AbzblrW+eud1Rd
IOG2vKh/ABPdEtjkS+WpCw+lLVCoePGUwE9JiPi2oWtPJlGbbXWJV7uZ/R2KFN+4TG6UtYoM5hWQ
GY8+VoN2A3qr8PV//HhJhOEqr62t8fhk4IyT91wUGbquni1VesSp7ErJmv/r3c4u8ZbBCqmabKyy
DVXQcV//UmgoUnnMtncuHONGNzSYXawmB8pKiHYFJwgQz88A7agCFHa0Za7iL2U8V/kUWZBOi8qy
dMgBmxVwUSbXHSmGJd3NWZcyQavrGHK2FcBqWUxdRZjobJA/ImoLBtKCiG23QWkUiZm4nk6oa4TR
qxoof6z/T5Ww4BguaPwhZNTBKgbzNf+xeQ9oPuenKFCfEWx3MBgB37bKa70iFmPn2ixlasIImpLr
HKvY7vq+5aBJNU3rY/ErONsEViG4fIf3EsO87y9P0V1spZy166eLX5ttAb46Rxj0k0Sp6yPPa07c
oWsci4dpagh8Y77Lp3nPsYkMfIhdKhZsPS2zjvy05bA0pHLvez/ly125l6tgccbV5Ml7nHxBTJ5r
Yv9mGHbA0e30SGaTz60KS2R4H+2o/AxHXlTj3Zm8tNSSqui6p2/LJYkeTwN4oaxA6NI+uFEcP8Tc
reqwgGIjUZSC3sCJ6f/paibVvqt5ARF+tqnqMLxWCFWuzdz0SG6GimHBo6Fck2IN5GIloBGqnMzA
FLVIycQshnBOGstEL01xShmkdPRgYfDwFzxxUbLe1U7CjUUGj8ruzNRUGcT38i/c/3zm9D4/yywV
0Cs+Z+c+qHjJzEDi/s3nv5kySV3dh/ZHLprzoFn47HrhwZsvrcOpJ9Ptmvnyy8EMlR+UVTRnaQLl
Pzkznw+AmPl+LOcvqASE6rjx02AkOOXI4R9XP630vEm6BiOX3HrkZPuqLKQsA/M4Tv5zzXBZlfEH
B+uCQ78DljS02R9WtDLtl6Y0ljcQ3dWKvLpkw1vKPzX+5gRgp2o3ANGZ3c+0AB7odUcw+9Piw/qK
5FBIGvrVOMm1aK+RZ3aigPwVWqr62BISOuQ14qjpHPSJNvXYzQNIq6tl+wsyuu/K7F+j5qDFRoEO
HZke7zLv+9ccC7BiNE4hyoN/mBEZhMvtNjwXopHWTqPPsLNp5N+oxLVVd/83/cTByoy3UM1kPa3K
+nrD9P4MikyUueGjzBTUQrsQLTJlMluEC76RkU0obtXWBbxd60m3J0YabyufZAr0bJ971JHm51RZ
FimStR//4RIulELfTuwETkNccZfsMr4G/iF1yeQ/Yix5U74/d0BApfKLTLzCc2YlYCBICQqJiqvH
W4I8/2Ck75RUZZCH2fLv1SwvLk49BU6QywKeUdol25wkKj748KHOZKH5kLR2Nn/FjAytcsQRVmiO
nat3Gb1PxwGPltACVqtAQzGuyOky06rg/3KpLde939eLi5lJIUzeQ7gbs50YsEUAXqbQu6BMOPn8
vt0z3yCgQvhGdDWFO1amrbgmJq8+qjqoCgqWMY3d4+UTbJeKoVWxVD71m3Glivd6pPxM+hf4fTCv
9c2U+lcgqllYJxt90OMQDL/y95ILPgVRvkPY3rHDcmxoc/NzueWGiyYEjzuduULlGl/XMSnHIiry
9cMrQrtMEzUkp0GcFCsooHfBx2MJYAERGtihyfcG2ZPoyoFOOrL/ocKjAV4OcF+AiDEQN8y6jmZc
OqZCmVqeQLNnBI/4BR/mC4vfCgVGKwXvKtVdoBHxYgS1lAazZKpNqIGy2TN0F9T2u/bnaMJ0tvBH
NP3JXYQ/kQv0VNyeFvG1uVKxrBZUm9StqRk5XpOsGFhtFb75ZKkjBPvjvpBK+HaZwj/KYA0bW9b1
kULIk+NIFqfFFKMNFsdHbL6Pl4Z6IGYfOxgdpUHFlVNNHHEg/BCT310+ewHWXHukAmUncYekFT/h
A/SplrGEQgblFwuIxwPPwF1mghmjozGEJfcTuTByVleOlUPWYAf2uS2TbDO8DjV9l9J+hPTEelTs
BsvXo6XURB0GMadRYme+867CnoBmIAyrGK/5rYWv7tx/xtXZcDc/kbOVxrGwEpTEcs1CchGynTdN
yJLHnsanEI38vk+nUmx2w+RC8l/qNQ0lu3v6h7cHiNTfnZDoiNmPeY/wYCaM9ocrgUvNYY9U1I82
qsKRTdKxM7zwRMeifh4AiKgvwgAynl6Pu7IRVNtm7l9FHNGbi2OMVNCtDCubNRtZlcSCWRofjzjq
8AX/kDIWbwgx0VsyYr4HTJuwlCpsCpgF9ibh6TeUuT6DqdRX346W9NgHI1np6uvQRaIo/z265EkG
WtKh1UtRfm9tCv2sgtKnAy/gyJcX2Wg7RU1Rjb1oFXt75CVPyoBoHffZrpQgGW87Adfy832lnihx
6kuzuyHYGfGUQeiCuxDfd1q7GLIRjgjv1wMTnuohMvTEYnMOgtiLrEFSbltBriiFkKx2YlDDYNjA
zZMo9C5Nh1/GtcFY3pgUecrwJ2IQdR9kgFdJh9P48RSi/sjnkp+vtJ+NMIv+2U4n/F/GAHKwLwBA
vHYg4J2Ko/8bOY2RKonpgVNOg8Sa7CUWoykbAqeiEdhztx6cxhn6c8HfHdOiLzxVVfhfvJk9reRu
g866IN9nyvE4cRU8C2HB02/jogMVFsOEv8ciqU+NYLPNutueZZFhNAsIojJ+Z1UxD8tK5tmUMMaf
0mxgftmMw5W8m3RvdaZ7S2CcLbsNeuddLAhneivoJYnNPYE12HMlS8VaNoQJ0IIEcFlkSJuVzhya
HeWxDEHcRaWfissOCnf4cAfO1yfI4YLRhGwCaxnmqVLRQ9Rg/ymma2PNx5v5/BgdwDjtS+QaC2kd
FT4Ot3mie+xht8SCPbNTsiRSspH4XbOxvg8PDb3V4JUtPZXZ+1jvARxDAk5jvbaKeuQg+zJI4hgn
mpV6XwcN+SBJWu3NALOv8yIPztMTNj9HsvguADNYrjvJH9LRFrTKdTdKBdwU0IWROiI/vzMISs+T
ybi6x+1a7e1obbMLIPVEfFdQhk20izufWbxZXKJq6p8gLJ2Ucw1q5ZVc9cut8sWk+Wgd/8SZzBrM
ApIDuO8m9Kdz5vT+xL+9z+kWvu0pgTjxQAIeXdmVlLLpWg4ruy93LpxudJQgj+CH+2wwC2nIq8Rk
pYF4DtGN/W0N/bsLkg6DKvT4idBwGdZLhu6AhmSunzT9iHhJbAjFNjbJpXQf+zrTtIN0BIYBIFGD
2uMBP2aCNuDIWATBkJg0FB2YksCUUdfcuuXUDTXFahceoQ1sl60PYYZnS04aX78/aA/oTLZt7jpn
kneLdvZc/IgPu9gnDeBbMfAV8VGr9WGA8SaKO9kVlzxoKl4OV+ZcSz0YRqdNFyagxPUp07a8Y2Rx
BuoNK/hCHom1grYzF4WIsb+hUd4skGjWEKz4P5Z8KEcj0gwfnHJWtDRrMqil7JMYT14ei3BqkiW4
Aj40VHaBt3NMvcZBBAgvhWu/IwCv5qXEPnsUPYm4N1MvnFF8RomtmzIIAKQ/POAb63zT+WBDjnfH
0MIcP/VY1z5hfcGb3obyomYHnpor3FAsl0AixPt7Ro084CC5FobascPPzgCFVcAkS3Oipbgmjrwv
D6Rvs+V0IHCF5+G/IO3eSZheFxYL40j03gFMATyyTOK7Tw6o2OXGHo2Oxf4yd8/w2Iy/kOPJXQ25
IRAQFTu463Tr41c5yphwv5rt5xOKnwpmeO8UuDzIfNerWtCXA77a+uQbo7be0hM9TI/e7EEQ7JH+
HN6bA4VaXEN0uvTj1bExWyT6zZkF1WTvB4XtoHT2FoLb0g1/Tm66hZsxIR6kl0SbNX7YzQxFr7P5
BR302F7rt80Ukv5V0g3a8EmO3NAf67Wlm9OVKofIWRKPEMQkteL/ZHfo6xclx9sYKlBNvciosq6+
Ckkp9gtUMlcI3+f94vo/0YteRdZbTgx+6cFzbJFE8aMuO/NGhq/8VUaecKdRKPRTeJ6u+Bg/KBAA
Yn74IB6QL/D1kFiSNAPD7cQpPRkdUjDf7Zts0XFBY3nWw3KJrvYAolT4bhTo2h283MGeHDwUWlWE
IiXD8kIlMhvdVOPNjpGiRe3Xp6EoUs+tG8/XCjJ6joZCq3ZqsuaKAPohXkC+dQKTbR3MKqDDaLZe
LkRnBT6GT2ZBemMWGItOHgBlMyX+euIyI1Icksh6+w91pIpaQ1uM19mP3l+x39HEmFVSh7D1ps+A
qHev0VsyzOqa4b/MlshJW1RUOZeeuBX8d/tNLE3/2zn5Eu+I9GcVeWHsltCdbOxfWirsul6PpIzO
bpLT0F8ktGsZBBcWgsa4IgJ+k5iScu+TLEVM7T6WxHOzwTPfcIieiWe2AtQriPsphZ8BtKHFpXoz
P7xisA//3LDodYJmdDnQSlN7+7HSqDgFh0nxMTCODLJkC2hfLHLpjLcHGZNnDPAOqAkXm33Wa5Q+
wC36hvyMK0tC8ex6oCN9XYi5KuKzv7Nuxdj+FntyhjcuSXVoI23TXIlLNLLWSsisgPVSZPBvX8/8
/MJlCmodx+x3d3vm4Bp1GDFwk88dhYPN9tkGU73OaEooPhNDuJewJ2fceln+7XuenjVJGqgdo4uD
RMGzeJuAQ8v/MGu73bpJaDOyIEzcxzwjL16vcaYCi4lgz/vX0yuE8gzPtRAMQT87/vVKIDbmDPM8
K23lUyUhOYFakqHcuSrPTZEeHjIpdQNNEDC6wJsbRNLfqkhEFZLs/HBio267ziN5ksEi99dIWVvJ
WvicjGWNbLyugx0UFo+lPtXFJuf8KA0dqviLbKZJKj/R17OJpz6uvDyMuTtUqAQYtZ9xx19gtEkO
KbdZjUlh/Sihvif/b+E1KOxBTBqFOrYOf4arNPokH3VOZWy0SNbz3SJToPMT5YGAiASKXcWC9w3z
buKo0eMG6jzuvyK9zl4mbe2llOmtVQ6XlHGaTTN2Xd0JHFi+xI4U+ywkXVMrzokPBr/m/amnSok1
v3Z+FcHFYOZ1ApAoWqfq0S6mUBtRTxhEAu5wolN/g1w5FLnp4fkjw/U2A0Q5GWyb5eADirwNGsdX
EudgOuCD+uy414B6IcU5HTpW3oBtWR0RfgGAkJXzTEpbrbJnf2AbjEYQPSrKeLyhSAO86W0izlgG
4nQLnK06uE3HZEUYExJcnCq/Ci1GUzEi8aICbnyiUdiBERKHxoxql1ns0RPwlyML+qj4rzEUNeJ4
sJxrmUE622By0lwx7gsEKB7XHt18E4j8S1lR7EjqQSxUtu5SstvhnC6/5s4BX6JVBoONcEScZisU
hONc3CX5+rARxCn9OkRxROT1t7JM4C1epaODsMqv6AQa/bPLFR60XAvZQlwCnXFK0XR2yPCYU1s2
Os1je9dOUxVaWg46k7mcYdb1yDftOoPP+ktjoOSyCbYVisYBi2Vniy0SYUakIYqY+s1FTtUIVXw2
xkSf0VVDmuGlkGj2XenW1BDgSUrjG5lCK4jNebZgnPyiyj/VYksMR5zuykIGyZZoSZ4p1O6WhUG9
9+YsmrbGTlPdwxcULJel1kQIcabg/eM6D080Gi4qPxqZ+kxo0DjAarPlKX5X+a1QKIFUHwj0pjyp
X0kBh8fxT1EGhbMLojr6Ksp5bxebZtwuCzl7agcHDkgSoEr0hCbMIpBRYrCt3oKcUdpcL94uL6tA
fGjyvRp7a8LAErVNi9yWGWMY48daXsYIacuLxLpGMwkV2SbiWbVftfvPDIIGzlhR+4gBCuhwQ4QI
FvdjvlvwMuO6x7kEuzlHUlipTAo1Rz/uK0jLv14EZ1Jr8nLHBhx1Wh9JhXTg0SHSHFY6/btJYY41
67acNnJRoX9gwa5/wpamoASjb52K7dtlnZSseYA0zc6+inuFXe0WyYlBpclyC5vb4FNBNSIXKanu
dTeOPuBo0FQZOSwCgVwbtVvEYSV5cxKWXmem13MY6g5M3Rcq34JdXa2dphRPoqMD7v/nUtZc9/Y6
i2EToTdUr30HxcfYKE0So6y2AyVK/HmBEpIyIHjijVcHrsOUuSJ79sbAiXkgOwl8h1zZ31WR9qny
a8GzXXaEZRAX0xwYNP8ZngMCmul7sRw2DD7RTRqmYZk2AYKDcR85w9X3mytlVyZ2goxIUxmO433r
FJp6dHnDWrt6uHVFai2MgkySbcmkc3VDf3WgPbeUYRtfJxtLQEqqEbwHu9SY25nfSinvrFEqQR1B
Pqa28ZfZPtgUfDaI46sB2FnFMzYbSzIx6z+0v1hMejjuS411pIHkK/+CwiaewuL+UkIzXIk8qTYd
s7bzXW6onpckuA1D7DzbjEBncjZBty/lOjhywtM4UVEWlTHP+tzjr37rSWmkmq3hY+PnWcafppJk
36etm1HC/SWCLxFKYGPxqrY7htgGfjlkuZxc/pI0aKkVDgDzErbzPVHU+FXGx8GQG5G3u7OtGPNp
xe0rY3myTy8tFoVfFN75c1TZSiqPpPoAkXmuTk2cAmaHU4JTDQGnKoA0EcTTgfP0ZBY9w9o13bht
gmPc17JD/lTzQ0wHmpKcNJbRVYpW/N8e8EITQV5cRFa4nNpbAKYT7/nWuHHnyKvS4I8qnfuNxEif
ds9hq3Dp+8W0icqn6tlq5I2uA6Z3A/rn5l6WGPfDXLwv8M4NdnRdzf/o5ffh1vOnl5VzUvRyC1bY
VFbdVROGR1ZXPrJVAENNvHnDh41s/FQKGcM/UktFW8OEjl9PgNo5GWdf2kfMEHV0EjGA4U8uQJLK
uYGiJj6wksYlR9E2FfYAARHEKg99AJ7iBnJQV6DpLUHq8ZSA6r+bGb3Msmv2gwsu5nDoivCpEUFT
CoUbw4L1yKar7ltdJOultIP5OmYQXVX6lM/2V1YgDWAk9gLH3//TXIcum/if2sg50nra9NBIk/Nn
h5z95SELtLcuDezwIVhvWIQlqEUKaDpHxhg5Rz2XCqZNWbTtc2OqiUH87OidjpkKBjH7stn4Dq4c
ZCaQ4V8pnl+a3+1jQjUrRgGYztIn8JSvpiRtyLb07OTC+H8EkSQBzE5MW0skgjLFyNFUnm5mnkB1
/AN+DnWC5AQw9D+I3L5itGBLWY0ZMWUsPaZ4r/gw8WAC7Rz7cvQ3SD3pVBAFY5+YSWxU2RT0zY4D
sZ5LN4By+owU2SC1LZgsdn8lAmKEZysYSn/qW8FcW3FpWBXsAyXY3OSKIJ7DqIbF6dRL1JPOyfKr
7RVqVzBalwIKDqOHAbNl5LFlWP93BfaUKIQh08qEty+nrDTmnLfV2dTs6WfCfUIWntneukKvaX61
s8jfid/CLxxzdRvtnOWVzEjof7OZeIIPSMEOS1isUR0MpjEEFsBK381x+CbL2yCKHfiI78cZRXPD
1rdzj1GPfZklVDd/OcEPlyrhMYKutKV2RIxaq9vnFZrC9QsFATnZyccBftPczEsHda2oaBUF9K9P
lMKFVCUA94NBSslcKba+mAvlhdqd9Q4Zbtni6oXsJ0CquE/qhs/yKR8jmnPUpksCGbWZLNkrXGvd
2Gba4qFhNASugZVxMkY25lRHuFXeFb1MBgliWCvKCXZfIHPYTJatXtSevsuHSHXAyq2G/VtqFfDi
CDR761ul2z7KlIhSLvo5wA4Qyd8fcDrflr7QMrrgJCuyeUeIN6Dg4eVqClYNxFe5lmu8zMkTjHDg
e6gLMYy/vCciVi6ba7/ZV/YPTrEqn8MWM6PHp+kChMvfMQgFNQ0r4BmqxWqi1ngvAfq8t+SMi1z6
gq/tJqmWcZlW9/SRqeyIdYU/0yo0PUPrIMCvyXWPUe/2YFELpPrcITvaszssqQUbnLpi0Zp44J3h
R/8PRYuVYOdeXb+k37YAasRxJ+rkpHpJhYrKL3SBe3x3TCXwdy258iKGrHxt7/mYZgEsxApGVP/H
/jT830D5QVq35+uh/erVrKBHfuU3tWVzcFNNEBnG8CPfKh9qNq7yghTKVSwemMxQiLBkrmS3AKo5
WzsuE3hpx3+3VnlRvp9B6zvPgJGCFygnrRKklCTJfn93q/oCAAcNxze+fLui5euUyH6Gdu7AkO3Q
sC9ov+ucW0r27PRtmZL9XOEevpBVmBQkUGtb5laAexY4CrNYCsMoyz8vYX1J4k1uD9LJuk62GGYA
1f6pIy0VX3vm1v/VT9K4K2bGl0hLzNcZ4TBeEgL9T0Nd3d7cx7p9gbZrO/oai2Z0jeie7YGWTg6V
3pnc1HNM5LY3AWGZ82rrLsJvrWt8KSeXEAXPPJpzPgB/IvILoBiYoSNzqupxBVNVSabJ6eSgl82o
nIXLCgxO9xV7q8vxNljproeKV38JI3WyUp2yLeNMA7nCrTw497fx2joF2g4Kd95TIQFBbp5a6HUl
JylLXMy3085zWNFMnKqg2FndtdNlr6hsnrg0vupIaY2LC/199wEx8zZpw4XmySttgGlEEahX8a5Y
UeolpVg0I8mhBSCuFHm1/8B6oJ1wOKrbRnWU5KH8639whilfJyr94xp0R0zEAmLtE0CHh9zewuUk
BmaIx8pmJMfbS7AHKaqAJOhXZmZxKmkqilYw4GkQV5a/B/SkOpt+hrmgLaXQdqHpUYDbvt7bdDKh
hj18uDBlvx76uYULtYfeuiHR1iUOb040RVxoGmCns82/wBOueaaBmv1V+3YsQnpFNoB5LAhgMi61
VRER7/0czRw+AI3poNOTU72DyeDNEwy4s+aVj8Ja4N8BUzNKNfcnSDmpXdQfbqHjXnwn6GLol8ep
HpqFV+tP2sJO46DDo0MjnhfbNvTDIfeGoP/+THc3b3kwcDMk8yi14ghE8pd6PS5iNGBDJZlMvxnZ
qtB55frlf0YHY9bilr8azcWF0TqweWIwUcdupQ8emWYvtE4AnxyIcWgvbm5KrDKhxAVUP0aI8eQj
7TCfLxZX8iu0nvvxBgHN/13qsKTdxrYLzNnwk1BntJGAdbNj6PJ0oUaAfg3xmAJGN9Xep256MdPg
zlx+UK3rgbXdf95vZ8UgYkRx2N98Vf1J4w6OvmVj5L869jO2JhUwlp+e01Y9X0pl01PC9yyzirq0
ykKUql5CrzSV9uB7upj7dG5ThYY/BYmf154Jvg13XcJc8L3e8QqOBmg7umal0lukf6W3gN93ucBF
uklotT42NzmwPz508MCcdhpuXyUkINX5wO5lctGSKSd+QrxPmB0a9q7EMPCEbgsR+5/wQ/jzH4D4
vpxCX0MPnoHl0U48n6RGtrSareps0LPWkjkaGQZi2tjaJ1q5rgKj0qQFsaWMTu9dnu2khufzdAYt
kDbFAQifiLnnU/qefFNolgmI7bHST/Y+xWSLWtIhaI7U9kquXt1lywpTNyfZvYhiiGqnTwK7leqP
eHSLigfa2wt38t5Qi4Q+n5JVqzjd61iDGbdJGDRC52VPzIminEeUeWcG7gLrH18z/v3LgnLMte4Z
BqwD5l08Pt+0WMOBjjvHiF10xOHKfVi+GT72r+bGPwMNRSXfOBEKgZadopd0JR5dwt7Dqhpb95mG
BySJZvEcZjhNAClAph8W0PZPJ2v2pNnxiGjX7EfJJa2+ZiyTRH2V6fY/nqHZsNOpahA347AXa6SU
0BoIonuV3vrIRzztGXRU3KbND1wwaK5nAPnXPCyUminC4NfZbTqnlOWdcq4jvO/IyOkIvXToE8nr
a5cuBRL8SzsPxPaLgvsACo1pqzoJUyxhF2oKADihubpM90v49/7hLEpaSi2E9jgc4jeUI/PSO4xz
HtTn/zKf8/Ig9WO64X/tEuo7YKfNlC7NgDuhLtxE74RZDadt7JrFsbu20iZ2PuJZpC7nuSfWz3bo
CAtgc86bz8RAXs9rChMRQCtlgEQp/Qr0m6d2XQ1B/5+huAnfknTaaWsX4UPSIyXM5t8KOpcrrHcf
Tco6dZ0fPW4F7wIGicAlJx8fQrEJi15T4u2fzeiSHJY35Je3TC18cbe56V+zkjGKhYknW3YmAEc3
EtoSMJbmRq94GmLcaTE+7TncL+rgtPWx4nNlnniJRUbO1S4clewmpJ8g9CnQpHOhufpWzA4XV4BK
ic6K7E7Im1xFLYVu1Yl80k1390YJzIlpM1E+ZpUeweT7MQXZDAYZOovtWmACXjyUYqxcM+0r9mIF
cNOwNRFCGYlianhnp97mUTwiDCkyxO66nHIw9i/fs8ulxGF2lf6x7WbrciNqHSSjdHqp2i9/eH7g
C13EmJ/wqPq1iOoBmXHGmC1pLD9x820QYR80VHDItF9oKnV685KRyO+AfGrb/9vCK62uQcQM6vWZ
cc9aNJtcxmdcl2LJaLzhv2pswsYIOFWVL0FDELuIL12pRbWZ6mzcIj7MaaFdZ5MjoV0cvwOyRd1W
FoZDP0OGkbeDLnUGAHZ3lkJAA1aLcXhPk5H3TGab0szc3XwIvnbJUgkBPAvqBZZXEXEO2jtGvvLH
cTjXGtV1JoNU25s8Y7jTetS+UdclUJd6GDKMYBVtNG/xHaMDvkVMOh8EVoDnMV6SR4Qk4CL9t02d
2GnYYLXMFOqgKIFuzTdZx/xlS0wim14esSaCdpWVZuBd+OlR2ER6hVP4soxU9m9Edz9pfXLjcyau
ipuYkwGD0zQ+ZLGa8/PKyBCvXgzQDq6+SvOsLBKHtYjmvmClbmdaJe4HflOImxCxqIII1EuNYxmD
41bmAx2EViNUEd9PtuMM3P8ikhCtL03BEAdYjwZou1dgWd4UocbO4iY32yb6QDdurYChKJd7ACRZ
J/+FUwvkDWQ4r9OqJSUY4lixzsK7KZti9920C8z/o4dINldPPqTXcLeLNjnBiaR//RJDI96Uhfw7
o31I+VH9+u09lYKwdO7oU5Gihia2QBDr6T/pA12scCWAzmVN+61QyZvQwhWRl4VjxBAs0xJ+3Vzy
WaEyns73PIiC55iUyhK21MgBsqvjXLNLRDEfJRXYtj/jP5Xi2nrAaBQRYoNmMvEO2Nxm3V1LAlnG
M94t8+xMHryLnD7vrb9qwCXaIti0BUl900iGizFstg7ShlYDsuPuDM/5dNdRef4scb+l5a3HROhG
PnDiLYg0WQmJtASP5W5y3E1YeiHIDNsgVdKWM3jxjhXLf6AROtV7l0hqZp+A8RcHhhQxKW1+3NuK
2F4Rwhicjei1t6Xzp9Ubc28/BkZYrXWXsz2aUbPgJBA1KaWYmFWOLDs5RaWuSMeIAebkQ8m/LfJq
q1RYuvPQJ2sbyuSQxJNBnvMOeg0dwUeECVe6sl2OUpB04fiUKVoyd/P1lg7dFS6ZIWEcwg1lRlN3
xJyygcFRx3igW71LkHWyzYPn9WccHXf0tRi8lg991p6fOBEfA8+SvsG7M4/1qaVC7aZzPzzdbsqH
85ViFWMZKhhjyDuBpI+pand1EXOVAZssppAvej0AwScXuw6f1gmWrNqhAYN64xHxZVfZn3EHk1cK
7vWCNRE3EzGddkbdRsmIlh4K+Q4xJLNpfrVsSq0MjPEqLGbteOJCwSXRQ0ECyL64fxD4yffbVAYY
MQj3vl5l+zWd3SYiTAaI+EEf507PfMeeRt9xJcxLseVUapLHKFac9YIbLxMRM/BmSJXJtuY22fba
B8JRpharwKnyLsxfMqopx1wHnHssHbmA3WbnGFbjxFYguEhsCPbkcTAr69puQk2zU5Um6IR4DbcU
4ECWJKf6V/JCcX78BDmmkmpB5bZlDTwyUl7nbH+MYSepYtAxtGYKbB1dh7TzHQzjEi+g3WdLDkXK
8VHtl9iYD6KtoDud7njKaGeuIv6QDrYUyZ7buZ9+ZKdomcmiGv1Rfczg3l1mXXmO7DChbswbH4i/
IpQteflD5fT/6r/u+b+xyFQCyLN5wBKf6wqao62WUgrzXChuGniwAceDpb4wDZ50ECapHuUdZCtY
UfLbuuiIa5Oq2S7qtrfgKtA8j0FgBFX4bMEErtgLM1dSNmP6nDFcL30ytLuLhModnEy+zhE9telv
5dRBmKd4469ehXr9FB7EthKALI3nGhRMJvnMp5J//5yRWs/aZCOWS2+pulEisTYSntvY2qPE0ert
FDD463T9xoIscHezxiwQN3MMG1Kp/QnU4gtIyoSRa8ImRwLdmCnZjpUu858DiaXNwZMEvySs4pY5
1tPaFcWX+bhwUzxZ8qCNZ5QbHE1b9RF9kLw6DKn7Va/TXjv0BF6NY2hvxY95IKcuyuemasBBJRky
5itu3Anf3kixrdS27V2ZNlAAkiVVGTfjdfJqW0l5Qzdj5fRHIvEpWPMAhDWOtKofhfVFle0ZJzj+
7ZxMCsxIUJ1GxTZBKXuAqdz3lHyHeMKqWSBDYCHeUPA/CcS9eC1UJ5jwfaDiASrSEbVixF45/QyO
HT9pm6Ajc82T/CYxS/m+JUhp4v2wQX3sK+JKCS9pJtAf5g40V72kznwimjj9rHk3N9eEqURucsYV
xPysiy3nqukumD/j2WlgrZp+8uWwBgU8zZrZ2IyoIDkADLN9cwl4MdfEdJ/pk48DU2MMTHD4s38r
bgmMgOwDaAUqiRcPZsp2R6h5LtPlyNkwQoF/dMHZ7aD47el9jCHTU8KJufLCXNfvPCiBCwWaJT0O
qgO/xxBbvWMKzNVZTPzPrUJZAArcBOK77xC3k4XS1oTaGgLBpQSoueiJX2XWXXdRa3yWKa4jttcC
ymBXe2uUzGiDtYmd056gcNUC15N3SY7OL9YXPtcxhakVQ2fYVbxVl8bs+1Hq40UQtwCxUSkbnYWn
d6mWA/yyHCnMWsjHlpDmBrVnPYGbsX4a9Hwqd6p9+RoMAD2kIAGrDDxVIA7SxaSSNtNItPsqFAwa
lAMqZNNF0uA6FnlrvCv2+wDUGo18d89TSHGJzdQUTS8XVz/8gw0jDIee4lm5KgmU/EIgILkg7fSK
vc/YXUFWdfJumiwZzANHVvpluC8/PFTntj/s7hYjy3AtUIxneQRFOEKztRf2gByeE+MWI1NtRFn7
djmzd3T3F+UhlRzuDdkY5So5r2evJAt7Tq6Rn7YAdpWIYSLZibE0Nsmm9zwhdJoHFXZGv8rVZbqU
+j658EYaI1lF5us8GwVIDc7D2Fk1ntOVtlTleO1WJVa8L2rMSAA9NVRl28mjoT0PIANjaFBZIY7p
Q9Wk7uakWWMRBnoWsxlonerrd8ocTNHzlK9E9WKNEv5I3lmXZ4gHH8KpM1aRL6KAQv0sd5gWPP3P
Ji4tzvGYmZ9rGh9Fza5qE74DSWHl7GoqiRdRvmimxKlicVF/ISsJ1ZIxQnLHQx9cCxtDJfaNnatV
tL05Ha4PPRHnM5oMWJxH5uqc70WtA/cQlp1bZhCIGZoClQhoc4m5jQCJ2VlslohLKWptVxziQsBJ
IxielI5n4UGHFA1pC4BY+JqemLPiataxHq4Uj9n5p2AlSNXoOeMeJWxdrOMdPiDB82N3QNiUw+wJ
66iYr936n6Qw6o6ji5Zhrqk+91blh94zwy0ZR6e27mMbF2dMyKMt7z+prICFyvSKqGxaZmXpNI4C
8RLjhwXnn9Po/0c/jOdsWXKDOmDJ4znD9eaRjvOYUGEEjz+GMOGCsJDq9HAsRKrz8a3Qs3fItPN2
GnnJgIqH0z6UNn3LrtkKbQa84SrAiioY9bezEamhFLD3lAH8/G3KLaY+6rIu1fSH5FHvPhKKPVuW
G/7hnHPlXDEIfHLG5Gh2CAOaxCkYLAHM9PY9sxD6525nre0tXwSX6MaqtY6RRITTOob5KmQJL7T3
PvVUc4cjR0CykiNjtFBDZX7X+KcEwa/hn+VvUNZtCmGd+UbQms8aUa3aFSTJYZwnERWGXutrOh4A
a71ZwCIYAkdEWu/GsTGiMiWh8VJUbBXW/kvntkHkJxN2tEBTz5lfocPKvNsFS0gf2JgbXvW+gbNi
MtWwOMi66Pm7bELrkOCLbyjwd5fmwls/3XdO8FfpHVTyaf3rEwG1SHESjXz2bCZb/XlzbMrhBU64
aqwNOUtyGtYoc9C0/+QCAISLw0z3bqhfJwEaSl768aN1aZ9zTKDn8RX3g5TXCotTkELfVwYtnZRI
HVvSnboitrCMkGF9BnwbymVRwaNZkmWrD6ADaGA3XJdR+S0Az4PmRtj8Kl54XXmZ0Aa+tPg5ilAf
uMUCpjWwGgITQtQGMxRSDsfuFc9a2Mw8vkA19oKcGVqOf0iZGyNEc8E01QIH5ONbPy8MyFfAhUqd
CfD5R4yUVAuf6ZxX85zIrVuaKmnpG46manTU6sntpxug3/TZ8iKNzZiZWkpZTqV3/N56ZuZpLU3P
AbPE1kCNLGN+l7bGyaDu3vXRFUSqGc8m7hiLgPeIGvMjZkiL7fLatHw4mzd5d2s0abddx0BrBa04
6P5+0Kt2brR66ocGvlki+yiGJA+Hpc1ady/0PKtwclZpQJJF991nHQddvGM2663x+hjDOofFQr6t
hhyJXMMWY4LJn8i1tCgXAt2QDQBbfvi34FSUYPqX2c79QsywLlo60g730dyftVsXImZj/TvfEoRx
RwFbSszL96zrw3KYL+75CsmaNChU8ExLBHWs8lPXYg1RnimK4FGFN223mVlRwGoZUaO14BrZz+uL
Tt/sAm2vDDNCM/2S0gHRhQFqr+Dv+WvOkyAuhjMwCMLIR/kgP247Dyzjvblc7VTnVhuBxjEFUXn6
YgBVollWEHUhIZT43OS5a3wRhd+VhU2GAzv239gy9gYXjAAzaApUSdepxqX0dgIzKw/DITKNBlyc
2jXOfQX8N2JMgVrwQtR8rq42+eTq+Y7bW/kfePlgzZh3w1I1hp/0LoHryBxpbk6kXB+Iqmp+xHJ2
5mRUpKiW9QJDQRHhDcEZLyv78+xsF3nSSHrFtM8Oajnvgb0lBMnxqM1oPiHGnmD5QYBlQjQESl2Z
wtROTSPb8u6GMHXSeKURbKHZDvipAOk+a0W9FMjzMavtkCwNnnm3SFL7qJdTMjk8nG92Te7lu0Zj
NuslhJOkrh3NVJpV78iz2c0KJ0i6at8TAfuAqTNDntAbV+1qt9eCRr+RA9lkPhS3KBKYnyHucw87
zruQxW58RxE4DixMLt1oDeij1Vj6dktlplC2Quh6BOq/zWPivdE0ih6fN6TWwaulO8eQ5wSDH6Tz
2eP27bWLaB+DwGasrrvCuIxq9SFcFvlOe0Bha5x11LRutA5v+oVTYcJwrYpHE7Gi1IzZe4PxRasW
QKzMUH3r5QoX1iZe8Z/6SepPJesV/JZeO41RB1CkCkCZi6FgP4r+EiEEql/HhbA0GEHD4yz+KKbC
F9gg9nIu7fZZHHNiBXMSeMz0nHCgi+VnjObWAI5hTTPccHPvL4yfpx0ckdgLKnjQqQ6e0u42fFI9
8wWvDXUISFy6gBrtjpBkiYfHI+R8Oqpjdk9tBxuEaJx9QuIuD8hSSrmRcgmuCsZ8cEB0oCRkcjGm
hdadluQzQ4B95Xl1P6tFcpVB0lpUMjlh3piBZEIMu0wXpMuryXld1Kg5Kq+cuYFW5nYmQJgyPlTQ
8TYiCwS77HKZsKn4AQRvyoWUuPSZ1DdCxUMUTaGwkKguzRv5N3ybSEt/g3QCSploGqSykz7htWHu
c5qVG2F8rZvuRZDJS/kdsjkmeS5+k+MbYSbAfMAiBKYUfWKdQSfX0r94vP5W7iMcBZpbgVxN3iy3
/uSS9NWcV1GyyM1FhrOCzY1Oi949TH1LqYUO1o85f3ZLUzsge4WXcuBJz1NFH5njfaVlxUn0nBwO
EvyPw9MKBtR5I4JQhCwGWeDxeQrkB7/EdnIiTUFujfWHRiIGjiNUuMhG3hcC5eiN1IOrBSDEeX1m
VlgTFe4b82m5fqmOli+fEYQgFHIHD/c0JQp1cZ1qVMUMnon8tduSorj9B4HIGCNQNIc3UIU02tgu
B6zDZSeute7VeEuLM3Br4lU+hq51Vi/KWtV8/KoLq1ysRAAKdtpVxS3QAzVw+os1tvGWqvo8notU
RSewWC4W8PPm7IF59Qlx/EzKZo6TQ7rAZ7k9JPudm/+mGxb+0BTGGhjFww8z1A8xbJOmnP1Le1NN
ZKKRnXeI5U7xrA8EjNxd1xjPpdr89D7W0PvyuF88S7Ek5zgOZZpXJKggfPXTlicXR1V86YjOWEmY
onfq9YaCxEa68Pqtd9UOTIh0KHbq5YR9Nth1gd9rrsCA0EZrO1u8PCqghE0RQ/Iif6LsQ+09JUiN
QIV+/qM9zzIdgu01bTyYOvebtQitKgYEkiR1sFQtKky2ISGnIa6FCfd+l/h1agxfvb21ylk/iw6N
1xQzfkvzMNL16fHOWdV/euT0X0mMW8A2kQ8f1KaMooy1jGCv/kbOT4aF7k0gj2eYCtZyf5iGQM4H
0LhhSHRfWlQfUQKJxmErCaU1Wq/T501EECB0JuhRpDAnjuvWNLQU0/m5ckl55Hdbbp90xigI6ye8
bu+lGk23I/p4DWwUVhtDlVj0jUmW8nBlrW/1n7AHs6T7KiqeAH57Zw0Vd+5m266AwUETQ8yCNhrU
3oe/fMrw2993W4FyDpUJuqiemmMS1hLWRRxjETyholk2vOk25Sr9dbyNNDKFmFGPr5GEOno07BM4
cnTiT0UP6Om2jv3p/OGd7sX/s8A8NgOk36c9PunNwIEkWhg385T65IaQTCs6wVCqiwNwXycW9gGU
L0GyDBPy/vcuSGvys0RZ0xDScjgnn6tzaufkfyEgsjjk28fyfR2RtQHwx5WUYk0qu88SY7KPB+7r
+yvtQDY8efq5nHyDr3UFhdwsAvoIETWn+4M4YhIwkpqpU2ilj5iIg2jZXzwQAeItPUo1R/gOkTWj
zrJnUNLxijEtRxxkNO4AXnBN2ok84RZctaQ+TeAFB2NDI8+2XUDxFlaFF++G3TFkB+1lLGzaqaSk
nbqukzefqiYtUXGt+jTRikuejUA5LYOH5GUfuqMSC+U7gZQfE1XK8ffSGupJpvIzffDOcyKBk/6F
JGLQ/jwM8MlM1fH4YgwEgeS0KIAZgaxb8Gw2P/sxqBAqtRlyk11iKd4OuzOHE50NlzBhMBUCLFhk
gYhuzDEBrj5yAD/+COuT6FudgYa4Evg4Em4cpZK16a4YaVWQJR+MSUzKXiqvrdkHc89qoENn3QGN
5Y66JCBrIInUYjNhWa5CX8mvlwd91JJYUrITdpOYya7dOHeW2Knzq8f0/3NJlZmHRKsv4G67A5eP
NX4n4zjDy0p+qUb4voSGeVsPXjGiocjgV6zPFEet3j9dli+3Kg3vmaKvbWiP/abRS3AfOBaD7dVj
JVvEnoGx9RwgImCNEl8LynSP0+wPyXYPc8tTVjZKQINsnEl/OjrvH+3TiHxjzF+8FZkDFyqzsaWW
lf3BVpQ0Iie2I0Um2g02LtXAbRBbjFolVGjRFHw7Jbu2vpTpmn6FOo5wl1GQeNvj1F+0fQoHyt1a
h0hl5WLpEPmhzZpSfn0FQbd8YqIQsR066Oyn4Yc7G9v2hJytTYQPC27Nxp1KjDq+Q9RIT6EErrmM
cUVccoGIQaVDmna0wgvFjy9zZ2hy3eAUGR8WUWuDpfMQG5WL/gNLAV1PBFdScKjC1FXzzkPKgte6
D0bWbihA9gJGGZQpQ1YS9zV6X1gAV0rIT9wZaXL7TNIP5lrd+UzM7RTeGcu8SeY/Uyb0jXIoWCeN
qDjME/XjHE787NEFDyG7twaheBmXFyyRSNDk8gUS06J4kAwxZ9GcnIquhqouHYBSM7FdQc99WNgX
hkWPyv6mLPZxg6F9W+L4Wy0lM13dkO+Hyl3taJ1AgyoSsUZu0YXE0vl2ZkaAAnZlSbq2X3/GXVqf
t60mGpcHk09OqdhPWq5v4xliQ4l9o1QgRvrBAjDyPbOqP657twtT2eeHG2I6IwiBtwN0gpEFs9/M
+x5a9iVH9qvQazxVho2yXDvQujTpZiXMYjtiBNopUAypITdFNe0rnTaSyb+6YFS7P5BGAF7hMbyb
D5V+8wpRJJSoWxiZ4JlIYlE+ew6n77pB6kBV2kvPuATOZSxDsSvsWk7Vm8rETeqGgnn+dDeOqQ7T
/hSaS0ZrrZOLMZCCpp7kiPjyfv+Kr6iz/fvXYT2WcC3WXAw0aDOeD+3064UmqCfDbo1eQiYufy7a
gmtQKhknB7jkJTZkANJ7OiKThSfM3lFAyKWgdhZuiEc4gyjKc6+njgM0tKau7TwBGcmNyHfnpiST
QltoG8I/KEdlzoH4Q5tmxewH15gEYDrtpN2vH69RgNV3A11pC3YCegVccFczlz1VEAnvm306mj1S
YcmG78xdMAlfsGEmTPDjMFy1h4Dii/NA5zOeR3sN6dVRy5YQ/Fvkf3MUpQjX2iGVRU29o0Wk38MV
S7LiPNRNJLC2n5pdoIOkOClS2QVW1Q9mDKdEcE37jetnwpefs5Nw16Tt2IFq2FjjrHo7+43jLJ1E
mQ9ooNuEI2fuINv3g5aXWX0glvEDWO/KO36YPnlD3NC+RbM20p6HQwGZceyHBQVKo4ctd6HiqmDX
/hncNXXQ5aaz0AW5nneQWumerhZA8LvJ2rOwuBOMRuOAAss0UceZCBOTkIjYT7sIyzXenGW4ixIo
1YOiktEhdRahJ51s3528CksRedK7BSGnZf6h2sZku9XcdtucnC3yBRUA+9ZzeBbVpyGLUiiG4WZT
xFj1lhddgaQwnr6vqP/PghZ55OiuXfed4O5WnHDEwgbwVZJHVpnjBxjbLIUj6dvpjufzpebRkwsd
VyYiLQLT/d8q8K3Ps69Q8Wum+dBCGuoVzQMSToFtu4JAFw57eJHmF6fqhH71tKCzHQjoMAT+WuP/
mXMMmLXHGY95Vr4fg6EqBYa5cxkTJ5eKbZC16nhOCrSO1M4b6azUmYfF9JmtqXkPwjpBVpVaLZq2
wQAE524e3ClKYLwlkP/V4MnfEQuy7vC3KfOqhkIyzpBw84KqlinaSRiSsCbm7Ef95GaLxH7YlTMz
0s0dr73J6IkYRJz0E+f0mJaaPmeV6ZgCEqspZFdUD4E/ue/bhTCqBx/R+Z8Bglrb9l5t1Ne7gXzA
UMxfmLq+UEltUe9+ex0Y6vNIiEsI3aG9L1JOw+6ggJjGjqqETzym5KeO7x7yJehuz35L48usV4oB
HUHBZu6o7lRBN+/TCgTB8Zo3fw4HVMV83iUmUdTszxiR0awGZwH8+RhGa/bBZhnCQKmfbKBCXFIa
Tp1sVLVqTgu9pUStei7XQHnD8WwQoXCFBdXj28PH2l3Tihrg1owoU6PLdNtRh4fg5vuanWZcWP/Y
ZgscOKspH9zi0DZcvcIfDVACEiXiBldY1QdEkYY1OmFRUK+2Omo/kHmzYjbkJ/pZiNUUAPv3k+9q
ynPxrCRXtyfPH8TQckBcC1BCz0tri6qs6JYgvlmGruICB1LmQtAgQNq9JqHvwwUR3c1WVcQF6bbe
lVN+ikj5Y0H+gHpxpbTBQvOQ+/O3pN1gHX6bn9uNm6PQhIcSSv0Af6mcT0Fb7/xw5mHbWW+XzXCr
1VQZYRTlzfAPSTibGq3iG5mDxelaeAcJtnJh4ywFiLXT0vhYjcOVIqDkBVANzAEt/WGIrM77NI8p
j1kuLV4MTQFWNMxRnI61xpaZ0JIukpcYbG/7PnN7VO3PSPtUBeRtnfjt3QKIFJjKbW8uql4g/7cB
+i2SfGmmo8vmWjKgt3kwoWwcZjh455zKFzN0CQ6HGNT/8WlaErPR2hgVEvOXjJStgX/70gloOquc
0H2vSlbaHCQpIXoJcAsPzUPIh6X2RLYA7fZLZs7l3S0ZJpNlagTejT0QmlQ4JKOfhoF+DX16132T
e4lIOGFv8hdAGpTILCe81QmayhBMtIhxcPd75qrY5CmOPZHkBm1qU8GR+VcstnXzhRBKcdX9yfRL
NbwpJPKUs02hcNcbmam3n3BueV0vlCKa3SgwDc2TefVWJgonS5a6HTN9z7e7avGqu5WNt0IPql8z
WUIzX9rVV/tiFPt56+7GHOPV3SyOyKEeRLyacl4MLXBAKvVvk5wh+32aiNYjg4xQmOyPLbzdamk8
FG+uYvTMJkpyh3nrDXydqF///o37tkhGkKydm5ktIHrWkgttdA5wIPBR2SoG9b1EBYjR6Gio2XY9
uzud7Cvl9PD8RNWakqEwTbUL8YgIce4RGSfr8VKvP55h3avxn/O/raYOtyaySqYE/m2N435lCfaQ
pIv/la/WHjhsolXy4gc/v2vIw6utVqEKX4tBSW+Vr4V1YbBV9gu4KRq8covxDbOzmSWZzA/ep0vO
9VMdInFQgUY8+63EDpsvDyquvFZijxSlRT6v0MCGhhkZWF0paFl1snwdZ1FOmJie7rILiNYBIPHm
LZQ4nk9GpHUEuJisp8hjPPQKcK6vR+b8ABQqp0cg2lBjyb7U40z1vvRzWPxNkbhF3lXudd5cCqOz
eTrVhawJ9R+gbrFQQeOEZpEn4GvOPnAVov3O8MLLFraTSRk59JR23sb5r5gFqkzS6AaSUIiyZ/cA
wzYL5GQrlBsw/ECBSo/x9PRLiG7IBjnFM+2xZ6tQe4M8xNRa6FIGd3uKwsp8SSmfPyy8ODVTz704
hlnxuGeesEQ7zkK106hiQIXa8QDPSO/Gi8NfaBpvgn2WGWiHj6dzicyWndygNcNYi24kFhdws1mD
D8uaGDurWsJ9ScepIbpu17Xni9o/tVZNOWF4P3WDS6TanR5LCkV1k6iup26zSbnoLGce6ZpcNPu5
ksUNAXxlZ0nISORtmUVdu44HHGQdrPQW62iqJOdmOGA8P3L5uzPwi0o0ae4DdKVU6O7UYRmxzscM
3x/9zKcGn9VLIoEmRHNP3OJhXuo68xqsleIMo2DyHGL8+XhLEXjEqE8AiHp+jHIUEvYSettzH5eX
Z1ROAdlLpEKEh9djm7i5whRMvHjSoBHzZQVb8YhRKrBHfuLv5L/AopShRhCAXML0VHOqd9isDZw/
bGdUnK3SjaNV4c2DvvhFspLvnZNavbtXbdZUwHKUh10ugKrojq2qIFa3hXa4m8AgZAXCwtbzeXPG
nH3/wPc+FW80aBtGwJkyILeBTV/0+18g+EOpLt8yRNjxTJwr+wf0i3uLw0m0HGvgnAD5sB7Q3SBR
g/v/CQIxX4DLbeuKC8aqvUYYY1O4J6rezp5ghAPkF0XbDIrC+pHEPH7GawqwxaXhCKk6rFPiFKqH
Y29/PMC5W0ggYb23Qh6XN8nUpfnqDVhFhJldvFHv8qN0V1ZTJY+pbofqtq34Kf0fosqSucMhLCzW
Qzowonfh9bnKzpIt4qPCJnghfCtiOM5PmmWP0k8IWFnIhd/Jqss1u18ffSIdx/KpO3aTOyCzWq9Q
hp/ZFRWeL3dxNI0+3NhLPHlhPFAqMkPwEbg7uV0iIykyibjFHZXH30nvLXTbZDL5tgueoUFAtMeJ
DpJ+cA9jj72++6aj0dAb9o9V2yXx5VECnd/1VG9dD5nHjQNa4r8jyrQY7BBO12naY0JBviC/lRmw
BXyPR0trG/zsYKq9xyXPj417LXs0H7iQyvzYOyq5XJbCR5HjYKpYHwxil5l169Vb5LFy7VH+Q7/t
UQ2LiuVQHi9pnmctC4ANta9xCOp/iNSSY+8mdlaeC87dLNxsvMFVP8UpkTs7VY1d7CaPvLDG3oAv
x1+j64Voy2MY8ON+sKzy41tlRYsV+f9Ik2h2E137sWYGGhR5/wBPcrYrK2nYUzUSvjCX26NH2i30
/sqYgiARXub293rBrgGHFqdqvBjZov8CKsB7ZqaXtkjhem5CTVybYhWxxqCz+6mO3MkevKncYZW3
K1Uz2VLIMm9QJ89/COPeOH5eaQPk1zVJEa1cpTOBBfwHI/6M3dPqVphnEOIVuOdFD3lKjZxGBAuO
S1Ww3gifWOp4uVDPkuW53uriy+7j98+3/RA4q5FaKntMHOxr9CmaQPNx2XoSSW50nPkUNW/sxoL2
XS70ph3M/EhLAocshu/L2WbilGUD8RGjkfq8YL1iKvaO9gtSj4RcLVRh9p6DtMNtyidI/pIHOzRq
5qHBvnf+wnhrHZQEN/EQTdCKYF76/LnyIE1peI1fjGk54M2jAX7YvnsmzNEyAJ0ialauJM4GoQvG
f5Bv8sKQ/nWhHvFEpp/0/LOSqfF9zSLFUpc5t+hhefSbobnFHuFNNKvMSMQB3sjJW8e7HKk51NiA
IekGTS82MKeiRAv915PcZS/LB2rj5UboYu3nV3fZ/6OL5BjQ9dMEnQ6JwM/br6HPmMihcy8ek5MM
zJecUqgFUr777XRBfkTp/4Hk+7UsDbDqrY2CtzfAhyXzYF1fNXqq4WPhVCI449nsz2nuDWMdXr1T
Wkn/TK1t95x82Ol0AmbhnCfv2jc9IlVai8Jt705do/AwVkQquIrQQ4XIAwfpi+J4n3JkVZ9l4xRu
tx5zcUmmbaXaMtQa+aST2ykNkILYTzytxi39dWE8LgVyToghzOc2E0U7dMvRBVG9UYVL21b3rkAB
CYwpF5/cUbh48CYzw2folm2N+u1o9VKfP8Ip26XmWvg8SA4T/9cPZWVpUp7lxL+lklnqwROsp6gf
Lm1ggcV2PUvf3wHjl0WtmsMB3+JGtlqkLc+M1PWsL44SKkXjlJkOzH4upBan1XUPemQ99hmQ2eTS
Bq08WTepOZVLPF4I6tM1OTbnIMQg4mXYUS9cNgiskOyWRgr+65LRdth9iM9SW8Qf9CwfG+u4fHWD
ngfvl4p4NBI9y8AaL8RbwDp2TQwLkw9U+jiyT3s2qL5YvYSCQCphnVmrsyMaqzu8+eMFaJmR/aEc
q08odbhUWseQkHNj7dQd94TnCNjCExy5rhsC1RQsOMLxJCkSGBCFKAKkqvDPur8elAt44L6pKq9T
VwQcVpyPBVur0AZQevVzD+QtAO7bvnp3itd0SwGh506fQVI4Tn1DOKH+94KRmO/rRs06N5DV5+FF
TkEuhKvAQzaIvY8PjTHanzxcpEugBLYWNqll2SuPborQUiF8WuHWnQ/BQoxG2u2yiQ078+MmW9rw
pjvNFxz6nE90jRMhQp9D3z49LK99ldlCksyD4HGtqmg9oa+Qxd0vcEfg6kH8xmgc8Cc+/5JPmstc
pHTi7/7Ubc+UqWHJqTvODYQV85Iw3mGhRxyrEt6bgRmRGsdX6zjtctj/j/nwMd8aFwkf8DkxKFAK
6Cr0lTnTuQwSQGTNl/0ekV3P7dgJsrJH8kEhlxC+r9wFzyG/0+Yi1sJnYvcxy9lgyQzByccOhVmF
tjfh5VdPGGaG3dezyaqmImAxuehwvLXbfh7jpmTdAyA5CSeSH5BnialnClKmVyi1wHUOJaGzEP+2
HIM/HOGkgSfL2FD2z2w0nzNzMT6QxOv35D5OibUV9/Wd1cM1ECkW5f0BCB/lfTjAu7eaNpvYF2tX
Ln6UIfX9dQaH3ujQE61XTpw0EilqdFLTINlU2dQdECnyoBYYzzkzsqqvpUaS3XsMMWL5KSgeexrC
M07AzuFpq9ZhXXTpAajxjdoCsx4f0NRq3CFi9qqCD6dDlEAFm0BYwCGUvwuPqydfMItAlvcY646l
78rilCF3uiC5mOOHVzfl96JDgqhrIdtrwSDOwbFVXOEyhBrnhcETBlRucthZ5BlGjdippaVwRlsW
U/zGpzoAOQYN80vsW+KXsi9Nk+M/ah0t3/s0li+L3Srd4+k922RAvve1/4v/YjDTKheeNr+srzM3
eQps3WLxMQeX5z1L2lixoMHLcSoj4PWnyGl6qaDiNT7YvQVfZmYr11eeHJoDlq1I4bXJkFF62Byt
rsmMao4EBQeglDCP2G8i8r3W9h2lkDQ2QlKqcRb+FCM3fsxUKLKWqEcBPzuPHwxgYzSoakpjk96B
MDoh5eSYHiHRBY6ffoX9WKUuUHboFedNvHRm4RQDPFZMURoTpXuYdgXi82t8YFjepWFIOOz1w+TG
4Bc9sUUXx+r/e6fkgworhSXbQvJxc7t7cct/0PYmY8eZU2ZU80oriZUrKBpPSM2Claim77Fg9WGy
Vu2m3A40k/Q/ehbFM+A30Txpcu2CmWEBww1kZNGxS2qIAJy3aUdfHpJRM4fSjxywDGdzv4O1dH0s
KbcTTDbauJmbORGVD3WRGo+8ove1LoJqJ8/14fCDmmwOU7+up3N2Xl7NScDwSzyD6ItvfmMGwSog
0vJmzaj5yo6wOK3cXWeHDxudP3Uy2Ig5E1hTiNYiwnaQlgWxD3wTjX0TrGNR+/PgGnLeqN+72Hcu
79jvKvCHpuVIYFHXDVLWdNeRG0kGZn3cbXENydzT0wau3AGgl/syaTlUujgccQCEHD27AthTuLO8
r/HsswnMH3ITH97sgyDusRXRbYP5WEwN2XwmrOMZPKqqGADwZco4eWGNETouKzYnMBSIt2kACEqJ
qKo/OSo1zhhZ5V9RhXKnsd7RrGrhy7XVSyeslQVJlP2qdoX4sleD0l3ogLwCP1jhtb+maPR1lmsb
jJKdng2LfP+Urjz8gtq5FV3/k5uXpdXkV+SKIkX+9GZxJ8IgZGz7M/SbDSIymuNcWUmjW6RkK2QV
gpcovl9WngZLULUyBfGPUrZiKBUd84k4AGPkwZImDr5kLoo/UuDjX5jPyUJrGIfRH+G/y4DrU52J
ZfDYldtAPeRh4Mq+T/VG4uzbRoZdQeMJSnqqNR3gziLsS0UO1MluefBk41Ff61YzjLsjjNv1RVRV
WVDVux3PDcml29QLyYc3nMVc7wjhKcY+2oIdfY1wfKglKgmVvZHw35Ft+ch/psfdoGzRDKkNsrgP
couK8mu5IpvvtZ687uJKggB3r0DKCBnDUNI+krFIVWRZvhXJdTU0i5aw7KgerX+cSWhWkmJtcL0p
VKC3oJpRTx6z4S2/Kxkuu4UdhhhEhxoKjaQebxvVKac6FiZwtMOwxDDhmVXy9pQ516m61B097mxZ
WBEg/eoDiMp0PR9d7LP+s21xxYJOQxwUA7cBiu3+Nucjbn5uNHNgbxFpIqXe1WkaCbLhuyI+pbKo
UwNOT2T3JHUrNEJuDZQiOn7miaHtzP0eVwl6dR8KHeO1Hcd2KRnYwA4r82UN/qB+oqjfg8Y3Nmrv
pGUX7I3H0sH80PldUiQUdUGoEtvpCyCLm0eSTnSkiMDgtXYrThCWrRJmGwukK1J7VqzFpl7TxCFG
wsOJFmGfkqEllx3tiL4YychA+ujDVTp3zF+qoLdmYMbYvI/87yhXn/N2dRt8u4AFGMPLnVkOzm08
dgSA/l0Kv5JDas0TJ1iIY9mayE7rHEQDo6uwc3UHd7np6wK1b7dFACKVhDnxfcY+K0brViysbot7
3BlIHD2h5vcAOSn8Brzgv+/AmAeCKzNJZ8WbAwkP1OKaRLvBpPnKvN+60LZUzQSh1jXyVxYbvfs8
oHFxtB8ynWlzc8NCesYBAWZOPMVLqM2+1YcsyQdp+9YG723i9ZbdGOMuiJ3GJHoyV7tcXAYp6/IB
MFA9aXXKUFnve4QXWnvLgU2qIaQfUhhclSNknUDWWUedXOOkLnYZ8NmxvFsCMOmJMffOmrv+ew1/
1IyofViXQintHZphFQ/r3qrg7OfsNztc3d/Vcn7ck9RPBpQQkMQEp8ySoE3waLp6mc6Oy908iTPl
5sPI4Psq4UqjpfcttFwjj0UPvxOXlLVvQUXKU3iobIIS3jaO562/9xHBnej9m6L4clRjOVJ/nMWP
TkncgEiAVFa2lBqt+KqvgLU5tyFvYRt1hL5Feit/mC84DXQXYoaVO/iLQdoDj3Aij0yUfpn8LP8d
Qub5Ucy/lWT3sJssTx4k9/QYJsaCJTx6SbZFDPyqCA/tEzC2ThNVt+BsGaEqc5sYk5bDr3fYNXN6
X+6xzPs06jNua5wTwXuXaV7Sw23UsacRySW2Kg96yxJFVjZdD0UvvUFZOyHjAlSSGz/rQ9SFfJyT
vVL3bcuEzE9huIbiJ8VqPawXjIVkwbZU1IHYxdR+Gnyxh/LJ1wTk5LzUlluIVhfvilE1hz6hXo94
eEOz8L6niAi31O9G9K1Vxwsw7oAoC7FduOvjUL3EdDmi6b0NIbZY0M14Stz6PxeU3ikb87jkb4ig
cljsNuwtynlZqBCgMbbb1NIchKy1dSlXmyHZ+sj0gNteiQwQF8g1LRf0XUkhRp9wdExqL27btykp
lbfa7pk5EFKQDKFQArO6QB/o7/709MTlifePX89e/UNKzxRIhsSpkj8R1aSwdMUydIyQGtFOM0Ya
kU4pTGw9723VJBbYY5GhnkpNpz0tFKywqO7ZUdcP8B2Wu1TJF+jhlwgx6yvh/XofdchckwSmWB22
QEOk56YxYmGzm/rjkD8ucT2+xtaPeVLOu3iKPfboHe+41gYmF5ct0b509eXkjZgM6iUE4HvlaPOh
YZjzAWRgfEyFtQdAvr/UEQ1V8xPS2mphf3oCwtMfQ/aSyK0IKKUzmsZWGa6Qx7BCx6ECfdXEZUvz
N40MbP5N+ON0fe/4YX/m7RFGP7a3HycELdYDecNcDGtyOMcZJ6LJhYBThYdwNnmLCl+zVpMP8CED
4RRBRsNsWr+IwzDUfoYEWb3Fbj2WAzt4+4STpI8gHMFR+5sA2n/eHFy4PKIK1u5jBLakccci8Azf
J2Y2KcLa6sA3wHWsPXFxMdvp6+Ib6mdJ3nkqb1Y/W930qaVoBNZiuq44UG10ShXDaLAWyhbCnHvE
H9hxXEY8r5rvShY1Gy8S7hXC0LYdx3bp4WuoO61F7ZziUIRFSJxdQq74td8qlNWdLJEfZehEWoum
fSmf4iq3x4ShFdxJY9bOeWV/BxGejtmXjRaBSN9IE+YFs56nPXJZjUd+aoMxUq7OA//IduuK6TCT
MwhMW0HdwpaxEZthJm0W7avmL4P1rgiJgHQZnTJ/GoDS/B4WE8bPYBykTYCDNaDGuLjvrV9EX4JT
jsLKSqERrCPWsq2LIFD2JftCv6WtOQIwnLD5JJrB3FcKQqTQoApn1ahlfJ+Kaqm3CygZxY7vM/kZ
O5anUgk8o5WyXx6WYWRle6czdUBO1lG0teaWuvix1oDP05Qkb914OnVqStPgWcQ6jfKoF+dU0vPP
/QYidvVaI6VRooqE1aRiZPvXDRQNkqVzMlDXpE1IJbEl9pgidK8w3j+WIUKQjhZo7isn77YNYB9M
YoazXYb3iNNdrGr5l47ZFgiIKLoWULbG+GkDmxGV2Igh5Nnao3nf8jb/1EtgXfoLcy2HPPGWOpDb
hti+II2fJUwvPxeHDH0Sy05jwSSEfIX3KbIsbedan6vW3bDnYzbpwfrTCYUy2nHXvNNHzCNApicS
VAcwh3YG5Pp+730ohwpNxSBXY4E00U4WW9PwvQIbuskYmM46fzLDt3xNhi+X+hdxmKXe8RCFpWfm
9YFHsahiYl87vJHQXZUCSpDcIA/vt1YyuxUeKMpGbhvUwZJ1+aBh7IYySVTHgT6g+7Mwt68/WtnI
+Kz1zvxORJzwuckF4te83lDvbZ08eZAI32uXqhxJUFfSa+clOz/JAK+gbzsqbes45o+L4QZ5HiKD
b5Z4/EcpwJiNFswlOjelhU9uzyTPg4zBzUhrgx2JQE+rw/7Zf9Bl3BbSR95DUasZtQFbBKqlCeEF
BCYOf7GD4DXPCX/x9Va0IDEzBx2VB44YUCLcfQYKItiAXubVC8urIGNH06YPVQqKaNrG9xhxvFef
AqGwg2LW6/kG+Bh/RQ7248oQ1Wbd/OYU8T0gHRcw41tX2rN3HZnz3nuDk6APjOiv2Kc3RrBUARpY
34U7AQRfqqLlg6eCt3Pcq3UzG1iniTT8TyR2tTXOxaFcZu1A5CEayyi6bWnR0+gbnaFwFGxoT41X
D2QeS7tcGHo9YoZO7gg7W1MWZvHK4VfwwXnIDQ6n5+eV01cYDpCBIxFzepyO3ViVNDezbwb/pP4C
Gb0a0C2ZDp4AMh1cJvwGIwWZPXxTLX177WWe3z/75yreu5a5pQWyVZiZELsVyGOCHULyH89mD1h0
+s2Af+8hC0N4lG1noM3go6X5WL6FaC3Z6hv4pQ7EArdwxPGei7RCMzdfkicy5vXFnePQtGbncVeN
iCfLIcLKRI2la8fXnI2oZ6NCIagltm3R++m3IosdIwVe4pIvveNzlfusSO0xH46shVskrqghv/3n
DjJYwQM0WXsMY1AtrBeyeSnbBWHANnXcZNG/FP1V4I6N6fltRCUUc0sVVKFN1G19uxH5evU0egv7
oFO9+M44iKa1TUBTsOGXcLizqaEMeppozlEUVhQda9HdOyTOxtLNHpPggmlfcNXYN3157Fl5lVgi
DOYrq+zCDfQ1Gq+vPGipe22m0u/mhNSkMNC401+u063498KV3IW04mUAy6biCJE462hALEksmm6Y
AI4Mg7HJzfp/Rx2ZXDcxkbexcznawaaOmqsn61ibHziSDYtkAlxYHWLSMDhc5Qw6wuev/YgEww16
Bjo8BL7Vy5PRqPiHd9+Vmrh+febfh1g2gQRLMjmxZbryOt50sFblv98dBpB1L4pq04YbEsEr+Cej
OL+31re7M0rVKWw0bHSLuHXzchH06Ty+vGaALk2NKZDyIVLmspthpQbfUTBB1MzDOwWGWspjTHpa
BF+UexuA/IYxTr3ftFAX/QRnt5dNtyFOdWwYlB5xe4zAm2fxFTvnt1PQtV8WGQ0Ja7Rdk5/w81Qb
kMuCCW3Sh6Mnpgfuqkft8MdJFp02m9VURo+EnWZggC3uJ4WTkg8uMlLxbQi1EaEC0Cxwwnw6dLyJ
aHpdw0Xnmfvl5UwH5FBNnt/A92Fb36Px7yEf/OkEmCvmIB6wZ1vRe4p5ZqtS/AFsY5JMo9WrZEUy
pY3Oshxxc5aek5ZP0g8/Ra80VQgUgw/b1I2jXAbPv2lvLBs1FJEx69NFgOaRfIcv+m/ldsK1c4qF
JeGAweSavfyImQRX4G6IUFHkJ6xl/6MJDaMB7TnvKgHINDNmx6Um42bOHDDf6/bvZwyd5vPICupM
a6H0U8/Dsih/WwqOnbtXSXG4Dgui59qgkipLGqcxZDEbNdj+XqLOWpdreWDrLIMJIxacWCbRwHx1
QE7tj5lT8baUCYDt55lxU/jfmxsJRjTBFABaVWR0OTjqDGyOBowfKA4dgRZlWI+Ws5AYz56GqjWX
8pxjcYQ3iGN8K2rLfdP8ZJWBkLrxYGA8JJ3YGdJzTjl/aegJuKV0QlHFkYiL+gb5JdotPYA8BRiO
rX2ENyK/dv5vxIeFESuMssVUSYAVVhIqGcZU+9gI0O72bB163h9lZ8mxrIXKFujHHj0vwI70zbyj
JZgTsltRgtWLHwLcT7G9AVDHzyROFy/9O4vXQ7ktNcIO2SRfshMTa7Q4ctmRHxD1wP1CijJC2Qbn
ZQIfOH+FFXxmQNS3m1W45grr0cwp1cv5oSJSLM8ejin+t63K95gSxNnP5Cuc7+MSTnDmTzp7MjoM
T3E39ubQ346/dvHsSnsgaUQ+mL1RsK7zMgl8eBSBLOYhKlPDiasFLb9vEjetRpEkOOhUr7kATSZM
ZHVBq6wamWfyaocNRciQLomfWaxkXtlXFRYvV++1IgjCLbopVC9JCuKeeiqM3nuXkYtFktefrJhX
YTi0yRuUAH4l7VZWNOMkFNB4g/9/zRJkKCMpX6h+D5zQac0FYaxrFKV9zqTYh5CxaVqKEx2NwpTc
hYgxGKZ9AZgsX+OFeSqZi4FawueqGOH4f8y5sE6BDw2F9s7n8fKzAW7+2UsuRHcL236EMDXFYHNF
B+vZ9B+ln+h4IU5SrbAfvuOdquZifoJ8h9pxe0yCJxUg/acGsxLqj5hpO9nHbOdCKBwJ+px/JDGJ
TWEUZzVO3l3pWexpziqbRw1TliXE8c6Uop+4/QVZsc7OdhLJpdMI36pbaNfwFogK7eg9yykp+/Ga
rzvCfpYSd5hZPHtb0czfmI72Fcrnl4gW7p5uz5QgV+1i3pIjOIFkYim7A/X/8BhMZI9vFuOJ9Usc
7m+8NZ+eE6in8EaGtqcNXc9VF4NA5CPgrq+hnpL1v/ka1qDUnqy+XrnxuuUvvEvWwK8AQP+JJvuM
tJFRi/Z9uLTs6aduE2t0G8XA2DO5TMPWP1tR1MYG2pEAbto/+Qp1e3dtM2uUphD0TtMgD0pysLX8
WvyqJe8BzrHw9t46XIMtLqvsuorob0IHA9NQIKTW+2yAoqMy7X2Cu4uMYhuD392RkmyIcEY1JVxb
Cpaq+TT+mQx6VABgUrtqHyaTN/BRjul6qfzq+2ZFErksUEjJx3M6p/SIJmmk8/8JF9W1Pm8Bwpm5
MhUL+s76J5+jCQ0LvGyoWiG868CRRm366r8OA7OtMukMcnqt1gF63e1pWspMuVCpMzDdx+0OSoM0
yZhg55vHD+qnesXRnudZbo7WK4A22I8wMzYn8s9S7R7GekM9raYuOnliqlqXq1Xwrke+wXggqCXH
C//lySpam0HRCjeLBVLCeOjurg+KhuR6lUJAHsk3Vmt43lHmOAkWagDPaYH/ufuA3NNVuslGCZ0J
f1+vpRuoVaae5u8duWipQ4DQFtOZ5V1zUuVC9zwsmSATq0+nhfNJOfa6Ssi/T6JTlz7ZN8CobK0w
Qn7VXTNhf5d0RyrN9HxikGOCbxJGVSt0/R4hjeSt1LAeTgpnQhPMcsD2WcNJmaRba4rQV9zVe4Pz
d/A3Z7QnngM4h8t3H/5tvejLekI7FN1YDQAwQWAdL8a9jIJZ9R4Z0hEhxFJuFd0V6WN3gnODrL8T
Z32NGY/ResZyPxYWay5SNg8DQwRbXc3VEVthWspYmE6VwZ/VYnAeLwUelQM3hUcpx5cK7MqaP4PT
hqo2bwVAaijpEwq8UQDvGYWDsF14HXYQLJRNpuWjwRBLKhnnBfFDmsbSxd2clug5wOq+WpwUaoZw
U15fOJgJoB1V+PX/YX7gqdoVqKDFB8NyiT67KoItnKvak6LZSb0ufaGfsk6EOVgQtAV06uOwAdpt
lsncKAJ/PYD+eflyZEbbvMsm+k4fsiZF7dMb6MRWKkTfH5XtIGs6H7VVqbJiPnthSfu93d2pHV5H
a5sbpyBOkYwG2V0GpE22QJ5S7JWXb+3W1W0Jjl84eJ0N8aSMMxmd+Uk002R8IGu6t8c3ORSviNAs
jnpWAUZRLyd/mPC3dISdSmXnqSKDagLkq91yEApva2ufwpuCStbdeSWbkmerBnCzaMBX9pNC5xAW
OrMciFtk+ZWwINURigk417szgwPbzZQixAD/QLB0YrFHHx5ZW0nSK28Nam1koNMxToi64d0zzIxC
DYzORSIYFGBPypArE6dwc3mswwnLzRv1Ox5LOriPgRkLLF9nsErJ7Czwm9Yr78ZhVJyPA82Tfj3L
L2nG6D+LR8xul1Nxv8N6BbtcgYAkAsm1NWGG+vIMTZwMP463NWzSMPzX8jOggJhl+vFEF1pUrQ9c
/at33x9gsfxJPQOW4VceczhMjc38eR5nUStVBER1vSL+lq1yHBomCCp8fZ+3AjxXsjuX9QE3VQj6
BqPPY5vYk6IcEDKkSIQGDyYfs6Qvpn90QXYYez3jkf2EQ/gICfchumk8FhWMA07Wrt6sCsGNR+i+
5B1TdwR+Y8XNSvd4FBXISv6M14xEpKa0R1Ve4kuxm9xegOm075NRR/xN97MRFF8syeyBQZP6CDKM
tG+kc1TmSji6ygWUcXMovz9Q48RggmezSqB8D4moXim5WnT2LuCK37/T2C+insz9gOg2m8hT9F7O
CiM9Tv80T+56vSqfoDBrvBFtAWOgMmvYZcMOgqNmenR57tS1sCT9AnV+973etqTyNxVMctqQOvU0
t4Bw5uM4k6EXHF5+nbz3ad70vDxLw/w5B4OSW53UXlIdOoNvpX+OkNMUjJkceehgF5qD0pRyIxCU
7vP+clnxHE5adcd7S3CpbwiJd5+8RY1Iuw+3sPjND95QF0rs4Ii6+nckQNKPYLey0nvKIGSPY7/L
6oXuS11C+YX0ehFj+mr4O4BdVeyHnhilSxq40ObUh/1uoV/HWcg1yBLp6NAAQ4P5y4OpyKm2KvgP
eMkg7LXH5F/EJLS3w+FjMujM75dYfKW6RJLfakjyVCuZcLz70IpUq+acE81gDaNXCmXmalxO1Xta
JyYPQFmNhzZ7k4/rMa12J41kaBppXGFbGpbDlbadOIcKSzDtD1ceMN4XmuwyzqYwPyGnL9O8mzag
sGghzKzTyBcfvkpAjeBQJGHNhz4JVqeMGvk4HD6+Gokg6ca43ZjE9osGr3Ssq2IjrAhLeGcfxzjp
iVlZgvzOqmvEf6FXhZgPPByyim2W+BV8Ixb37ni5VVpLRtXbJpOkUcMTHdkl21h8FumNlO+Uyelk
EtUmv1D5EwnG4T7WtHfc7scYe0uAicyIZU4B4o9vhgYvOYU8AZaB2p/Qv6cthXnQi7IhbUilwh2+
zmVj9KVm+SF8xFW5ALpHiBNFeshVtv/e/IxwJ01EywUWTHM0EePoa46mc+aukSIof7UfwoHT5LX9
rM/E5iokHe+KBILmv4rmspSdQ2ngRuIY65dT/pUvzXpsPeNCdIS6R3j5yms/U1dxtZxkdnT1W5W8
RfYCTwp3schnNb0HFPteCv7L4u/PEPaESNd4h1XQYYefI3CTdknyNhiyyIACCtAbovdsD43Jfv5V
LpJQjxeEaTJi4LU3YozkMBLGWbxwSqVk5rkU9HMRhdR2N6x52CHfEPoChEtOW+RTr2XbuKw9o9NU
Kb+ukFMcvLf6757xusvkGv8twlNMctdBKClsym/tfe4qwz5hOanUdmsylJszNNLeYA1wd0RcKpr4
OkL3EStiLNKz2Vjk+WNf3ODx+Kmu+gcPy1PjQwADBt2vNKtMm5so2xd6bmhoexyC7sq3cFILRvP8
rPtaSj0n74h9W+NbFeVAN17tN6QKTiTHHyjk2En8R2iCzC3hALzbemeEGBABX/PTvC2Ym1EDszem
Cpx80Br3NmPAcXqV5tpJMny8kcZuRpe4kCETx4DOobiw4d7DCtWqIeMEXNl6/EB8Jl7EZHW+1M4Q
eHsEv8ejpw9nbm9y+9yRjOwDhXlro1Y1jLoS1ZKiVLL0Dd7Qt6WkGJvRBwj3rlqaimlPsEmZLABj
oEw7G0/+8S1SY/zebG3ZmU7r8gY+9iPMOQ/faCAoT2UefhlJOR7idM6Vw6+CMDqIS5+cocYofGSb
TWIymaDVaQ1jlxAQ663ty7hRUvd+3j3ZeNjQz+yfLhOAOBOMHx/rrkhbF2qZ+4O4wm0DHcXwOzl1
g/O086YvHgPWPY+G6U0V1CSGbagvI/albX3xAZoZ6vj/wfmKPirqp3oP49K+RQTC2T5qDyz/L1nO
c5x9+6IpTzpTktAuNjdcoxcV9wGB9p15yiZu999hAbTpFLAxW75K4qOG6JhsQdt0ceRspabqS/eB
riMvTs1CbTKm8xqVlOZ5ETPPSjlDbnLJbeVD2nrWX3Yizi6zZWnCtvZ7+adgueEjs93+C7tXHS5b
x0EOVGwRml/skTBMdYBQIQI1WFLuvJzuNK120q4MwnxHKJZJmRiehsc5GsyfUUFlOYbZjc57bdZ7
udxFuisWNMhBiEwy6pQ0NTGfHPc797qMxYiL+zXJTiK4NESukSHuP0QCLbJGRPw2FA4EU7VzxBJB
tQTs6G4WwS3PGFEz1ETHunoaMlng3HSMGFEjTfVaZjDR0t0sMqLKWGxgU9cmDmbtA4tZLs3OSpvR
9sZ5ezXWzC/Hzxern2xv3pz24y8EJiaV7KGC0ox4UmxtLgqXiTt5N3/WZqKwXafYbRI8gRE+s78d
Z5JvTJw8COLMrqDswJryJnWMthFBtWprXX3Vi7XZaPynK281HjkEbsyuG7Y13riyNk6M/C7eQFfe
gVoMtYBW8U7Y+k5dwsZNO/jQK76W1T24GaX8OAHmJ8i/Qtav6XKwXpMP/dIUn/+00IWcP4GGgJC9
MKFZ8+cqJoNm8esmjTLeouxvkydCGnm2dyT7FjsaIZ6V2Cr9+6SsynZmdWNBaHnXi7hAx/4Ty2q7
S4etfkN5qztGR027bTr/OXVDYjdZL4/+ODBW5O8NMKScIAKcd76CHkFbLTNns3uLEBPldwPvUAB6
42pcaUgEhFTL3w1aQj6SLd71aXbZ9jMeMHETaZMSndmmKMLAcmHwqh/Z1zjsjC2tmnUqDJWfOrob
d2XEz7rNG29HV9k1/WygIqfJ81+PEQ2Q1sepPqrYWHVPBf5IR6FkGqbHcrM1hqioYu974wtrZRZK
ryJpUNJ8xb5w8P8X6h3IuASUeYViJoQV1Ddu+cNxsgRw7MWxWjrzXGA1uVvziuUpEMKSFokH8oD9
MjgFqa+s2+9ZgZu4xLp1SUm0urFI+pQXU6n/ttmFUcBZyZl/GAUHCySblCw6Bv3bCx3qavLxhfOm
+iFOVcsgrPGYBqdiOYim/H1olowp1+u2KPZRVnOJWPbui1Rn1/xBm3Mmnaeuil3nojfazSbrlCdd
Q2hbxcML+ONlDcE93KGPm6ceiNAUM3oNLw/jzsKv7qa83uxERBlvQRBY4su16PIeVULQ8VAdDcFu
sWTf+0clP5lNN+UNkf8KmBA/M4Vbqzvmdcm4bSeeUXDefWxVJTwiZ8EJBl7zJ4CPhNKvoDJfeJC6
0vgnZUfmlggvqA26QD3RDCzXu7xt6WEdNwFt+9EDvCbskGStpKfcPbyKzOfskjlKVail6jlbyLW8
Fj/PMMNENmYi6T8ReeWbZ8RzXfwgHvCkoZXO1dCWFslJezQ5PJy0pSj01BsrddGWMLCGMrsHaD97
6Uih6GvFIxp6w+Qy4qM25U023QU2QZgqLCHk0/eYqaWxntioaVhtlAHl+jorVhwhehwgywrJFjwi
Z1Hf0nvDUMasB7Taj5jDGQ7VWzypJN7xpEy/1rAcPe1qvXKu370dIntuwYsG4eKkKZJnV6HJuBVN
XoxJKfFXByOQTMtiPu4PE8J6cuzinJMIlDCyuGq+oqRjCyLvpOhxNnGiVyE7udCMiFlCFzq4wEO+
unl7CVEL/ZLSHhtlPIxGilibevKHPyh1fcCALScvHg8VedebDr6XA5c5ZTBw6YWAfyoeY4k7dVmz
g1R2DZw90m0nDSshRftDE2gI02TQKpg0InRzw9YmJttKDqeLNS9VIkg/v1sSaSLUZCy0L9NMT7Nk
OyDuhtlQ2YH/T9Y20if9EJn41c6iAKRc2bbiW2FJbLp7llMU7flv+K9eJ7cNPck+lH+GpqUm27Bs
dsHbvmhIo+of4MTo2RO3en0nhcknH73nJL07Iql2DNb5U0V+fea1u98NQqkguW5CqgVyNCL4O3n2
PzDso48gH3FEl/F9hZ32xskP+bsrIV+p+cw2RmDYY4Uan9MtVQJL8AtN8jOOGQMJmlBOSXgYsi3t
eM33vxzWo6yQ0JxOzlcubIg4Y0cezAYDQd0HMQ334NcCxERoV2I8lYHwpf3Uax2jZglzpQsfrMJt
lrWdkRRYMNTNyFJ5GfvLfZLv/frQDBHhIywOPZSaM8sFVf1Cym3JVCUCDT0AKnvCUZz+NjEcmUkP
RwOdyRyXVI1rFQOqXRt7/9jhtErCrGgRETx2A0mQN00Q7vMpF3C1S2JJX0RQt/hMVyQZBW+XlhdA
tw5OuQaVpDdKS0ouBmX/PfXOTZyymdbWL6A3KUiCva+7SrV7Sw6Z2yjdPaigKkidXjKY1sP4fc7k
i8EjhH5pO1tScTtqQAGp819RMZALhQpDi5uP6UXR306uPZKf51ngbKlECbmmOIkFIVQUQV/GAcFI
IH24OQuQQ9ZcuuuNZMaZBBhBD4XfsSUrKvuITN3SkrmPEphd13kBlR4AmTIsWAjxPX5No1m3QPgb
LCfTlB+Gw1k6jCrSwoL5w+cIwCPIbwf83jzUAL7K1kbAOF1tlz95S7ExIuwtGuSmZHk0cm2Of2tx
HfHLLmSUTZFMhaK3pFQFh4M+wDx9emckLPhSMNSoWr2eoQo4Qyn2G713R30WeQD20xrAUrUSCl1Q
gQs3SiHQWg05i81hJawc3zNy6gtbrb9rHfA5tCP+En+5bTi3lGdY5ysXS8hHKgn72ncrmOCTEw2C
106LnoYGGNpWwcVPahRWE9xxJLV+G3oArNThRgvuv4xt+hUQlJqLIMqyUK0CXr9b6PcDsCitoSYD
i/quWCwaO8wLaRZaS2tvUg7kw8movZ6X+TLseQrjlKRJEv2GQZ0PKJmMSjtWvns0j0D3bs67XcyC
O7pWTPt/e+0xdHr7dorYgdotu7GRA9HAZUHeEhiNovAU6U9sVAS7FcXhV0k7eYnvqQl47sdICnAL
hBGcayiJnt37O9F7CKkwASv7+smNKkDIzeGRD2K5bSE1FrRlPXOnn6B3HOkhJjw8vebs9Fh7qXr+
hvUU0lAPh6AzlcbkG3f0uezXjcZnsYUkuVHd4LUPECjHxai5NwDufMqkC4/bmupKVDy0suFj+2eF
ZFNUI/QO28LQyMGHBUWRJriICWNqoI0wAvYjBWmYfFlxrKsfN7o8UYoOP64zu8LE0+1pvhHJsmXs
1dxISs+NE+g3WtKg7fb738sP1a7YVUskTJ9lTAT1/aPS8Rpb1hOxrlU7ZE+lJ0WzlBB+gQkOUf3t
aHf1GYvCaD1ildGZvycojOGcKj4q0BUfYBMU3w+JpKfWpEE3Nnf5wGyuBCkrvecS4LcmZNf1L9M7
Hd4gZ9KQqLSfnfWFPRctYhJZtt8pn6CEQ8MrZe0Qjn0nfOikd4+pxQreiI5u3uXriYM8o7C0M4jA
IMq5tLL366qiWqVcq2SzIVN6qEx41VdgnyNDjrIVt6xlwT6uxh1UaM1+A4QTcq5jeHjCWS5bP0NS
3svJj3hgfyVI3aj7u/TnvoAwpd0/4N2vs4LYaKSWHGNsNVHBGHoTM4DQ/MYzXOTtITPp1OLuO6jt
TDTL4SkG4BxdEhLtdBUu97t/5QEVBoxREgltCJu830CikPbX40yd48G7oAuJgkHdTBu/LTilWQ9J
Q/2avLFOjJ8Iuae+bgoSSSIQNABmirl7QWkq14F/yNKFlpxHI6fGiF6JfLPDuqb9+7mjQ3AFf61r
7J5FM8ewUlptM2e+TN530XK7fszu6drfEQ2fVdyrTluRc2vMv+3G/p5HcWA3ec/Da6gegWsLLhe4
up3yDBgqWZT+g8QamVz4c18e5P1KfcfCnD34qRYlknYLEinQXYT2ZzqynlQGTQjvsjq0VsYB/tBu
kOAaJXh7wpfGzKajTb3AL1snJ33RXAbBJ8+SKdAHPz8JtxIareCsitVGWAco8d3aH4cb9/E9u6dj
2qkjG51q+k1kN+MVNj+lrTVthhae0FIckP6WdGTKBzAiRXbdQO6BuX+axb+B43sSb48EA9c3GlGy
kNt6UT4jCjucKivD0VF0ta/ZDvlaixvui/H1hL5FISH6soxtWnSpFiAXi8RnaXO9CR/RRXEoEn8R
ryWBQjOCzhs1DEJZZxqtoETOOCKPjF5TWoimF5TjngAef2VkDIrtcXI0z/T5nhDKDORtR74cPdQ+
cLIdtxlAVBCKlwPVT9UMgSQolLgzRa0etsizchJSN5o6ydWBHFksGxzfmhrzSHmZzE3BSQzgAE0y
hq5Rf3k9MCH41uT96ZI0bSnN1MuR9vwkZuubCUFOsUWKfdObqpnyAz9dO1j2BubCvfMf/c0DGDWX
/mZat4PRuwspPBnxz8CnJzfSEcl/alt+oABqxPEKT7ly5ZwfKYQVrF14nnuyzTyjU3YO9RAi8cCB
+si2iBOM8cgexpIdmfgIw6MY9bWu8PNcz/8VjfGarYzb7NrA03HrWZzLLDCkJ1hTnmCejlwcgFnY
uSPQE2uswIY6Jt1CMzSZte7/OHykyNlBsJodQ32GoBsbBxwwDo5wBHS3MEFofBhokqsB0m4O7oXO
7vlyPciGe2BtipgwA0GsOZCkmZdlcyf84R9ekaozUKw6ZQc+8E+6aNpGNVWMIZnJEOvpN1EFLyUz
aZel4pfnsF4ysH+4xJe6yJeebaIandirbgxZp6DtxkXsT2h92XHc8uJUkSH1FhOs9qZhWHFod7C4
E4nvzk762BqyJ4vpjuVYOuk4axE0YiL7wpc4EaEuIVWtwQz28uXJbVkX9ZPibVfuboJ0MJozVfdK
tsukvcl2UzpNVmLYUpoHsK1WyZDydnK+Mz5DrsyL4oj0sqUbBjDf87GqLpbbDdl5Igdwf8Q5kFci
lEiztY0ZXsIkRg9MgdyYNtp+JcImKXqHF7LqMyh9URxxc+OfheGkp+BXeGVUH1bgqfT9zy3q0upr
3eMGkX/IxCRhi8l9L3ac4Z0MWQNV7LWkQ4s1Y2I0oY16QhWA4zVLcyyyn5SXJX0RC2G1qUBumfvc
zFMqf8mcS3we+ggSuAv4vwgNS6tdtl6LDgXQQYDT2xFa2XnKMdc3/ehZvBvyZHBaAhLstZrq7gSA
EpD/bbejfqQDd5sodMZTjgJwajz6grTPIpBi6XGe8eCu1Y/0Lh3CnraSLqwyaLbr9QfN3ePgrIKC
xwulLtIY5kNjZos2TSUpfHwWaVq6F2+xAh/K6IsNR1X+Fc+mpCZDpgiLfSKgDIio/qxVencV8lrZ
EpkNo1/non94PSCesLumKi7HGpfYTjkVu63UMnNkCiUvoeGvCVYPgFe2kbErzodc1sxl+X+zVPaT
RgTQazRn+tcYwYRKUwvK65NBJVbfK6rD2BBUboR9BivfFWdlWn4OHf1VrlMMfuVIEJIrG+hbte+b
jqnmS7147gJVccLs6rHSaHNDvyjhpWnDVQkhM9wYxw19nkELeJOF0bjbUn8g3woBzkZy3E3pgq4b
GTp0B3DMMNX00x3C5HejSmtMg7CdbEUPYWETS54/92Bj945FqbWau80pRh9ffR9eDCkta2mt3nOz
//R0IiEspfBiLMTYAiZr9dN+8qihmsNrJkTv+HfOxFKpFyCpbXvpcv+LJ9M0lcHTrrEQ0sPxl4n8
UmR8XWAfZl2WihdQRzVnK+rp3VKt58wjaS3DXMH2EX0ZO/BMCyHZAObXWEyGF314zf5QmS2ePxIN
+a2z/W58L6lAUNcqznQ98t4lot0xjkx6XNyAElsQB0mo2GPBOFdm/dfgnDU7QG+qq2+UYldNOoRp
xBdFtH5kg6LkEEXwaGyq3IiI9XB4xW8nCc6KoxcWYpJXh1DuU9wNq3s7eySbp1aXJAEm4Slzj8kI
1LSJ/iOMmi+nx1Q3s3Nfl6yRqfMhHXc7vnD2Is3rSq3fqtHl7GWOoPQg1jCplOkJY0RjF5ndhh45
9XmxlBC8bVQ61KFEVQ94JrIhlxqR6qNChePVUJFqxnz746RQbwjBOON2mE5Es0RRVyXFjzDb6/ui
12ZdEtYzzBPnqPA2idq4DjoO+SSTux93X4AaHWDfwmsiBfALxTps0joP864vdHaGp/j/FMAnpr6h
GxH3nP4wS1p5NyCJE9plJrPUedSCtMpJ84NOP5rObkdEKFC6DDHsblWzAJ4WEW5LFfdiLLyhvubo
ElFORP0JIYTytib2+SusNtoerg7j5MCl+8a494Qy88vmvEz0SfS+VLLlnVrqHQ/RpdmgH19dTVV0
zrJe1A9zoa/u6qAa288Ffb4D7Ed/pWLRO/AIOz/oOYv3tD7cMHrrl4tq3AQVdB9U76Ux29kOXQ3p
EhEmQlb46RrIQPcmCxTIbBogrpal5FRzNEflZ7LYMOzswRjayBLPD/b0UzMQL/ABkg6V/xD9gkp/
CuR7dXtl2md7RUHe6/Y5yCEQT1jF2lhBcxcrcaHRtj2LhbEtzYbULn4tKUC860F+xLkXNg/y49es
pCSLWpqKyNOHTSLl6gfJsSV0FwduiDNwU1Enxw+mP3JW7tQBcgb1w8/5v2l1cxZNNwjoOkr8eXGz
5lt1BJCVFoErxtMUd05CU0apsv9wfepEUXQ9EpxFr8TIKu/QM04nhknXg5ILDkXlcEXTZrDWz2m0
M7aNCJfb7RQl6lbhn5fn+sMufG4ziLlHfermrpcOJzuSgoU+bErdvDB8xfwpKfJnICLkeAaC1+uy
Xh8BwKqu/b+4QOrXzuJX8fWxYU0R00t/eyIG0YtQYwKPC+pelUySkTAvva28ZhUw1dWO83T6eI4e
vqTS7ik+IdgwqPwMRSjAp8QloXET+YVeZxKloLNW+mF8Wu5saX39l7z3LkziHJeFNGRK+Dn/IOw4
avgy/StKs+V23empOQD3ZRs3Nlm1IyTI6kzr5bDscTnuxao1qFukgthm3AnxwR8cgbG2l+i5Ld5o
uAi9/jVPX/O6ID6sM3Q7OZ4gu3CNrCAEMovlvn7DlEFJulbBzkEBYm/c9N6odkDzhqbT+306faEh
xrLnwG3L/7cJ3phIr3D3gUaHxAP4JmkAzil2rFYbnTft0pzlPG4fNBZQSbLL5yxpEBSh7OVOw/xo
B27gFVEPB/1tOBLUf7OHETUUQ1H2jtgB/w+YJ/7oaflD8QSqB/FJg5seHuTdvMnAMN68ii50Uu6h
hby5GqMKxuENBP/UIVKWWZeqGENQ07L6HktOvGsnNeUWL661JoJVUPD206Lx0BK3GMMDRyalskLo
BzSeE7cAYUEnetRa77cV83+Dv3CckfO7YsZQwqHE7ykfdEJA7s0CZHhZv19F2ckkQNUa1f+Uv2sT
rfrjIC8CHulMIghvnLjoTUY0NXekF+RCvueH828oOTSJ3G5lbvQl4KM0f/WRF46C+Jv9fF5e5Q8H
SJKRQWJGEDbTv6iQ3JyCXXWpVshBo/gvS/L/RLsipEYK5MFhf7nLKUwUujtAUTcGREVu+8CifbuE
CEIYjX25CqHSx6bZSMXoc4uZcy2BOYBL9jGlu3X33WdGl79FYZA+MgJohcgaFqfLw+Ex8r3uSHJW
LqoVhFztzhpNr4N0VQIringSeG7CI3shJI/BAIma0VTFdAHPM//tNz1/+/MUt/GhAEJuNQ9O4Dmb
vU+jT0Yp+s/le/tKAip2GRT7PGHJQYyvwx1MrZF2PtTR9f1edF/TjmGmn9yPGTrxI10Emm9sy9KC
hD0qjgKGuM1uh/8AeYQHdF7ZVnA1ZTxjLvE2FlDTKVrgrJ4q4qouXduhRIHO1I+YHlWaF03TrhD0
iMmKbSc6bPx0BATk81YsMJlegjA/DdVkTLmFgHyM3ZpKp32VHMSt1lPurg+xr/DJcaKKWr10RX8I
3c18zxXzWjXhGKpSFgXuUQaRIz998QKc3KI0BJWW0EqNBFWGdreGd2kwNbkrRtFl3yVmpIZian+R
oCqqRJ37KyLQn7Lt96xgLsbwyXyecVbDQYbmxLoDLFgewjwnjlNilgDUIWjjNc+uSutHM6gj697i
BBscUmNQuXc1oIIx0RMSXKYataujOQ7vAYJIdSuQRbRHDSNN0Jjwiwra8dpDSkT3x98T98O/Gof0
q70Az+5BRsnsU1sjBcqfa/obaY6Gk5kXw/w/augflw6f2BLr/+YhN6t3XhkDtV91Y6a/dZANElSa
mcqR6K5o3nGtXG09FwLZM7iqTR20f46xxp2SIPsL/Byii2IP8zbWjhm9SGubvCjjl7zQCUIJaKuR
rAjU1VtC1LjeAX+GQk839+x4SfRxOP3PVZvcwqJ+Zx7GPWirS9UUk00pBLSKgahFBSJ97VtxFo3g
Nw3Wu99F3wVNeEXMPm2QHg4JiNgxmLyRqdKQqxoTz/ISDNvMWXX9KnnQfW79C1YRRYCq1f1RCTJQ
6rADbbnPof1F+99oqUQJjQ2RiEQsMNPLlQ3TL7lmwlXRkSALcFWYL04Kc/kJvFxtAm2eQojrolaw
IR9yUCzmX/bToYtM6wlnY/Ik/3AWIMg5ZuNzeuIT+gqI7FaOEMQBXm8j6xR5KyABlgGA3U7is0B9
2aHdz5z9LEVqTVjA/4bKAcaggu89bf4eC+cQMRklt3F/bf7DpnrEBxqvd8zUVXJNv6aaYAEGhT3U
QTUMLSxOfajwv9pCd2k6Fs/eGyakd6+vi08atsXkIa3z97FF7x36c9eBpApOQoPV1hPxemmbxzB4
2p8edS5pLy+TWf/srkSHgsMvVS1/W+xlUUFjBLUL3qU0olKEFKiMULYqaQ7L9i4YNOs/O+2bIjzV
wzt/DyG+EdL7GvdaqnIw5td45hKJY/099i1L+Dw705p4d0ZR4wrR+7pF9Ge0+Kx3V8jkzthsThgK
XxQV9E4OGMCjWnZ9YunzoUEyscabNJLIS3jeKIZdoivIzXU13gWVFO+SKt6+v9WHdw3dGZexTQdx
7B+L5C8bIpZBDoXvp3N3U4YMu7Mcs4WTbPMB2MczYQRlDI0sVy922Xa+hdiHP9bp36tsuGF1svY0
VFuUKYXJv2uf8hD45xIhN8eSeEF+Szv2lU/XDQxlW5JJubhMwFpSFQz/pYKTWYcr8eZlGZVS5AFv
rA1voZkgNDC6LtCGTpk0gKA3oO46wQE7CUcRnDElZIM/wKQNJ7FwqlYF7ZK/AUbYg3VeJ31mgKeA
HtoFtg2WkDM8hN0AskeRbcj2GfWXVncZkUNdI+l1Cjy53NuXYXnXE+nbNiu7gba70CUm48bfJ+Tb
gjsfhHIaUgpXnbd9SLODD+bTkqhcjhPFOC5u5BD7QAWH5wnFmryRWGusiZOPnYKAjhKVLerNA+Ie
vl1dBG3gHwWM4ai1HpbRTYsQTLinDhBKa1xllCJrMPS/hseQBJxwp1bC3KAZYv7KDXDmgCRBqAvV
wchDvJKVBtWux/J6mtY2M0HmVdBmQHsiLrU9wCXvhLTXiMXzy1RFTBjG43Z1FUaamNjTmnarNutX
/bCcKcgAznJQacCQUloOxVUXnsOhemQRPQWrotlvMpkqxM+aacKN65awO+miDbGumtWMG8v2thY+
z6vPEMMSmoPF0J4CoB4uspEPnZxtS9vFAsY7cuIrIKu69baeyGTRw622LUWliZjrJYOc4DopJ/8u
sVBau0v0gL9itZBweKGrIIw5E1qDcMB2pTzKLcwMh3VoVnJxdIHbagsA1JDv0Zz5bBFYM67LtB7p
iC23beUQjc3+nL7WLIaT5ZNO6PIswQ2tieYTWp3dGTU597M+3WR2JQ1voZwZDKcXhqZ/QTEaiK27
Rfv70IomrQeyFR5AbFS8yVZMBNcXbaMcU8c9x2Dz0EBoEQaFafYoiRam4B2K8fH5vS0v983qbdZp
BYK84QG39JLcxGHxoVUaPoHqXvmQgZ9iuNf1FTTIKT3rjlJ/qYe8iCOAPai8Rm0cgWEY/8hx5Wzg
SY4phCeBPGjeKUuhbxD0uD63cXUDDxDyxL4B7VxvLw6qF0dnmGg7NHl7TNjk22rj/CA5kuSpJcY7
Us5lhYq+DHIzE+3NlOCg1NhQjX7RqMM2SyZD5s38pYM9GJrRR5h6znnTNeWhAHgrF8hviJakZxaU
2sLk6MN7nqbq4sLTMHJtk0kK9XBdq4EZNMaOnI342ZkQaoHJ6B/NvkFLS4QwvyvjVimUe6lMGLu5
RW43IQShmEjueeD0gIQ7RtBemlpKxnLuBErbTvo12uYCFUZmEXzy3VwZRHEENZhmW7lxMVV2eUyg
Hujo5GmXmaF6GfNb/8pL6G/LmmvPvaK6aBh7vePsyo9pVPXQfwDR4QFGdgr9/oMa3wp8r6F07w9c
VgGOUvK722dnqbZQGVx5O1RsXdD46ricIBoVrlztoLq5XzBo/8WarT2ZCNV2qMlnG4a0e5XBNFww
fKeVkT08IsSJbHCP0tzGAmsgs+3jCrZD0gDhHf9/KxbExRHR6epmzPkW5S7Ts8+oYa/PJv8v8wdi
bmOlqkvX6oaB6vLRlA1jvOWemavYdOwkE4xcKjJyA0Tknb8bFAyXWuiVD51ZVbgXVqQhQEGd8bEk
rD5A9Hi56m7qKdXACLyqpSWlsSTYswE2YqHaz/1KQxxk1svc2f7142bDa4Q5RMCqldac1Qbb9Xp/
nTeaNyIewXD9oR4WB9sLOnH4acl25pbw/jNGWBFXCYi1Je/L7Hn5HkCqsG4gdDSHbFaP+tx0bqa3
peVvDdpQ7bedAiEegeN28llGvuDt/lcJlXyQH+Irv3u/G6ScKe51F1aejSTF+Fa3ySB5YFEljpzu
8HzH0xlLRW1wJHsiHNUnIFiljVAPp8ZbjZlfgReOdp4XywtId2tP619yKKkRaA6cbK9UkZ0ecuQZ
pywrKPo98AYItKZjTP6OOoRTdNgZvllV6wOJ+yH8Qxcl0FlmQFIMTl9ImI2fcgpJcPvPiRKxVlO/
cZKvfsHWXbOyxGUwd7zkxN+WkwuWCrJ+9V63R7p/7Wp/3g6swjrKg9ZJqq9+/RqeW2h98QvcOehs
lX9KrifZEUM6gZycCcQSTwYCxXsauHXXAkjCV0kRJ0pnPD8HMPO7RJ0CDW2NBtaRQqHaesSITl4n
Sf0SfLFqpmuF7ZJVmAgiOI6r7c3UTuvjQNvG/J6NirkPArQId229Y0kUEhb8Hd1+PqM9o2XH0urM
MOAQOpNN6jjn64lhdZfzk9pTo9VBXhJDAb5O9xbNAlT+0qLc4NOTtM93t6pl+exQasOMAIidALud
ObIZbCHkR/EVtPtT06mo1CZyYnbTJscTTmS/l71n8/d4frW142dyrb3DhgkVO9+MSJbMwDDWYQvk
NWMOXxYxKsKKKVjoaoagufsCbNlcYAsD4Y5xLdm5xda4UOgzekTYYOC8Mws9sM61x8omCTHyk4LG
JExu+XvV0V+Q4zXievUacO54cZ9kTuZ0/7IX1MFywSOj35YFuujwQDCEUDhh8Fe1GLj9KbveNY1X
+FJK8sfcGXjRKpd5VZ2be8UMwRiI4012Mq3/aoLFBUixJqKnxiv3FUG1oUsCrbq2k57ZFRZmAVdO
3cX08gVxw9HjK21QIoIt7EShkrVZFXpO/JJvklUmFDiWcMnQBxeNOygvkjhtz3Ij/lMYraUofMrU
sUkmeD6VRbA3jwnpm0OY2mdeffkT4LyEHSfQntz3JfWBTLMzJ6PSdgIFcihSED5sTKXNuFJHVJY9
ZqiKhCliqxQs8yPoJrm3IvDlP3NhLHtC0HnahFvzIv289xNeOqUuGP4v2JZ54JcHCOwVOo9xG0ad
jwe3qktp7TTFmEU94vrddEIAm6gjt2OAK/SZJlNIiMIdTPeyVWic+wnG+6wyVsWLRhhzoZmaJ8Km
QQtQXUqUS/tssvJqsrbJIuqnfUQdd+ZdegnDiihwJir8C2+p6cadvsQ4f/SmluTWKt568jyOJGIr
OCusJLlmOIA2fZaD/lO3TzJKhNG34nOy7I/aO2T3vHA6DgoueR9cHyDKDIt1P8aKheoaFdLY94mB
nO0tWqNXKmSCyjyQgTf3eP5VV0ES+h53ufdH9xz0GGEWo7wA7brSzWeBgb8JcXJbWrprHCOczkqJ
7tv3Q2h4AMsiHQJant/NVUzKaFLP9DD0jIqBrrSyOa0uliWY77yi2YYTZFnhTMjI48Buz9ZXef2+
0Tc3B4G6u+gL3811wOSFLCfXCIKlhqi3dFqZ/h31LIZ2yoJ/Iul7YO2nl6rd7Vx+/ChxOzOChzD4
33xFxGCfh9Hf4bsKMAGxFy3RpREJwiZ0tqE3grbLEUyxwQVHbifmIIF8M9qah6RTGKpkxRMk5QTO
0dN5y/Q612/9ACTNoH6qcmSzLwsBOHz/0x3uBDfK95YikhnAtYlLz94rJxPcbb+yTVDIn09fAGJh
ixaQiwu37jVuK+AN5zUevMXPE8lX/DC0hHssIeX12Iq6iuj8TZO22JzvKSZRr9xs0A7W4Y2XDl0f
QZ+uYSSJ3gNwJ2euc3P6yrvlnJoJ5fNKd1n5GEASY/FLG1WPdrRsldYG+F/jpf6gzbeXIbN94N2J
BEZv66lrk+uX58FGecgj7Hknl7BiSTy49Khh33d5W19B9s+8pd/XptBcSxiuL1IiJEqrs37CSyTD
oDCzzjJ3/jN86UmBynw+qFe/uoxe73rjhgr9eUhg3vKwIg6bcLGAnUbHo+s7rYFMv73IUVPnwSbE
kz3pH2lcRe6z7pe28MrLOm+0uTbHELwn6fTVsxUjjgETLgex7btB6WtSMzwoc6xakhz3U//6YPtS
EzueysJJpEKOuTGtdBkxVXjxHjQBoUd3ozCOEyb9DFUvUxFneCQf13ueaHuDC3PXHe9QqtlEZqwb
DmeXGC4etQIlYSPWjLHSnn/IJGe0bjkmUBu7avwfsvtFucoGYUZzaSk62MMTbzlJ+ULCFv2cOCRa
fSwOGPeeHZth/WF6ORhPzMEvWp7zExbbKhud73PSSWPHTi33r5DpRQQIcrcl/OWtQtHJw4j/QQIF
/KaqRAA52oTiAhVQhfgYtvMM9wfu9+8PGXoHnCfp/IVb++osMplHjqzn+9SCI7S/Q7LWRWT3pgY7
1bJy980/6/sEF3fVD1qfhqUumsqWKBmVnIo2KSv/x3W6Ydn41RWusubNSPxbxisj4MCZtXZte8cf
FVbUdCMdNNt4GZoruU1KFe/Dpvg6QtlRw8/iM17Gtwz+3mC7tbk6rp1qyp/GaoMqg3JNSXtrE1PX
hZBqpuWehsqdcxFUGiqZb1yhb9WJKP6ztfLidZBeDM8XNccdHfuFX2LcMFa3UnwKmIqU2qx0ocgP
XYj/tGF+vLn3zR15fghBZb/34Q1aTn/3rFij28MDvduJBqUzv1vxv9DbbmIO98hwfLuhG17N9mzV
ZC79mlUIm867cMPJm7+503ySIDVbRNcWRAXtuw8XmJU/upCu7h3sSZ8H69Dytyrc1Uff1roPMhFE
46GPN7sk4NMSKw4WUaIEbFC3gLqP3PbZ/e1GYXJPxOCYxyFINmUH49raSG5xJ8V8zl2SEaCtNwK8
Kn3AUHjEDm0TKA5OXHabWgB1asRzp8/+LHAbuxYpsraZkSwRC3U6f0wEJnQp2gvqpUwFLdvZG3uP
GN1dswmg9bbopEQjkm+OcZNrRG2NM+WYoUcYnqJyAWYCs2nmVOfnuzW330v+tBnQ2fIkNigtXZIU
2Y4wZxKMvteKoKvV8LV/gTH5PitrNFCF1T8DJf0tVs60izOOeiyeSKZjFSE8SWjS8UVOqVIvBH7P
DL094g0hWAwHFoE5LB8oIDtcipGm6mZHN3D64wURh61UjZGTiO13n3cW+Vbm5YvwLCG6a8kTv4lu
VfCPVF3n4+hPmgPWgmqYOgXswbkafJ+ZgQr3nt+3ts8fai67nj07JIZkPezyhi33mw19+7pFoViZ
Re/emPdpt/3hU/dv/gQGXbCXOSvnVe0VVMaYLui0DoXUXZYkS3pCsgx6hg94i24YMFr9Q5vawqMb
fPrrZ+/G8NtgdcPTEWaZasySqS4wpMyGQPRcGsErcdCpR2dVJw1IeEHtj6+WcFGFlPz1k/Uza8DR
4FPtxufT8MyFpe4wf85OyMKrXOpDWB+SnapKhrB/Btc+/wlV1VWuhNCkNibk5RcvFKNFa+WfSy6B
2Kcb+De/4VL3mmBMjKnOZ6YxdirbCv3DQsZ/S9Q6wWAA/Y/2dKq+iHd81uV5AA9pkjGt75Jw9xkF
3mGeCj8m7uocdk/JZMXVldrq4oHj6Erq5ToKqK3o9KUQWptzurTYbKtXCrcE/0DyAty+fOnktJPm
QL7lWPMxU5pfPz7KBz6JwZMoB3OX1sqKI8cJv9R5wzlhPrZEAZ+w+IPL3F9RP5mijFU4FhHFADcc
4glnGjLK34Wcmh2ZGEWKV7UXpVupdmmM9umDMGvIYxiqJJGyzUx3qxjmRe/lPytdzi+czaHMB6iB
CAd5T/Knb2j0T8B+wN+LYPOu28XTVHYPC03mvp2Tm4Rh/EJVPxvXxJFOYA23c8FOUg9zXMX9HKGP
LWDGO56mgvidCTaPMVSSxXeG8554E35X6l0wktkfY4C5u+JqGkvC9rICiAzhHx9X5MXbz5LHxafd
pi1YK5Q/pPjewMH9wNVEwDtuqR9HFP39sTe6Y429trAZWCutAz5ZZkJiVEjypSodT/hEMcriGTX0
Qe+moGiwXBwXjAo7KxfGwE4n6+v0DZtoEP17QMd4Kth59+7pFANbNd6KW6DgIWcmT9a5YCaTy70X
sLrlBOqYCEh7arZneWxpLVHBmg6XDLq4vMqu7seF85T8FydNi24+s5oUvPc2N2e+Lh0HQ8cW/Ksa
WyXnFmZ5zH4LHFiF1Hgl28aZjo5Zuss+AjoiJyK9ONx0NRV2ilrh1RxmpMVy3aTOEXsxUvqNtgCA
MipGkso059W5ut1eDit3A9cNnNOOuRu93CNSx5/D/tRASqezZPm9s0J9INLCISrpjaitQrkHuGlF
Lu6p04U0fBegWQC1kklMsD+QN4UYZhsrZugLwuy24JMq4BMXwMgrgOm/ZTZZJaZWh9GmNKFQJI/y
9YCI3zRQR1n/AHTa87x+LBG16SyLQmFUCEJ9WBFMSjlK/gJIlSYymcF/99yIAhP5+rJzCYuduona
T5dCQpvd76KuHypFwXTU/FKgjThmagaJX5Q50k0fr9yjfIQF6IqupYkdT9V8IGFvtelJbuoATUq8
nkM1bcMA0pG2CzctNLMng/UvIswCCyBcCXYOJxdWsLtdOhAuqleyUWa4AmicDu/TQvwTGtILE/6v
IXfhT5gUd7gHL0RTO3PrrY1myYsFTlE4us82Inilhw8KyqejF4NHR/zsvWyuKtWUV7Z7lujLqDlb
uBs7YTid2r/+uL0bmEFHcuTeNh0BFVQJM3UK576QlZEnfvJv6rDu/KIUwwoa3bo4tlBH1y5fCkD2
SuEgf2dBvIp+uWCdKK52QkmZHYTbyFL6efEm03uow9icn/EiMHtVblTfBkM+UjkAo1A6eSpDpTM9
GByABK81hrb23tGIY/nxaweYVXYkcICniZ76x6N3Rm6NoNQ49MTPzyH5uP016u7fgPwjmMLa49Er
tQS5HAHktdunSb5NC4Bo6NIOEYSZ1IRofVBghL+Mj5Nzk3dofXuaNa8Pz4hHZYUJor/TpZXDTkog
H4Oo6QsNGtIW8NREBX5ci++2D6VEn1CVsYtt9hq1M64ambTWQRjG1O7rgjj/JUkxs/y3ZyRMx9Rt
Jgcpeo/rhBbNG3GbHL598uhAIRW79BIaG9NvKGqaAAPeSwFbv2XWRlh+0QF/8CFiYX+/ckaSscPT
rCIAJTu8yiFbFKjs+cN2HqVRxAjOTeq78BHc7YcblQrK+5bw24Wg6IwgV4nmRjiWXqSoGaWeLedB
ozSxHjv9HN0Poy8G2/x4awIc+ZpdY+4SXHLl5ID7mT4vHLNCTDgIoP9vyS8HbZnHGJrzLshjtPIL
/xa0cqPFqNxCgxE02pW3yECN7OT4AFzVu1NhhF/I0nR3PHHQ6xhsXVLLyTUu9DMEshLD/nh8hoB7
2ZlJLnW4KkuZe0vg5ySf/0TOIUxabgrq7aQnd7bOSoVW4Grwkyvf3YYrt5ZK6Lw8svynRCmMAh9s
rto9hoQjpzpYUwmSIrzvLZo1iXvRhILBLRPyEHDJ1+HXrgTm+ZrvURI7ZoA6uFlslqTDheDAEPNU
V9sr2dtOg2Y0tcB9l9lt0el0FRMNktkVS4McSsgzj5qiVKNdKBtV+/EFRaGph8F16GqWkM9i0yQV
jx/h9qQQ91SLgsbVL+h7aNP1DlOP+hnDX6FT8XvUENb/DnlAFxraVPe/Yne+/6KyQTnzNpLlbhc+
fi8ABx7mRf+zqAHEGK8X2SFaYMOL4bizatyKtk99v5i2d235FnVR1HYYpUEJVNsb6PDE6z3LzrJR
uw+l8QAb1x16WctTzknoNF1wKIPFFkx9ad5QW0XtQarBrzp1OxCG0fsGUmjbs1iOxy8jjpzMfzkG
HkVDzyTE8fbXEk6kU8Vdm+NGMSWXedn9FH5Na8Ci9jAQhUOJSKdhFfNKO/mqNJ5r36+NxevmwNBM
GdJry/M4gIPg9oN6/txGVXDMY6ra352njIdw1ezmAmIuGhNu66c3pJNnX/4tAbOI2R8KSTwtv5HO
uWuWK7uLHrwO465bBNrpzzhEh/uV/m4lq6bfSoW4080gKcp0N49sDskwgiik9ql+058OwwDNMeI0
N5RmlXRC8mvDfc4BbFZMrUxeM0GG/TY/LZ+G8QYlJ+mDwK1tuLMe85ZQlR8cVs4VZP3Cs5RTSXuX
Jj/uTi83K1iFbtltm58FFTHInbd8EACTEhfUn/VohgoEUGlYGIeDfBxD9bERLKT0rqNfZkNBpFSD
B4K6Y4H1dkNmiJyrX+1NO8xKBxtim1TOeKk6xPJ/cBovVqGEp4VXFP96PYwsbhcaaK3CyA8Xtfgy
WXwhSqKeMJeOoCm03yNjzuxLO0s/ObBz4A3iElfllyp3Uwy+wmz8VaS+WuvcOssDEASlyB6BOxFE
i+1dNXTrg+j1WDV9COBXitSYP8d7Gk/2rAoM31Yi2qc7Sb1TO2RR1JK5F1EVxMTb/J0qeXCyirsk
MfWbr13mV5VHKRczByukK9GBlxYXPDbIsP/vMuZNRUAfEy7aJ2nZ95HqJVX/OdA9RfLcPOY/9A85
4azoa4h35RKcijSRNgbG/+Fc/pB90t3OjrfYXLC5M8bHMsusHSM9k7Fa+PEUkpbZ2adKWba15dbp
iKR3itVB7nHDi88oeWDD9tI4ZJ2qLpIcl2fhGdKFS6nLDTc885sCvnnKfBuhy3zgWE+xePoN4rCZ
2VIeow5UjIGWvGyZd853ttO+xhT108+I2z+XcuwLVKmt63Vr5r38/hhx930zsB7jJ41MNjL8ArPn
NlxADBZO78yo+WoYi6GclcJL/1ZpRRoNvpEGIO2d6XtJA9pzOI6VcrQQLXgYbGzjLCQhrEyIG5Xo
C2Q05NnrADccdy5umlE0aNLbvvr308CaWIiigAQB73X11QzV6BiMjKQL72OJ38wOnaUsRHaWkVBJ
Mmd93FBdWnUaIKUpGS2rs55JUt1WNAHeTdH+nif0j5OrGF3wrp1p2Jura1xnDEw2CHC1i9bpQRHN
2Fskd4lIyO0lvktqTmBJ8/dvlP1IyTn2FeKeYH5tqDMNTEuWGVyojm2ZW7tKQ8Vy0+1j8BSXobLG
4h3PxUS3NG9kaYXJ/VPRRgQiE8tzNmbU4CvRzefgmGuCmt/urRu9jUctLKR0oIoLRNIXTog/qy1B
ux4SMRaC+A3v2g1dmc9TnSIsIbDfkcB0XGBQ2v5If1E2CHjqszcHfDmis3BZb3YDAajDxdeLlQo4
zg5rySsZT0avNXe/ZRoOqFwNOZj1sC5jSdnS7pXLdUI0nBsPn+FCsOzwBpd0jjHIWrENX/F4Cbiy
PcpgwFXv6nKJdqT5VdY/QkqgA/nUvv5H8lgbJVP+Rl25omEfiP05a3gYcUXmWkRjUoKLr4oUcokw
Dzmn4Tc8vlzikrZLbZDsSZ4m8qEhWxleA8e8aWwBslxVEZmlqh/E3MffBFIQokbvfER3EvQAuZe+
/seZL0q92G3q741xY92pCzsY3ctIA5iwpLwdBw2FJp9U4mPuckzN3e+rPD22WX1vCRYx5G8Myrve
anSGoMs3mIBSHPn2U6WYCPFLwCbgT3tQaZJO6NkSCAcdfjoTG+d05MNF0WlMt+Trc+Z787vHZEyt
2/FQmteOQ5Hi7tqsLLmF4l9uYI0d6YjHg/fTrckEiJAtBLajUYcSKXbWfZ4Xt5Pw3923UKkO/aSd
+kiq1vMihn07H1Xoohfxz//PQfI8XS/SZmaJEqQQljORv9WTazN6DcRWxn2XPdgzhyjkeVmqkC9e
UACl5wTfYc7xjgJaCAduj5YEjfK4ATN/22KA4FuiASHBS9FYREsvAf2XhwVZ2MlHiFLXWDJtKZsv
x3hM6SZB/OvUbRCqvsppEEy+HmK+Xv2O8fUIMU3qJp3e4EJPOHgD3qpOm0M3Xiv1viwI7GEwlSv1
VWBS09vePWZ7a17PHvTMgFKx8eP9RcyyWJhKOFTWPejtzG6MgGCpybrjLcsE8wvZ5+/OHfnPmHQ1
wZpN9SV4tj8RVZ0+9oghMWYIdxzsYlN77ar1qItgcY1vNofX71bkh9ApLCeXyc5E1bsu1p9t+VSa
7pFLB5HiESRZyHYgN1kSxieuSQVJeTcCx+TpfbJm9Azc1AXIsvflOsRUyFeWxeSA78be3MJzniS9
S98xfalYslurqDLWOvQ8Tcikwwb8ckFqD9GFCEd6p3t/Le3y+7CkP8uWvrxMb1dIRpwrCbHimRTk
ulmKhj+S/pii2i2yrEJbRirz2neDUsypbk8j/mZzp/aap0LK1Orj8PEghecudu5Vssv3wQEGo9Zh
ZWm4QBFfcM/KrWYlQbcn5t+IAy6coCJEkGDN50n0oXroyYZZbit/PUXwVdU24gaoJ5z5eeBPqJ06
dtMsXBSRGSetSy1rvmB1T+bKgGwpobb2NcZQ1BhnLOm1h6n4egI4FX213cMHOdrJbfNBCpekqksg
qQjDP/EPIdP84ZcVQaCNEWJwD7MMNVtauW2ZvCSDQSu7sv/G2MQemDHDJ7gNWqfZJYv7HJsl1ee5
KUfubLxyv1mi4/PLraXHUeU8fiKiMrTZk3LxppFD7IQsmVzwuAuxz1dtk3lmy2g2RC21dbhqkamw
sRsfrXoHCNyswWy6NsMtffYjmH2cRY8P8R60wxsh/zy9cUQOCRZUnRgo1BFHf/Y0/BRGT6yaoGLw
qwy8qWxjE4xclcvl0a4VQ5IKVcBLocbjlEZDLsWLiPmfYe5BxJnRjSI5ss7ecT/laIfmfLmRXlqT
/YrnS7KVyPkKWYWbEV6+ucT6xMFBUu7VwbhXbIqMG7WcBJsBURuDSuzQm2KRl2LpCd+xDKR61Kxj
sPBhseu/oRRAWOZU9TdiiGWYODrIPiuVlFp3u/bCHtPvcD+O7f8Igx2QMqhaqsgI1PjVnFTN9TaX
ai6oadFqu2UI/h5UBdSqzuiWeybj32dpE0a0XlVTiV4ULmch5nRYfTQ6HcMKTDhHaYNKjNNJsUSi
cdUfkcE7JYdDZdzdf3uYfnVgSFEAn1GqWt4WYrmr1W3fKzXV5tSFBeQxfb27zDueI6kALdKmXKMd
xG9VfAyTXAfi6jqLFtP+KIQE+U/W/jzvym9Mo1fqrC3moXoO4CJHfZw4hl/YItsAD7S3nb9uqohU
ajXkDH9tN0yQjHLpoLqV+Hq03pX9gMRSAKuFMlFKOQkY849QNOmrxaCwqvaOhXNUaU8/RUpAqRCT
ktpPhayQaZTiNcPFkN6H+UKxsbsL6XQa+ppK2srJV4CIbJezJZ91MreI5E7k2McBxcsAhTC5U9wC
Wt0lFHShMOf5Sc5JEkwyPJz/mzB4d4ZcG/16JaDtO1Vsza26qBcC9J7Yx8+mYqTx2+sY9EZwD6zq
k3ImI9N6XCMqE60/NnI3x90yN2HC3cZ/CjrM4junQtHuS9cwhkK3AvwuUMBBLsH4pR6iRTGxeMAg
f6k/+K9nmQzuedszCPKU1217MhBppGAUkxFZ61t8F8Dwvy2bp8gaV7MF4AgEMJVvHmFxSeHAalP2
UMXgkZKwslWCrmiOL27hiGJOAa8plNpPt1wVdPDIU86fwM4S2WK4WaZ/r+uGEPfo5bdDykGcf+i+
3iZjoPWHbznnUq1tH22r2G1fBM9TgzWLFlrgJPuF9Zs3v/B3dnI5ksOQ4ywDxf08enpQ5JIXFUkq
6+xf1GU85WIN3kwxHiUz3FfE9XQER9nRgn7sJTmuE6w5biZQtsp7+0orvtOLrW5It79MLDFAYPMO
E+SeErapkiKK7C4R0xuuucyLZlGD8cL3jhWgrvC3PYzZsNHVPSdf3bKsmqCiyttNcpqOOgJfDbIa
G/Nnyf5fn/ipZ2h1Pv6rurWuydhxGli65JDXYT4YwMpGrwMhBP9H96tvgLDE689XXoghygW01gby
/+q+Gp57mOmmxFIzbacUCgvRPruLsfhDXPNLbDikxOKL5CGSBRHXFRdeVc32W20M+BUfIWLohZPt
EBOoCTAWTHTpDwlDZzcT9kcHhNtpAO6NeGXYJpYf5pXwVPAm3hX9+HMlvMLSDAHzvM09Fp9j+Itj
tUMJW10FngIqg0eKJ46UqZqJPiPTqTVf1SZQp9T+hj+i8OHD0MwxgRy9hKKHYLE1XtwYElNSoKRG
BOgmUf380dvuwBDwi2wsjKtK/evEnV4UfZ5CK0EX9e9ptwbwp+VeuAhLiImBdN82x9KBNvYGZK/v
Ga8uJfka1NMDJeY4aXhGB7pxJbk1dYtIkjzBmygtz5daU4BpyrbNajxpV87cEZ+NJBfvnLe4Syzx
L953sqx5j1X/9pUYh98e0rdwBVLv8Hqb3aTqHiagzBvHFlsee07s6PVu4J5ZBYHven520d1oM30L
uv4PXc+K1Qpr6za+7pcv1GyFzVGagaMEZjZXv4l8kbj9BIqSKT8e7rHNRZD0QVu91dVo196yYnIw
K8Tse4RE6jWecrRhGQ/p8qRX/rMb1QtPmOvqKZCA0A86ArFr8elK4F5x1tCiJDRJapE/DfZ8RLpt
JZ8ZU4AnmhlYimQjG/yoyQoDD7pBt0gcKeX/tioX6zSicKJU4GDxsmXumIusldnJgj3byrEtZ8Lg
ulqDa048P6qUpy5wnyAsSuDK2ywkE4qG07PCwoxYtN2u58I/EUQPyTc5tybY3wWoDEB2R9YB6dok
gMVkgd3y6e5Xw3kWbg8f1A49FUIsWqj1R0Ys9+scAOkGDHy7yKDfX9z6izenxpKV90QPVH6JzPkM
W8nsFxQ8+Fee4KKdvd+Wvke+hIfL3anXyF13yYElvem5i7uRRKHI7lV1RF49Vc5/OAP3I5yS0Wah
1KgMVLaZnXNy5fZZghCShAiMy+1UrnGAK1sb5IVF9qrE33Mq2macOUYnhwZVthhUxp1AoRfcTbBu
FrQiYp+OCYfevsJF5xiR0Z2fRZ6ZzA/VIozDdqKcX1P8rF70YUAkIHf3zMn48+GW0JtCg47rYWjv
XPLdji/65LHX1eaM89Cgm2FeYBlBHQgC2Tn0cC9MAySBl+/trUKO4U9IYW3YLJwXkNjQgrWGG8eQ
xAr6+qFEt2LkpW/fIq4mqXm3U4qjTHICxwr/i5O3bHw+AeT61aCQGEtStJgQbBFNnQHoxQ2gIlgP
WSU2MGuio8Q00KyBu3C8mV8R1g1NbI8G0SzDUxmXWNX34RoYX5CmnAhe/E8TBW+1q7qi8R5sxQ4/
OB0oD7LM7eaWKqdfUCJM7Q5wlLiOxEIXziY2DaviPU4Z6vtbSzoSoyCBR8UKnsW6ez8GZt0RLWHm
uTGVOb/J8fh/ev4Pxw7UU+8Fw28tGLtUBbUENMO4Acoj4tzUDYc1tXsF8hRh2/RuyI+XjWgvFTTW
ZKiAeJfK34R8EUphn0Qyu+bn4ne2zmbTg1IJWgy3tCQ8Kw3oG9RyItuDsN1uigKURtGH9EJqrmgD
Bq1OCE12vFwUdc3kt+kG59TUBfJHBcFXPcxl7gQH8hrHWKkPof29VfUNSl3DqmcqqBp/dwIvSbvp
KFiLqbfvlID7Bo9rW184VVe3MyeQ0dW1Vm7Yw0V2uXvyEaxhBIddy8C9cUxFpDSPNZdag4lhasLK
+w3rQY/xeizCj5plMW0NXhml99tA3RLFE3L1G7MCN36ttDVKTdXm+oH79YMOzASECpBaL1oXHB5r
9Rou/9i/rcXUQdYyoZmf1f8PDXqegI6ETAG/jn9AVRDBAbaj1NfQ52HC8ZuKU+mVLoW3D3VCwdLl
7ivYAlByTcnI4HhcHf/HAG3yt8PrCNUuKG2z32DQ4fCPiJwnwUXDjr2yh+QpO3gGjIiEAkob8IMs
Q+Y6vhgk51Wd5m6wkyYMS/WkPCRorWIe+cZsFkm+CK8AweD7CvRd9PRhl0M/Nwn/n9NQu28mA7RK
hcbc3NG+V7ST19ER2ttD9Wrj9a9n+4yeB6mn2jcH1zImxbW+Tujj4lLdPnSHjSPAb8S+4AxkZaIH
VLodLEsPD1EyGQv5SfKYX8gjlUhyFTaV2pOiLPg2uTxtzZSYp/47sjdjWIgKT33NBRTtwXo7qBOV
8SWDFqc7qFtE+pJZFccv8UyY5C2u0E2E1lArPOT8ROK8MvNpD4jBIa0RTZywvQ0rUlzliSH9LFG8
OMu3d4ElIjDdQc6/PtHbzOrlI1SABaZBgqEK34jNpAxn6aw0WuH0mkgNTkBk73IoBmCQmQ22JBr1
B422eH92JnwrIQbCNoVNQafLGubvl6dZTp5TUVCJc2Jl5kH1bNTxqL7dlsui03vj25spYDpQqrcW
3W2ep5HzhG/qEbg1/TGfOO05t8EtGks4MaX3TAs+1bOsqXpC7vp3a2vpjgv3U35zQnVVxjwvlkjM
PbytLwGJgZH0HBs+mLkkSAi4Ff4GnFtgvYbfTfK7k2VNEccfReNgfvbBAYuS5h78TPyehQjk80I9
/IRAaBkGmEz2PBM/VppgUGNOShsf5bbAkXGVv/zBKr5iSTaIElrUvzGv6HlysnCmekcPBusA8EXc
WhIM6e31tDB8VsudBD/904gMB3W4Hnr+qomZy6uihMFSdNGQ6ku+23yL5hy93ce5MRK5oH76cfT9
F4c8sBSn0GxmQptGvLBH37De0BA1qUAn/XrWDYe7ZZUbsS8PJ9MBEldVvnejDRbmz2RvzX0exjCS
158s+vLrLtdws7g1/yRlRRT0L1uXOTZuFeo4SrTbLBxqztzEqoO+h/wQflJCgPetEz7v11E2Sitc
zYhngdnyzmnzBfCDSs4gUVeKcV4auHS/kb6TeDYkIYe5+zMgm5ks8RaUNraNAiCRrzYOjMukUxHt
srteQcZ1xGe3POLOYpd1ITA/CeQcFhf9Vz4gCaCIRuM3nPy96iCFlaaDm8V3ZHPG7FPsU/cjWw28
z+ry3gb8CxKqCnEf7LbURoy03RLMt7hRAsYqAhHOhhsnpC/s3dFtoQl3U3c3DStJMZ5mCGlSXWDC
3O2WDcPEHsCwO875RhBdNVps+DgZ0Ttwa24rQMPDNbAZV+Qf5XrPsGPlBYtjq86S4CCXArAaM3+w
EUD1Jpz18wxM4mLOEhfHqCRLqBSFi7doHMd/GqihUXQDiWDq+mIedLKjrXo56pVDJxjaUsCWh2Ud
w8nNmsjKZhzN2Mj8uiUQyblnSSPofADSpxqLPFYzwciu9YvJx1YD7GIbncX4CK7Vto8ozdv8PcJF
1pHWayouJWoLEliHv4LM7c6ZWIeDfHkO5FkTKgW6bw6xeRDiBpleJi9gsE+bS1qNmu3epd1hwkV9
4bPG5VVkvlI9MB09SvOw1SVhtxozOs4kb9Wmy/tmQEakdZ901sa5MIdlBbvAEl9FQ3h7wHQYa4FA
WsWsj/R1vrbIiS1MYCK+03TPnoVK7BnY5Sot0qDgPNALAsqIbahqgokpNC3k1VME9eoa2Q5m/x+W
5PnGD6F0T3AIBufBrr1rl1LwtZ0Znk+ixFuL/8GfTCQvdCQGwe8GmhhjG2mMObvJBFq7ONou+HYF
Pih+DKmt+KfADGydh72exnn+sZ3pf7NFRgfltcrDnk5slEEZLzlM9ScXCF7R4Y0BQT+3/86te00M
42rilpHxiGMExHwLjiB3hFW/KBbnGhOBLEgEzxWKRxHApyGWp8TSbh1WihmFJE76ukgidEsTj59i
059SGOf1CSz1tIiXLqz0DnNVC8kmgjONntEyPHxD06DOgYGQggx1tP6Ig0IXklWpu1SvfjHmGu/c
ShAuIzCj7gBNrp8rH27rWqkC+/0ehUwInv7BjzznGk3nVOwrcIWJqkIb8pCV7EeWRwQPrfxlhd9P
+TNuojxPCFObKRfyH6H1mS6o3BAG1N/5LrupFe4FDLelSoyZ2WgqgIHgz1konHCVVSegQq8u0eFI
ucDRkybuHnpzpQSl1JnqKmk2io9XrCfBdq47P4r2cnn9JRnphW2BG+MCtVry+icGBa/a23853KhH
tNHkSQGAKdKj8XzzwCP6gKMKk3HtmdgVwapojFpCrJoZDCXU6F774bVqkfEFFE6QomM+CpIJWNPl
a3/1g0AllkWIy1lU68ciDbSVPbME7CcQj3AyIpv5ZrjWRfNCiv+87c+7Vc3tJ6V1PgAmWnFRjNxi
90McVwjuFajSCE459uSDLYePoEN1/LJlUy47WIBAKiEzD4Wb5pq166jErI37RsNc63jLB/hQbQ/B
8ERzFoRWmCpEif4Uf4/laqDioIOJLRvsTrJ5WQk1OHvplWC2qcKRh/FmM/X3n2Tg0adYzlPyy2Xy
/5p8LNvX+Pu/yIW0y444J/6KO40cuQLGt9GzpE76PC8gZ6Y+l+OW4d60lgaM8DlsDbaKvobaNxXm
eUUK7qeReokwu4Qja4996z/Ta/73ykiEgpw4+19u5ZQgAlYimU/27yQCYqpj90RoAyUbpx9PS1Mm
l9g19/Yx+1d0NcLBJcjur0KIolFbkdeJa8RxyfKAKwZJZvQYF7raFykRR/cuJ4MC7CCh/riUc5IT
ij0ScJusesmF6J0mxdmT+TsiPbu5iUfomAclCVKi+a3C8RnGsPimZHbQIY3Oe5oseN8LhwwEbXwT
U356U+MxiiPQcjeIgXdNpYp40d+CJ+M60tcc3BaqeepG56g1rTmXl7VWQSRaW6YvN4evwruu7w3N
h6SAC5B0GhUQv5rXO0o7kvO87Ja2+jFnIL+lwz9XnO5fxqU0cGbruoVQLNZNqE++rjsIEH5UysnD
FXRjKIgY4mEz3mkQvuZ8lnRGbzGssqhh8RGV9Mr41sehZfSv1k3RlMkvklZizPqnYu5j3usbe0bm
Pr1QnPlkC4ukipA+IBlnzGz9uW4qH5uqACzXH+tRfJn2p01QX9Gdej6dl0HgEaTVL2RZFKdYG+I5
52LIpNbYi+SputgkbCYP4T3vWHUh4nJFLrhOBBVgrEa4vclr5RyA+XLbPS/vzXK2BfvRbc4bUUK2
WAKlm8q4TQG8X9x7ljLAeYyR2inDrNLjcd1qL1ia5O4CTJSy9by1br1ANZuzePLHH2t4AlmkoNoH
xOc5+7zh3HYTOYGAp4Bd/Lt8vd1GVGT0HhKhkaBbw4dgHT4Nnozn74HaTvR/24mxV9ftStNjB3VI
n5oEpKMH6FI9w1H8xq63qYBdy0//BNMlAjvzotn4zcbzhDvR3kEiNwEiumFgaHcSmuqDwhIJnRPT
+6D2iqiLE/eo1aFjTMFB69BLw1aF4atGBXZIWQy23lkPqkMoY1zvotuVwIKBjGJz9qaeLo6MXG+7
Vpcp5BsVJrNMbguPSH5IF2AmsT9ht9uPcjHhmvUcfz4J4ISieoFV95k9ZxNVeAhPA7AMkM8BoExh
nkxIvqVCc/rZcZnmnb36+muxqGoyfPZU59B0ShpjXyjFzAxldGeqeLZZX1LLMqtMnArT+M4tbhNh
kTpfWrmfmV56gKWNHkcI0DtdcJiJuomOIx+c+pcV6sZuODgNTdFa5o6ehLXobbX+92jDxZ1eFTX2
ZzLdmCF+HAnsa/pci/OtW4LD4ouHTh3tD+GI6jZ4B00wLtksw7vGvzBna6j7c30is2JM2qiGro6S
qGCbF7vKQ60pUJGeONdp+EWYgoVB/zmSd7sMEMmZTy5ve3fghC1rqwUDQGSFDNTsGQNAwPryoqKQ
ievq4flZg8uYIX2kZF+166y6S8/0VaC0TWjIR8QkakgFY6pD5zztV+ST8RzPGTowmjY7xanOWLzB
220S4XUB5fZ3/44R0L73T3VZl4yVbKuWrG24D3eiTzxgJd5dCH6aLrHN0yS9Epl7vJ+QMIDzbXKN
uAMl0OCOUQ7NStbpWbJ1ihgpStLlQKehJtISkW8TIBPAHSaCHSGJuf2eXvmDLVDQ6U0cZ9fOI4St
/sKjEXiCJwx0DAglKCGkLSuVGB2WlQSKG+Z86/J9eWzBXu8zw9e04LVIU3rLlc6HtFkjkCIrlazX
ci1uGcUkj2KfVtOkoiUQ4NsQF6Um5rqyLSeYyXuygl87dYtPPkA3frB+OjRkJa95WhcpwpznW6ty
Ixc4qHdmM8BjSL6h7SAXhRV+YeZsImCclvbBZjIi+WDptRuvs17xtxHwi7jKrt8sk9zmF1LvoXl/
bgiymZXHFmZNHJAG0+pZE2QQMnvGETymG6RBDO9cmkzCHXE7+VdF4gy15qWB1sbU/dQt/8VAVGBA
thdDtwiLN3VDEMInOPuOqLG2eHS8M7atYpT6yDLmTFiO1h74lvgHbQX+LahhvBoMw82LJSh4ZUap
CUC3Xujoju0ZZR1XEACV4U0SeCv9pgafB1bZYM3V0ZQGsWh5M3AstHm2DIUoDLH3JWV31m6HuHTn
Y/fYRHry8CtiqLsUsJdBWTRcnleO+QY+iqash7eLi1a+7GjBrLmFpvaT9PpKgsmi0Dfaa38JDKJo
mCXqf4+6u/Xm7xIRGKXVA3taUUckPZf7yEKxcaSccVgEB5b6ZqfzxOXd4obRJKXvO3WPjUZ25L+b
X3KMG69pM/k+/urHNb3DKEwjudN5PGUVoIQ9LMAniI9053ptc4cFVcaRtbnWTJuyvVAR2qRqcVUe
X7nAFKZWzjyzynVUdMc1jObkObdHnHHU9WCj2NOWFteojVHqpp+UaiR7rE9RFqjldq8VTRTdHnx7
o3TUkoLAfJYNvFcc06oJmUly7EOSZr+cItBM97Bt9x4DOtKP2l/rFZofILN0MuNJzaaG0Y/Hgo6Q
H9RrqlEdsyDT59jsAnGlFYBKbsGa4MTjWX2MLg3Eq6qD/VuQmRp6XMmiSApBXyEP11yXLHr2ktlg
zllePskDV/mHU5VkfEclu9iBBJLkGo89Q4vBUfdDlIxlG3HuQ2OqwT0S0VnIZrD4I/+N8/dSRBTx
HsyF3LcvMkbIw0O+Bmy5DRUDRFc+CG6dW5m8wp9zgqLxZbX6IyXsjnC+YZw6JvDhWGPzSkDklqI3
woiUhhmtKkyhc0iPp5LC/WDMszdcWBYdzN9EGlYNLzVS11jFAUyCOI2T1qe8x+NesleS/HwCvwzn
8hzE2hrsZnuPZcvxavd4rN8g/saTBhpXe9ChrCZSLtVX4NpMJ4pol2bSyJDSMNBCxGFoYhSQ27Z7
TbJhiNyZe7ciMajbk3hS28gdkdIHBw2H1ilLNqtOMWu/FzV4pqbhPzO/0nrAO3RxpJMh51dCgXT0
sllsV5j0oKB2FMrILgY65RYNndH+hy1RIUPOcZYaAU2qg2zdobluWhuDO7rJF08gCUt+7Q0l7NN8
faSMV+rP25mvexcuoiAZ3yw5L4pnzSeNYc/QAr5Bu/XHvOy/Vl03pg/8ALg0z9ZccplyStEEvPNy
TLQ9lnUu+T777J9yzDCCkn3CeFL/kdIxA50ndEThRv69drji4xr+uEZa79pEKpmBjdWpuiXY+CJT
SClYh4ekkfEU3Di49XedGksrJFdhTtiCxZhx1vTiV8IbCJxuRShv0nRe5z5L7eSkcxVdnq2VH7Qa
s+23LeoazE+/5mXpOhlbxJrTzdFYIXrQtK2rD/LfUCl/u0pbxlm12W+dFv3WcVNHOgjOCW8qoCkk
zMmRdfZRaN9Xg5iK0WFVM6Mtp2O1vyJvfvW7w2NOqumsn1OxL6OyYp9ggJwWHCoZY4IjBzCFyBO3
i0uiURJuGUM/ufhTYQeshbO8r4sD/wPQJhfathAmXi8ov0BJuuyIG9nQ4zZZpY/OtyofJDYt1oOT
xHC5a+PxTTNI3n4UKl6qqTjB2GjIRj0+qn5lxAEsF2TE5lSDSe8iv8fM/DJllICWLcsXvFLLwFIO
kCLeQAQy3yu3QXkJ90jKmcix+iCfwGRH6/1XXVmlO25+8LEKfA4+Ae4kQoLmC98VHIwnQyJu8Y4Y
G+PJH0sXfdjqelHapTgIVKvqE2g05GXX38xU/8q2l99QsIPmXMUwL6bTTqmMOwFLmjFKiLXzPs+4
nSboTGS55Rcy7FRPaUV1agaV/xtcWu3lgd4PnmDuxZAYcrgCuXo/lyhnH7jUfCyIgM1nwB3WUrB7
M3+k3Sjv+LX/nde6GrkIRIXJNvYvxhMyfmqSXX27RiJML0FgW6jaY6Pzj46ql92BYjJsXUKZGwW7
LCSu2mnALZVr28qY1Fo9qWyOnAV/9NVe8gWrMYX2th3Pl6zLHVEzF2L2NwpDdQKBjOKMLr1I73ad
0eGwceIyEQbA5IEyfhA0zFqrgjQ4yTu793P5c9nh3ffvj6/av18u3Y0ZgiJK4JoFEWSEmpcajq0R
aio0nDBHEAJqFTuWEu9qs7A0ktZITeqfdebniwOgnNtQkAUJfBBJ+D1DvDcvGOzL4ZkLaltKA1Px
AS3kgKY6W7SleT29zJrwks16703ACdOEXCfoIlowdQhMqZTS+EqrXS/wxQ8uxPR2CzEmOroCTcox
MUrW12uVam+92B/tOXIN0RACnzwXPPQrBE//JoKNWtpwOYFzvBXr0FHuKwLmuMfsnrDjCMwnG6Xh
lnwvOduANNuYRbMcqdQHh0J1pQZPA+o06wcGh8XLsKhMc2xvVbu7PqHDArfvuh3iY5ql/0z4cHdc
I9QzS2N70Nkb+FJdVvw4eUvSAlTki5OFRZWIDgRyp+NLQ85hMSLK9ZmqmualLvpEeHrU6TMRhWP+
u054B+SEdOIKnMLCdvmK0d6CtgUcF0L5tbrrpP7QP6+ZJkvsvTzwTRNHXZVTvuhzZn+e0SVTsM9r
AnpXIP02X8VG9ULr5di2lxEVOQqx2AjgE8KOGKoMpQOpD0PZmSL9REp6MsiIiUzKtiyPStpwW1Mw
vBE6jXHnxzUoq5xyaL+zGmmj65cMaIlRrCs0bFznPYh/FF7ogHDZ3GYgp5/f8ojfiJxc78nv8acL
1s1BtDyAqk5Sq28p2ouXQ3Zvil2B/FMFFAEj1144GSmnFZGFY79pmlpopk/nZ8LSw4KpE9wKtbZI
o4Ma5pYsnLz5ZynUY1vjshxBYKOZysfC/6BWRaVWfEZJQfJFgb7lNDGGM0VCuAL2AQK47Piwf8JP
sVhtPWItPVl2n2hZPBS2EDM0Fk/lIdSL/yg5Xj+8YuzYHYe410jitC6WTqbbQTKyuLZs7EPE0djZ
En6n0EZ/YdcRFyHrROPTDoA3tfmhZSJaGJyVEqKxjoOfMxf7MNCAw62rzvJdafN0WglEsQIhYXBT
IqjyOZIlbXmIWevBPWQXW1L8HX5bqqflw4KG3zstkCCMYZkLgYyPCItLtWSxWvV8w4sROG2pGWvS
Gi9Wvcdyf21JRnUkO8KP3T0C/FQKXUxCKsvNjgnvAB7t6ceyY96C00+M9edeTSjgaWfkQ5orMJ7t
HlNK1nQ7v3HtkGI8EsDe3+NUsKzgPWcHylEzcGDheBVF1orcTRGcEMpdy3bisGflkkfUFFlfDRQv
x/okQBDlLLkUgDaYYXqh0XgMIdytmBuvmoRzMl6rycRjjWpQpYCEneSZxz5MnvNJb8aj7p/uRn+E
xYifV3NZCtQKYxyBcjhToKniOHSt0hYlUGoFg5EV6T6dGyS4EB6PoTUqrzO6gqlgFCvBdGOLJuGD
qxmVR6Ccq7/1mPaF7ppkulHTbdQavesMuwHPEt35xmzI0bi9vF4FwfpqyzjPNvRbByYyuxRFDvgs
EdlwNn4wHPEebyFs+nmYqqhblNxBLNP6OE7Obw7qypAIQWTLUO5d198cyEIwWiQ29MQViCBSNYkB
iDfY385C8aYk0FbEL6wZ7+LUtAWt2i20cXj9h1WHBBxM1ARdtTqW4OYo0aEDdTO5wiAdb+EDWLk5
Nl9jW/5/pGy4IZiayL8okUU55MuY+TrDGro8qkob4WQxpU7M0wErBJ9VjN4ctH7gLwaDDEmDKt5M
UtI4UY2NyQOYP7NfmDDr/tJZyT9hj+IA3CGh3ugzVeXh1gCSzxB7WBO44c50xlGXkRq4Jtp8Jlc7
k3rW3/Ox9ui8mKw3X4W6BYg+zv+5a5mJX0WWgL6U/1HHoHwMYJgePMaW369GFaGX8kIvvF/wV3gD
86D7F0CFGMCC92Mzjg/nNgI9Y8KDjTzI0jrpoCNm4hURiGsvhnT1bLa7TBI5bRO5ko32QNkadBb9
VOkVTLrmAGPY74f3n9W2J+FgYtLnqZI2fgssaanAG7d17tSPqIcNyAFKXaXRwHkGqr1YduSwSJsG
odKjZ+eayGsGCBRlq1QPRZec27VG84A9EJi5wmHcFm1fdcq5qPGnvV8vngBry3/VZXLrK8C7RLaX
ffilCd1VfivNxgyEGmi7H6Tk/bKNSpcIxWTjKvD85yxhcuLV4cKIkfqHB8V+1lpnKB4zD5vfNgP7
DQ6U+eS9ULBX3ycVuo/dbjW6vK7fGxVKot2kw9KbUAUZF6VNN9V+8xncqTkxnSWCHgpwxdP3mg26
vR80gv4lfBYig0miMfJgqX3Y9jwWshhiaW3xvtwHF51DPyQyVF4dmGeCgHw+JCQZ5JK9Iv6JS22U
wq0rn0lr+TDx+nI3kQHnaURAbl6jduQkcIZZwXlwxsC4GtZyZkVsUzRByEFuJWXpOoURbz+HZ9gW
XG0Y/k3LCvy34AMRI/QDupuuamZKlasXEsrGOGo3g4wCmq12IyOObaFck97sZtf4M36TRSpU9Kpf
WdaZj+YPoALm3i6sIrM5N5TEMKnxthCHwAHgVPf3KLcyTSqIda6m0c910vZG+gPDxCTvZUafkBdT
99RFWOpKym/5e1ndJgsoaI/NrM5fsXcPXqK+8PxmmtjQl5DEAam0yAaZsZBYVzkSuBiZTjjduT1K
bTotcUS13EilaPuOCKqD3QKrNGgcVuk9eF99Ia3CYHObApX0li0DpIWZ3VJIwGGB0D33uqZZ8pP+
1Peu3NXGlrWUdgYt5tJL+P7FLUgkit36JARRuw5O68Ju9h53VyRcLMaZpCKAJrL2RsGGUOURS9t6
jM9EuYtTfbha+hat8No57xToeuXo72O+GEDKd7DHKrgBcxk+x9hfgAGy9kVFzLNlOzHOKAH4txlz
Y2gWyi5QLqYl7MmPfyJWcdKnIu67+O9M58WQ6o5gRz1hwPcjAwEsxFvkmHM1u29vev0fpRdEds52
gjh4Xkk5xEdRU4kOVeyXZNV248OVXEuJTnxkp5l2u9p41ZQ7qh92UujAat119F2O81Xp36LW3fcI
QHgSL4sH8RuvTw4SKvyjKcOR1Nrfy8KrvaCb5SWncQ0wyvrpA2/+EYVScQ8HDhjGq0xtSZalQIUp
qKKaNGFpxWNVP+urmq943F1ZmuLeTIdJ7qWpkhxSDIL2F0+//zHobtjS3S0sVjK/k4mJBFcRQKF0
QRQ8Ggw5xoLFYapiNGqFSO8sK8nb2cq4qRN7HZjJZuo5Wjn5o1KS3suZ7qnYiLh7wNsvl8818Y1P
tNK4Rmxr2MPTjkz2btX6JDP3hdZacCphYmk5t5N3C4sCx4Mr8GJjdscFKSXfjZiVpeQTMF9DRwqp
EkYkHuQQb0u0yULnyPyTQjyif38EqYuORFRbM1chY3tNLllrZVY+FXHcCb2vcN9x82dVldZBrcF/
RZUMHxof7VcVIBrMK6S0djMglIIFxK362oWVf5X7s62EykD4JnZQE3KBjjDbn9ZNMu/7R8A8ddbG
5woLEfTETD1a4gZvEQRfo3QD3QN3OP/Q68di9nC+gi5GRsZ/MQLRs0Wl3ndkQmVjTDW9nXZGbPD5
ATiDySVhBGRjx/XgMQ0W1Gaf6/V7QPGTwXOeN1RCr81/ZHoOVxfv8N2i5SvgmZHt4gffrpU0O5ej
fScBFlW1HU7j69A/Q8DffNrruUrtmB3OQ6jtNL6WLvfNqBHfex7feunlGD8WmwNC6lk/1+Qp1Mrh
8b9J1e6QrPZ9Ew/sgC0xn2fc0rj3IN3Sr9AVfy5CdPoD5gNKPYH9qkeZeRZ6VAMybf4U3M6qmbxF
rdBN211lc2TMtmwgZmsU0txuaxibGFq5lZaO5ET2pjkyiHzJrLLYVOGB9VmoD3w79yszbUCX+Zva
iiqtWIA8Lw8cFoLzJ8cmPaZN4RmXtaOfMgTcP8uA/snwk0svwViJXIlpjKTjsea1bBEYylgInV/N
peoKPpdgQcstezw4bbQTrRjGBpLEFXT6isO7/4WnQkeB4ELrnLMLkk9RGMB3RfSCQPerEuX+Mn5U
W1MrmAvRkYkh+9C/2YfAlRqjhms0bZTcU0yaiNo0wKCL7MyaEefc5eHhvJdy5JrD69FIm5rPleqx
jc5WgFh7jNyu5VY2mmAwC6fa0lPaFV/QTLFm+d/mv5sHKkcNPMXC9Vf4qOmlUz9AHzn45hdk0daL
EPt5g8QyehBpOzsnJ+58opp/XcFNs1W8QONGun0RHXw0s/5HAwxkvqt1tGKacGzDM3KLw7Tzj+P6
N29McHT0yLqr+G+PSTwIXRD23WQeAYLa6w7J8UMLFyCfUBd8Ed6NV3UtIu3X0mrDL7kBR/IALfdQ
Fb09QVIzJ9LA5XDjskNDz3OlL/xLxnS9S3rllVL6quiLvCT7rExGIBzlVADNgqvRJOETkWs/WuE4
4FdgzAvdP/GB/4ys695EJeNZmws016a6oeq0gJ48g7T3IfKOA8fRJUeeKAfEq6DNd7YX/DP671JM
G9UEWo5ugRh+yb7xLIqH79T1Lp2n3FH/qIeAYOZNmtTfTIBgI8n4y3AbesNV9sCHXsR2DmTz4AA2
/Zgu3bVbK4CF9LabgNcWuH/vctZe7d0a2FK+IOzv7rIbAtz2af26C+FhKTo4oO8lhmC7dds17iOH
88ARdMxPXFqGkslCbk5i1xhv61vDMNAaqH0DNaIu3lpKd3zHcNoRrP7IPo51cdXhWOwYbWSL/BFX
tfR+2UyLL7j5yR4Uv8M8jFBWLXALiK93J4cKAisfIm5eysX8mdFTYKzSInx7cGGwS2J1tpRQMYGH
DOIJ3NyATrOp0GiF7ciqWOkTrn3aV4hepqJz7nyt87I5aKPlQWt8Fg2cIdzEndNJOsdHwf4fAXn+
qx+nJWhO48ZK8+czFHWoFrkJI2V5C1Q2e+d44oH8OGJRvxmSAmMI4m1sZYZriTQRwBmHVDd4/2U5
HQbVdc4C7/V8GUQR3/wTdcMaVHfWR0HIFuEhP+83K0qQeR/z2CNpLWz0WruA69LZHzJERJ8ANP6j
//Ic7U4c1zWm0synztyMwAHLCjmFguaOLLuX/cATCS+yKypkUZcClpmz/LEErnnFm2Y81JsALOm2
0GmZ19m3x+O5GIWsTub25vI1WV1M+6PJNbZavTdbXapqybYJnTmd36gwD/3olDzKJw0QGiUdIWCZ
OCKM9UKFmbsRLaF6dUhe5Q+XLTN1oxtTaJrMpI3gqxeQSc+5uhIIARsGEDJ28fR6ewIbNtsCxxS3
QTHsoehEfMxSftqeiI/qeIHlRduAeL4nMRcfL6eKkl4kea0a7iFHcOqujW3bWvBFqMpRpJ+BH7W1
ZrzKoXmzGp90HSA9IjTIz05y4TNaOF5BHnPrnoABg7KXWpAvVYOOWUIR+/tFFE2TpzbkCm9H6Sk/
nSNGZRO4I4/IZUHy3Ar71JihnTEWEy+gbewC1xO+WhUSN+bGarG4Pmzvdm0/NTooy9HOBa4ieplM
LeVnZT4yS++PBFAL8cetnSQYmImcWVHsztXHss9QrzWiXkm2kL7asjLDcLNkjk9JAHQ0eNm55zz0
CMWTRIvfZStwArsZp6ULwpK+Vb1n1Fvdu3xpwedb0hUgH1LZE1iiX5Ww3VNWd4L8uMppUaj1znt/
5WxF2SrkwY0iJa57PJuLGw7fo0o027hf6HkPiTH+bP+/mryFLOsKSWZpanQAWkHWtVf549aU7r0w
8EuyZu1MDFyWB+nEyvnWUr1bdhp+9n6bulJ9sqICLKW2sdf2LAIJmxT7o5maw3g0Xnb+sk5LMRsL
UQC9CXUcXCydeZ0SqKNu/Ilv/RYe2QxgmyxPfe6daXsNXMFWSIOCza5YWErtk5HGuQenLtwHRsvS
OwqiCyIj+jMxV5ysqBHGPpxaNN1o+8dgt6qFRTqCIGIihDmYIKFn9Qo4MrD1RbUikMjNZyxDiYZ9
lJ3BkonODsjMrJv/lhVNGhI6wlMfX4YEmXFSmboIEJEvWPPiWFxrfjAb/rOXjY7IFpQa1V0H+3WE
rwYKzZCV2jLokysaIdwF3TZFKrH/uVPqyFGrZ9H3+pa6nnamnqOZs3SLA95XjpDVbUWkV3zmXR0Q
lWC0EpUzhxztvhxPyM9WqYDuXtqnQvFhNR4NbChTZnhrMB8BUGj3id02Dcl6frkZ4BVHTyxJhYoI
oWgxLKuwirAKuvlQXLKf5DAp5xxKh2PR3fmDy4BXiuXCxW0pM5t8ZYpixNI+x7qOgO6fBuVdrKkV
/TEClfF0xHxWN2QF6wJPJFrMufhNHZwRGhdZugA+qImyVJtqDwlkzMNwbQN3GwvFT14aJgCrxZU9
nYRJiL3Emtwrjpy+vz/bHC3m+qmz1hzWF6pa4GrMwP54B+3ipPHw6luuPGbrfxjG7opNn3wPey/a
SoIwYCs2rFa/ib87g/f4icrHbCpxYKUTWx0e4MIeIzw88ea0H6aDuuM2YvWfUvFXVoDZGgeY/Gi6
Qkokro9VN4TMuJRn9Isg8cQmtKZCGIj6UB2zb3piKD9yktYpMpn6QmJrFztyoIYaLrwpiaI16/7B
Q4rWsZqaEYAtUueR1U+LPBRUX0YIJGT5jjm2kBsrwrsfgFqR1U+f53ByNxgLIHsvTXQtQyfUyXwE
rsNWwqspv8w92+jqNYxpIcvYqvWlc4Mvyqb8rzRlwIQJ1pKb0uvyWZwQt3KPyhwyBMY5stPFZSFR
JSkRDBuBf1dmyuh23pyUhA8m61LJ8jucitSH7xY1AIY1C+Ei8UYiXn72r84bkGVRz4KGHUj+Vy2f
CUtCJieoM83NP4lcZZ8S6eJfjFlblhfm9rTzdjkH5won2WghLTx4lsxjQ/dYiJuizgT3tqIeB0SP
LJ3cO0OabZ2piza4CGJ+HpgF4Y457gxImfEm0PuQ0naVE+L519sv81L+dK9GVgmUz4WJKN8elmNX
vDW/dyC+nhZQlSkssSi+3y9MADKK8RrbfKnZQZzbPWoV+bO51XUGdMmIyApI1xG46yukbKBG/aIN
/2u7X7qZIHyrvuRvkTF3TUXzMM7ZnZ+QaqBCRQIIwIc1uVy81ckwcpFQskHIFGY4wm4meTg3NBKv
8B2EstgrweRhuT0H2eMx0JCdoCcHh5dcXmHKM4aGpvz2m6nwQ7YPedLINpR8Ihk9AJb/UCx1vY85
pNZ6hSKGTxEd0/WvlyQL56FE3wqtzi2/06YiO3QD8/HdM9+Z3ttk1qqeDn8137jDamElw/WMqxe3
LVdglERt0d5hCjV2DJ9JO9l1nDC36DCXvasAoFxyZZYr+nerdXMQL4/ny8j44L7AdkvA8OUOcFWJ
bv3qmHK8T900B7EMWjk8WiTigjKS6Bh1nGvJj7w+i7Jt12TyMfAWLKAL7LqEUnnfK60YJzuRizJT
AwT+axzVda9vFTyVtIbG/iOmBLJFj6y5wE1sOCt7WMp6qmkqzzY3Z2HdbtnYDJNkfnoBHDi6PXEF
zJ/FAMCAu4qN2t8X/LDhe3Fn/0ImB7NaXcnk7d2exJd4o3ZqD8V11Z1zy5Ba9uDCN0Z/Me870e06
XBndoo2r2x22vIZmeFueKIMIzS1HjQlXCu3zte0e0NST3c8BfcpC7JBwZ0dSuGqdyTA+C2zNtW0Z
e0pqTonsN0STQZINkbg8roP06/FTpf8ZOruX3ViJEEm+vKvIezqvRV+Q1UXhH5wNnqh6tMyjyGuT
0vJiRg6/mIF0DKKMarci/YRl2Aq5uRzweTfpFXCNUUOJgN1xjnpg4YV6+blPgKD+Ls8dF/LBupnR
hIT+x47rxFkzDddwjukXMg9QTfKO38xUsilXZqBPFAoTEQtJX6YAoUTROnxsSHhXRJyfeh4lrnRb
cuEMhZY7S3NdkVUXCnhQqt0OsbY9Ag6kzZDEaAm3oV+02BPBdpsNPEhIiPARufnB9rw3ijfIdq+i
E3QzB0thd8+6k4G7iEV48UPdAZdCtntJDkVobnSE2n5o6RwJvc5vnmvQ7ZrS6JRXZ6G1MFzop/fF
mCE8gF/yabokG3UbJ9MTF9GAeMPMg+k5/BtI0JHlqrJmHW6IaXcB9TpOfYnYpj3ppVAltP4voKGb
EK6sG1HEzM1MtX55cXV2Lx9RVlbfs0MEvZ1+k4LBfqw59zBikfp7kqA9N/oFesMrXi83l0XqVp/x
DZhqKNXWFfu2cVl9kz9+VuZkuiwOsSeoewz0hoQNf1SKH4gkmyBlyHxmkBteVdtYRqFkW6ssB39m
qbpmb6xi8PiVS4mIBgNCC/S+BWo5SRUrIZmUN4NiEnez4PnjYgYQn+YKIfesLt1b15fnB+23U7pJ
oOPW4MXfVmcXblPLbKljR7Pp+xQs05+WHRPDpUnhN7fyGuHgTh+iqoXWCdBy/tasaocF6dqg06Q3
8Xdrr6lRL83NiNYZtaJ0O496wsvf4sRrlq7QKRQN3/P0YSkq0HDwlUr28lZgq/GAZEd4vpMlcxwK
45d2bAiktTxfVpxEfqt2VUu9FYkIK52iWqhrbYwlt5TDZ7qE6WwMRFh+5Tc7w6EtleYTmZJR6fOW
5zGK50OrJhsnJdxyh3PmEEdJYbXkkol3FtB1J6hqhRsU7OSTRRAn/NkQ3Bmko/fcCcwMM2Fs+gll
wcKY1/hzgMEiBR0Eq0oY9wkqJjmY47cwLu0jlhgGox1im59c22MMkrRCnN69wu1OGLmTzCHeyg1v
q7n25tOJdn8ppaA/e5Wl8K38f1EXAwLurQlfR4WDJ+4F+MRM4OM5M5A/SZjNMSS6IwJkBFUwAQza
o2cqRlXZUmu9gltE+RNX+HLVj3j8ozMMx431o4e7pdRlhcv0qHKKcwZFoXmrvnc21rqBRm6hl2/a
bSXFtQdET0KrUQGH71wlyKuGIYih4ABm+Nwcwy5RPvij4lHfc3UjqCprw4haCuPQuRxIAf9Tt1/e
HZrNSDqlIZ80lciNvdkiVwNo9jNKZ6rG0DVcmspL7/Ly5JoN+k4obnDbUkHkIFgkEfs/tn9CUEI6
UEA+JZXeu2nhwZamNeCvpB6IucGeu4o4Ysq/gB+oewhErGGChIw9mTgwtstj8vJNV8Y6QtIFpA+c
2FgHYHg2tfatfLZW/sd1O1qvLC5S7ZFZiOBDaWxNH9g2qherKmsp4R8zLjbEdnp7RSvqaoXyvG/H
w9qTEGkUWKTKP4UTri2awQPWkHOSdVT/04riREU4QKzA3Wh8SRiLJTfS6lGMe0WefNDcHNrargVq
7ZT/lIx/yw9kzMb2JRxpBxc/Ro0LlK7Yi1ZnZfFQUendSAee2WHuDPXG/+bac6K/A9HkMkfjGeKk
mnJonR/R/idN/rWxX1gQ7nP/a/GqnoNcaD4WPliTRPWqSsD0q1MZ5t3OIjJBu8q5ZfWHAk4pNj78
qXCJyegGWrBcdoV5MTNFNbETEkD+YEUDeEYqkKDGA+1mQnIJDmO3lMannWe5+oTfYYfbFMLUjYkn
v3vfMfMyvRDL0N312W2+371AAqwDVLcImDT6okyCEYjHOHARvi4ijs1U51n6gA1IWIU/dLT0CyK0
m0EyKUtsUyR2I9LAiyQ1qmof641k/9XWlX6fqetFvdC55FdaDtUIMyIYNuvtqyF0ShUqTVil8InP
+mvZo7JLvjF2UWy5NFIsEE+JLj4ZZW2fqp+NXhNQCS5v6q1d3MfXN88NLLRMuhplQtktQXWxN21Q
Fl1/7Nhi6wnbfYcbgzZbBiSYQCmKSiMq0TzZwqbozIeM6eQ3UMfyWqRAcKCpXkOSXh2wRyBNYNFG
bXstKeyiQWgXJ4x9h0pWdSzAhda5m4nV0CNPQ9IfGyhD393fWg36hQvPV3Xx4N6yZuVds7WxmSPQ
VuGj1nrr4iUrjvP7MnrOQ/DROYGhBjFoQMSVQsJpp4Jbc/46xq+B5/crZe8nbpjHr8Z2tAQ+fFMf
/n1/pSqakw+5odKti3T+M3Z1Y0nepNmXNF/bSt65rzmFIKORebfrqZOlVJnyOhfA8cC1HJgzX6hF
xqYXZXsUvoLCTdA112cHHeBoFthROtJQM22xAp0BPis4MDK47gz8b/Le5y+Cx8YblOxLI+XdOr5U
OLDGJVTkVD974eh+ZgCBjAOMNc6c/pvo6ayUqqS2BD2aXHCK9S7zlL/WUAHT4J/0sLzvPOyVWFIa
IUPQlkXunplD97mve0Lsv6gryDR2C3VLj8lLoyoWnhXDoEOcpSjEYNJ3UOVdfB3JAAExhWUp6cY5
RwTPinMyERWfz1ziyGN8Q/bMHyRMT/6mdt8+JDL2GVv6uEgAELgrSjSbH2GS+piLo1UmLZqSNy3r
0G1GUSSgtij2FZjY1cxdh8tglGODDrgTPyENnTGxBUFBp3rVPdHcDAxPd/pdaDkWEHk65PT5aKi4
eftCpK62EdsjY7AzK6PNAOG+H9Pw4CghIGvPu6/OHZAKohNS2CPP85MCiBMHoEDga6tC1G2O4sJz
EOghXpykrOFmcxOckJHSmrC/e0kZBETwCeWq1d228CvGQkV+XsDDYMedkQPWlfGDcTsplw0a+S1G
WiKL2zG7xqwiJe1OM5g/AYk8fxFCR4kW1iDjoha4OTIIG+kJXQ0gLwZnDdWmx2djtu81/AAonSZp
6wc81GExD+pE+hcNHuBMW74n9789VilEfxU9Ls4E3cby7Llv182gXvohVIFcbv25PWniNSP6Urq8
Thxyz/s/Sh+llE3Ph3q5uWAY/krXVGjQnXtwhUKfC0oA2ACUiMcbItrxKU4BcwgVm972eK6J/0H3
HrsEdLD86mJ33+4Nd2QNqLq9Zti9jlPawUN2wKfyjGeYaC0MeLN0M2onkp2t0UNhstxzDkTn4IAQ
IWSiNTWT98R6HBau0DiuelBOI4yRjWvq0np6DFJ5yMEW2tvND9rqHrwE8V7KgMELnCt+N72YYgFY
7RYeV3FTp1CJ/+6i2zaKGORArYoIk0YUgd79cmB7bi5JyMv8yqVRxRzoUATy2LgANTZ/I8Q8dRiH
LTxEHSBKHuUV1Jq2bDEEENmkRkcKubt4GAnqksS8LtXKU01enYehgxmJpdcgb2mckAGHm+WTMBGn
4Ztt33KdntORdYo7DdjYQ1u0pYcd35nwuhvxKDjwgRKXX7FqoM9xJW1IRaX6C0hF9gEsDgwVnrOI
KdJXnDznn4kd1q0UMNyp1ZqpiOFriTsBn0NOMdls1bw4Tf3tigc6PgxdDet0gQL8jj5LvHZRumeS
wkH7fwpdRlcojIn30n2j+ehamAMcn5EBnHfMw8xHH/mEsWinR9cTID9s356IF//o9LhG9njbxYIU
vfSaUfjLjjBw6d7EdMq6tEkJtZjLRE6NXpqbmSUHsgC4Jed+TsZw8uvHqXNtOACVJixnj6B9FOI9
WHSElBxhqrqA18nroTcWnDo0lHwILTPfGhbQnSo+mHgj28mzavLDHeCa+g3XSnmBLJn2CK25pSbs
htWGwCpJh59xYxTwyOmt2LmBc/Sz/dfRy0x2T9iHgXTbAMGSVzbCIRJ48VRFtKEQqJ/lypyvJtcR
N8aKTVeY6vVKsjLEboPZjwfLFW42ijQDhWhyNhSYYf0ydfd3/YQI8qcW8LsTpLY0DBK0LkDRTx1/
EyYyp1vjvQkVgjwVUzTEERBwKDSk1Z5lOwiTdTriHF3pPOFFcb3fVeac2gj3Paiz9oYDSKzE+8yY
5OnVZAePLWFopt0sptbHR53M9UY/rbhb2kLOsBsIfqtAvuToMSKnHr3pcZWIh7TEQ6T4O4wul31Q
3vcB3RH2NX8hlFeqmX30yOQo2fGNB0lmtLByvmYXP9o5kANdWdNBH6K+iH2NV+nlFdFAxLDXBeON
5y5i/j6hbffY+aOQqhcHyKAgdQIf7FkgjRV7Z2Z+Vb+ANoOhIyrJZnxQwOvrOz/VaLUKowyF23q6
kqZYUO4LuJ1NIWcIZOqB9O9hJDToMLp0Cq2KMaHr7MtsB117syU97+EZ8DBKeSIn6dPD44J/y2Li
GFAVe3o/uorEBa4XuSaH+ILzEUpaZ8Ep8eNvK0Qi2pQ90VdDKhEek9A9JdxD4g1RKqz+Rff3pQXL
fykBzrsADUk+9CDyzw1q+ddkdS3kQTblAcREyUEbBoUKk4oK0gypPeHht/GZoyBuarkG5uQyauib
nCARB0XrSagFwSPiR0ez/2SqlCSPfoCP6T1AVjFnyiM8gwfWcYnSqTF6a2HMh3ZFpIBqlgj5QqHg
1YFXZ6vk/fifjI3rpBrabdeG6dmr2I1+lD7tlA9CxHK+XR/xvvzsBLMG71Qz4tpx40DW+/u5f1K9
4IfYIZqWadLpk9rNkiaHlltamVAJ5RFbfPNvbEKWe8ixsii19tRqIJwMcaUcKHUfbmfAUgGjAqxl
dj/IOaJmvXfn7KtS2wf5zto9YJC1lwW3X5s1laPRzvMaItmi6Ur7JJccdEiCWu25ypJpptuuTNyY
TJMy+Kfoz241PyYaF7xwlxfXNmM5bAPF75kjU4QpbRjutzS1wopQgJeC4h6Xxscf+qkjuNHq+VK4
TqJjpg85IOBrO+jIfD9l4G6SLYKjLWyASXdQkRh5MHntDTb1a34UP5QXyOje+mncfKAazhIgbX8y
97ol6moOwmYGDSzi57xWD6R0iPz0Gr9kBjnMmEedVoVfugsc0XZXDc/7I96kgsQpjoX06aYxedvO
BN3MZWfUVHe1/gLN7J6mjRB3QCLG8fnkU8Kv5vZrYlkpaCLA3UqcijgFZcoScXdEpAE93K0iElCb
q0bSzoaGFYn/ezv9IJDLdAAorZVPVaT4NoW2PUWnC0IkFJL+44LkA0pnCuABheRgFrWU8z5Gn+TZ
J44mVQWxisMd+s5AV60xWwZo8bal3LmWl0kHNdHq0m2HcuiIoctQ6FXNWNrttI67ZZccy8LvAY+b
TL/+qgP6u3nuYSNlGn+/mucZ2mAiOHpNLawiBpTTWENJw4jJe91Sz2N746RRFn5/lJTkbvlSI5YF
60bWlbz3MEixCZhtajUrnzkkOPhn0apkya8oZaJBuYz0+RDX18XKzg8E6xRC0FxCEi8OZGJyy1uK
LYaHvlJ39SEm0/STgpxlN/WQng5ZHnzLJyqTcO4je6QBf/4wfDYRLPjTMf5d20owFO/9/YmG1ZS3
5vmNd5oWkTHo6I6020dHya6atYkvCUuXUCrVcPt402sgPLURuGX/qZvNkD3+G4WluKikrRSE3gHP
IGZElm/CtTNGy1W4XIgnY1Wvr+Q75LMVcDvFK2E9Eawu74z76HXGAtQVlylmQPUb99yNc9bAn3Tk
1da+Y0TrVUd9Fho+KuxCWZxL0EUu0Vibk702BOeBiTdMoUeWEFEylScHCNBZSdNpcbi821hU8Kga
eQQRJiP7NuCQWqQiJG2NRHWtE3KVtIg/ODQ0n5nsTDmBe5n3dYK7ZMBoAQAf3xORl+xVtlkwXif1
Q5n8k1VmRNT5RpSrVJ2Rau+SLH6oRngfXQ7xeFvIYpFD4yW8Z8LG9waf21aIGxA8iMyIx0nC7vC5
/F72dSfTAhZIfQJiopjSzUbMmLN4O385HwB/4EQQ69r1NbB+Q7AmbzmWFsDUYLA5pPMEWGTUo6tG
ivne+HgLN1wwglVvVKeVnJkMtnHkYUcNnlN2GGTS+cwxkNXi4mBMAiy96jYht2fCKajIqxzc8HPj
vR6FyH3DT2tg8B1HYuxYem0nJdUVhGb0ACgqf8NWe+FdXkuQSD9WVRL+ahAKGVEi3/6b7urYIhbm
rZ+pez2L8Oi2DF27K1MxGI2giEGuxhpqjkhukgerccCeZAEcjsCHCusKySI+8MpP7+bY861DDNDq
h97P3fQ9oGpQLyYWJQmomV3+JYbX1C/xSOaRsDYgJ+ZfWV38NLAA/H4k1sFPrnEJ3WI4UXlMg78r
XNEKJUyfyUmscDfxlbgwIkx2I8e5Wab93UbAtA6fgBzYt3FyN2Cq9ekHcqTFp/0KzhDDINogPPjE
8SAnXmc5P4/JNyammAfXXDuTIfKZnDZYO76zJEfzZEg9VrgjykDmhpSKgdqzFlwswjdDFy0SatqF
ujHbz9TD/QnFCdZqISNAy65twQ0ygGh6wXegY/jBBnhXW5WG55Tcp2BDuGFmicZ5g2CQmpDsSrov
hZB9sINjk3r4vl8d87iw99Zb7I6YH7As1fqkRoxfcUXf3q7+ZRAKpjKJ/GbLFGZ4yvSqmAa95Bmu
v9H2jkmzCJzgaT1nezrhvR/IQvhwoWYUUV8YKKfRNyLvJ0+BCh/QtshpMHRTYCJovReDqColm7oe
l7lXX/Q7AP3genb05ZD/n42/lts4nZAqiNpUVY87LNpoJRDL24QcGTs6ZhvKfBydTQ6LGuBF4/Iq
KBEEAC8CyJp8Y7Wv742KKsFzWQnpASM4frkgZ64amG8+1VEY6/+SwY91KZevbiQlnPpLUdoVLYgs
xLcTtWxxKi0bLP0lteA0HOsOe5ys1pNj/j68BQzbQmPKZVL6ayJsqgNI82YSMzcWToznsEEPfTWZ
1POwthEKIJmUN1iJdEopUSxMvIxEdVF8EaR8RR1HzoZLHjNR4JwTwL36m933T0nfdwtwrCXLCzaH
bR7yGhGna7JFMx39pxI0uDgo3Mi0HgJ5QZItozCQpYmnTvAS2ED/UYbBd3+pWLBPrmGOdMiZIkmx
mvDPQ7W3gAZwbVO+7evpZ2BsiwU8maHIybOrJbwLMIVzuB7ZHsr/bFGp83y5oRLwQ+k+q7tncm2o
ugc5pzu8Ns2oh23tUeh5mhjavWBEDBQ+9cSnWWnCnVYe2Ihwes6DnwUZqifu9APTU3IY+YM0Z58X
2UmLKMlwOrIMU5YGgcYyNuQJ8M0Wb/rCum8loKy/7EWSkWdH4/veyirYV6KuIU/wNHOBxU1fUTun
XpX7/DERLhDa1qGIKCE1vXV9IWwRP19j8yutRQ9NSxYmzJcNPK9MDDpa4qWgWxeD14zzN1dXgteF
waMO8qw9ymse+ELpEAJ0E7LPqOQsYuhjI7wga7N/5pE/awCEsmStCRgNYbHZ/CyYs2HjVjLDTuFi
27XsX53uxwi1XKfjGiOjjkXa/KjAtaBkXnXtjlZG+DtqP8+FlRiwq+SFd3d2fDvjnrLY3bQIYtKp
SZ8iBySgSSOszqB8NWLMAep9XCbmFfIGAghlIVkuy84KAqgrBSWG2nGnTcAZjT1TK81VMcwVJfS/
ivBnXdKbWnmJ79juE4TjKEyfXo67mcewrqKir9tH9U4vvRRfbYLD3XLES0Gl2QYokldtZg021sf0
pdp+7NR+/1G4E1/bWe0/l+6TE0YGDmA5G2uXNSwp9JlI4fbFtMIu7aCDMXhucvqwP9sIZd6o1Kfx
CntCMWnjcw0QcubdrzblBuRFu5TTJ7I3g8mrSSG437/SK0pbxTeKMMcQa6Y60RCz6On6N8JvpLwS
hJ3mWH/Tbbh84aG1K90YgMDMZPHd6eSPCwwywLDWeiXJVNAx8htBAE+ZEkUyPpesNLB5+1HvbrS/
rNBczN4ye6Qumz1kAwiewVcWL4uVmcr06S/7+/j4UPLuMBU9mMafT73rQoR9d3uvNgpZf2vfdjSe
jCcF7Rh3XuIyVurhwdKIMKrdJVHdAFQCOXt+zn9SoGINZQipuHwGgc9ndpWLsDdi+KBpVyLnUzMS
MGRaAvCfqQ+NP1zfRQP8q9uClnfU0jlhQyBKKn7mT+Oq1Aawy6DmcX8nM/XrWoNi6pZq+4p+eB7X
urhkaS23O/Dmvvy5X7hwaucjT5dmDW1zmquTXdlNKfKud5DUhLydexr+XBbVR+MH8sqO9g5UUsBR
vr0lpgs/RdbwPC73UB90bjZFDNysaR6l1Y2vmw/wW6cHg9mMn/hBPIKBWd0vEy+BrPtSXJF9QDX4
i45yOE/t6ym93URY5ckE3jizkfja/M07IbQu5lTPMKZjO+q/zoJaO/z0WSL7Sw3KJhMsQPbPVEXq
C4N7btYPg84nP8Yl9TpPNlp3LCMzdpTE6TyJXaQ3V5oJI0JVVKqkDNp3mO2qHFlVNLkLdD2ZX2Uk
u8dtIpcJ/+sdVZ0qdNy7cPftlpvq0hpuXJqy989WZtXbB91DR+rJL1po5DAj6readlbfT49dL5wJ
4uRyjcX6i+klglphRfrKujRvSoY5Xq2e1L0Olojj2+8ZhjEA/7hblqwOFwy91+osu4aKzvJS9nzl
oCSjBAGtMawkkfCm3OzrMLlDiMJcbO3yLfROkJnniG0VW0ATeuiQPymaaNw0YLLnkhysUpaIf4aF
Brd6TwnKanb1wsLFrpo7NmLS+v98yCUnXbTQHDFb/D8j7Qk+oonPtvzcwRSLBgMlkMtawHcfmYNC
TQvHt0A4oIWf8gVqJn4kc/H2B+/wDesJRbKt07oMXmzBNwnS+qgTbtf4FRY9TANaPwluFIqZlkdh
AUoXirf+QyFwxorDjwVXSnDD8ai67EHHyJzvD1hKA7ju/LFESTz1W0AQef5BxwoahSs5zM0FpiVZ
zkh1k+mPxBrGoql3YnQT9FbWoTMgkiW5i3R8Duszak0h3nPfMxEK8maluxClwPi03doYozsbjtw7
o7XfxNLRDx88K4TK0TpztWObEIn9TO4On14kpEz5peGRkDrbbpE/arsTfVlI1RnskQc/yIGh6xjT
5t5hDY/l3w58OxhEZkMva3nsdZYcV296ZbjxRzKX7ucrNowOPq6q1aKAulDBboFdtrdf6g9uIQWm
zDb0P3SJDkk2RW2dlP3qwKVPWpaehhDbb8ws71aHwSp84rH9qwj3IbqoiCLM/jpvpn6aZCjcMgR+
9n6VG9QmzT49rNKlai6PGVFjRqHdvZUeliqaNfEtUg0mQzTFZPqbTb/jHeXZREMTs4KCp+/1Kkr3
sOfrovcZ5OBLVYw1j2fpjdPUanRxe/updou63XADu0R3SgxSaRchXze9CvcMRlods5aKjoHeRZ+g
ypqfGQOvcmC2aebV9Wbp5hmYxvFwsdgsIlBMfdkyeL6d9H2NBelDALr5dzbVb9UR6vsqATswLzz5
FdLIn0TC87BugZ08E2xngAeYjYVFnKeS2KyKJifaKYw5eM/hWBjOaMlcmCqMjsQxsdOLDiiflaQB
GifEis2ZH3OCiDo810GboHqWJsm3RJWc43pN3eBvjF3HhTOpaImXNRtA61BhLM61WpCeYC3tiQuv
NzdtGqzd9khCa0jJ7Yb1fUPhWG7hvmVgtXyWNviNQsnl7a0BM1MjLElniHFIuk1vU91MLZispg8U
dpLzSy6R/fOYFsnNWRwZOdV9k/vJV7SU2xogWi5gViizrC7sw3iwBfpIWRDY//zptiv0B7ZT6pUf
tBBTL+xAeLk9ULui2ooO8P54ApvGlfomQrnMe9z27z5Z1u202jTfx2i35tyM2KwK4R2OLGOZjff2
E4HlbR+SkUch/3sEPYq5coNlDLNOhsa0eu5ktezfxXXWFvWMM4yBEeBuXxvGps4UuEAlw27I8dBc
Zd1Hq8Qq3SORgV/3J2AbnBT715J9Bg1NCuTZ02ri1IrL48+qFRQtQmqlSWu7OEkCPP2vsx38H1sZ
DFTiJ9D3VV6dypzke3rtIAOfR/WCjxRnR4DcdGG93S25B/7M686cdH/WBiEQ3duSGwRL6tzF1+Qd
TpwecdFKcscBdVuBTZuoRTfKju2z9dhNWTLpO/T21w73cKWXVbvffdw1/3mlPkJmRTNsbDav0K4P
sbLcRiDfo2tKdVvKoM4JvyUl1IQmoPKqFZbktkpNVVFZ+TKF1QiTWfDOc83etXKs7Ts0Fht55pvv
YC5abzbzCuR0hMhpAZ7NGXjD3qf70yVsaaLrjqughJx+HF1kO8kpfFPmlZAfMJ0k9vhq4JCTEmbq
k3xmpHF5zTjQrQ8xl9nVISuihFLtlNYETK+hVa1xb4dWNLDuGuDqOU9qXAp8CVSpn6hsnjQVRrl7
cdxeZ1HT0LJTyt+CV5PSL9H7tooY1DGg/K10kTaa6WvtIpOFqsZJ8QnnhmZmNAaylyMnQ0cr+hzE
4pvNrseHQfCMdvswMwpCJc5jHRjoOy8iI7ZwnBRJm9UZptcrmmobrJCHsSlwDGfSXiRPTd2ozt7i
PWgtwh0jw5k/Ouqvzh7YHn281JatS0irfkSkjke5OHynGjW0Ab88tsSJqbs2mOybRLz0XRbAHRUr
LbJloiYW7qAmGDNDqj+lND/FWySOGaa1pQKRwyGWinL8ce5pLM+P0HWM8cqMHRPm3+AoCeaPX1B9
MxfV1C34DGmhomzdzoz/VDzMl+1cstxovVm/ViDnE8N1l8WuOsitesMZtfBlR/gddvOItWu9XFDN
XNsyWRCL8XYzFOChGrPPELblplchIKl0zPVv/1UK3pYXUj2XMJltv0MmXaGRyLCAIKYeq16u5ReO
PE3ucreS5aW7d7qC6kjYmZT7P+qahJFvaDAKPCNBLhbAdE6h1pFbYcZw0xdo90EdXt1w3iHM+knu
MX8Qw3PdhN6csaE3sfWuKmnEiQcC3LpFDUL2zGjN/NW7QD/qfdDN1R6aGIitshHHkGUcrL2zM0n7
0dC/fuizcg7fcwEEsucvo0O9kkSih04hGzgk5VTqQ/WL3scg2+TprY/+eTi91t6W/A6/9H+DCSoa
tikUEPGZjOJy5VKYDJb9k3r2ngJ5XEGMJOmsIIcRGPUkuyPZih/YbA9w120Ps3BuWv9/pZZf3R/D
wM3WdKPgXx+wtmDzDBC3pQJYEHdWDo2tz5HD0PmIAwmJrkJEfIq02dC9KPkerfKqy2HghfX5RluX
tD7+NqpEA5VQUgrI5o158CcR7u06sUnvnl9lTQoKaDg3p+IKQLYEk08beJCRG5WPEJ3bLg+1BxyM
seXzcxMLiLyws01aMRwAJa6+LrXJ6mdcN3SobqHfzpdLTTfaulCU2TCSX9ESQxBoLCPHllskEb2d
NFEsy3eugLADlnwf5K/QkNWerP2kFGaI66TEqmT1IXlakH4eBHYKpL4ZBakeQjQwdwmcPb6VnEZY
DgfgujQIkezap6qcSqOzWO+r2l8l3vhqhe3wgkzeXrxr8r0j4Hxma5tGGuadv6u/dQxahJuLylNz
400fgC3PW+nPCLM4TlcfaVDTmGY/zOkypnOjF4xUBOXe/hU41nBZHZvFqOXIOH/9IKvb17MC8yGw
/SA37qjtXEdLDgPUKuu6E1iUQ/BoD+5+PGrqhhjIp+A+pSnybNvlNkD0uR3vlCFsmzg4lN5xI/iI
HSXqU0CAElqN+KozKNLuCZukgshg5rBLHdQYFuSxoQt12I9thnqNeQFrXNeb4wEwMBc5GAAK1sdh
mH6DxW6CBBXVzKUapxtJkfEs09GMh9r/9E5RnL0HMYzjbxRNTNhwyNkp9xaTKCvAe47tkwdTDsDN
TzXzpOutwj+527h2Xg5xDBYOKp19mscaSQSulVGeFIbRyhy2bTIEtDDAt/B9idKeGyU+sN7fEVOR
rrt4n27E2Umgmg6CnfuvrgYN70AJbCja7wrV4pH+nK2zlfi5P1YNr1N56M5qfq+kOGFkYf4SFdsk
oRr4QGovqwovwppaXf7QZ8KbwaG7vQf75OIrW3DjDZreLRX8RAlIe5ADKm6uG9LpOjL4qunq1OW3
qELNcwaz6SzOFVPfd9mEYLiMPI7705gWsxSFRT85Sdfix9YBSYyxoPCMKVAETHY04a7r7z8Zttij
rt7+8V2q8fd+oeST4W6wEaF+jSvi5NW/GLIN+yydkQXdRU4SXCOp+ZmwqzZT69m/SrcZLHvo/E3G
MC7ROFdGeWzovh3mgFNIqQCmsC8bKkDX5PiLDty9bNku1aCSNxkPHas+Wdcn8fWP9EHeeyJ9iv1R
euKMXC59691xLr+PRhTnw1K8lgd08Zew8T/SP6AAS7EKWXB/REmP3BrgOwdnBhozaac9TYeE/dkn
XceCJgpRViUM97LzgEEzuugzvDKFR4bdIa+gIL+S6yNhSJMF/azcHOwyT08eYaGTZAWMz9hoOzac
RDGlTqtviJDFX61ZJVFQkNCG87y4Ta8I1Fjx1pANLDtjsEvzUfsAkyudglJhwOYdCmamI62xdn2Q
4TyzP4857P8HfCJg4L4/A6WcCaVgLpNONC9FTzugNLGxL7NtUfGLQMi61wIrZY1LK/+JmW128QtH
BKwYcmuwn0MUFQYJSjOVUei6fCOxAGO3pEU492j90G/EyudEjrFLRzjmBzvKJCcCpi39OgFLrtNa
X4akZCqYq/V2DCfHOnT/DsumouVYtJGvYZsoPL9IQrelFfUTsBW/TZzmndUFZjXMAVC6gHeV3GK9
/YiqtiqyCvolPzU+5tBOtXsxbPglgjtwT77ghZfdfNjtRaajcV2JFSod3hx3BK9UOoBZDrg5WpTn
bWDt8seHU9gWjZYxXs6b3RCkS127I70KZS+vP0RFMuAMxsqxCFCaVJ09umt3gQwbU4cgF/GkycRh
/21TGcx9JJ1iuLvB+Olm9jGRzllxtbRcHKZfHV1agwj8f/xTytA7AmWAmTVwbb5/xO4+t4ohwOko
GIBWWjysg+7XYkmnorUgMzCpy9hFLOIq8QSEex6dCbr2chcFNAd7Izz3c1vCMXB8QZJh3zNDdAXH
BYTN33/7nJ2/bpKx5HGlDVXVmX0E/jx2oJ+xkz5xLlvluSJUiIt6kuY/ytODYruz8lVmjgxPWu/U
gk81JRjG06VWpaCNMJAnVPTPMunAbiSVmi1Od05E4d78gDbsRGFaUldAz8nVnDqlxN1YHdQOLER5
PueNDowhoMG+6RjI7fM/vMIxDI7jUP9HZpkYTq9EtMbGiwP207VKalQL6eirCMm8kzq4YTfYIPJt
GovkS/AtwPJix/2DVUZTcQENqmIcWVMlx/fqPAsNz8vFqvpNymCorKWG10XBGLSaf5Y5/eaBDq+d
4mkd8ki0gK2C+pbH64MJo7iExBHVpnDnV2aedmmya3pk+bnUlhpcB10YDv6b7qOOUuonRO2tDsVX
xoBN3oq5rjj6YstR7sLjJNrd07c2VgWTwjtZu/yVkOWqZq26GzOpWPSo39qrTDF3ZVdpbt2Rl2vV
DZ5EsDcgg9e7UKDI1peAt26cO7CKe8hAvYrUgo7N499xxWiwRWVW4k0M65tFsngFNo0INLNo2edx
H9LwexHfm4+pzZaG6unw7zBHs6p5bHOGHl99T6FLVWx/Ow3JTWjzBUmLuzu0gkFeVyBCfHLJ9BmR
uB+CzKwKLw1igB4ck2NPB3QXfpsz2eC9b/gotXmsCSakCYplnY8k+zV6kFRs1GYzAAVoJ/LJEpk/
l/srHTfPo5ymPOU6SYDFAElQB2z3vIqAuYitKwmQziifAcEGb6oJKiQNbmI9SkNVeExar+43PxnE
BTpd8M6R5i8OrfrOb8Kw8QBOhIdySONbJ7bg230EiVSgkckNFsD3FWOP8kXYPkp3jXffbCVtAiPP
9bq/XnLaNAeyCEwHxWhtmfz0XHGaKLmpYTBDyCoP6QJ/uwKzs5k6ZN6w0WappEZK8r6p7uszXl9/
MMHyarlC0DMxdj/sMJ3nmE03/PByQH1a88n1t1+0eZlu7DaFZn4OjeQCjbHSlZcGKXslrvMdTIg6
VBapab4KWB0tWKb0tJwVkqSu6Wap/UaptVi8YezXc4OJPsSYJod77ayPJSGUHrh6FqnaUtRGS5bU
Kuvnmvbgvd32m7w1ZK+mab0jT5Mf79VnJGT5j8la8PxkZ1VgTGc8Q2RTD1US48SJ2/rhuLRzbvCs
Nxw8qajOq5ekpEq2SI7ocpeeOaXjkVtQNQsrAa+1DP90hSlYPVviAIirAtTgBAMVUvoZb9Ge+388
pUCD7SVwNaSpDypJ4JxeBtIqYCk3BV8A+WJavKtxykD1eFAN8xRHHKxo/W+HcrO09FIeQ18Vpb6N
WTTWnJ8Ly+Nau0QWoDBSVlrMYCdSoepi18sC2o3tN+o9YKEce5Ol/K6+eHtUQ9WHaAKqhXVzlWT8
j6bIcNkhoRkCOIoOFsH0idmPOJLLIVfnxUC3AvN6WB3DjlX61ogyIhPUckfxT5JowTQ7LWXP2yCR
kibh20mxC1RVIpE5/VcLBxO6zJ6gXQHpTY8Kw2WxjxdD4krEL+3TYuwnF3HCoC0LN00oIzjEj4V/
Vc20GTHFmoQDm1Nlrw6N9iiN5BjHGm7lA8DsIlNkbH11u+n1jgDHS+/IB2eL5QmLHGOxSTVTQYhQ
ZWXI8WT2YCdrogKrecm65o4AiH7XhQxg8xkrTBYHaTOoU5OVIxhA9ee/PO+ebcCJrPimISVPmivW
rxufTsLF4qSrtVpw0N4pQIB5G1R0rw2kHMseaeADXv/LE/Cr3t/TYUPIthuvwKf1ILoKZg9wV+1f
+DDRTXnXWEwMvMEJyI+/8x80GsMAcTgkcHJLfHdwA6GD6iSkvbpcGzhmIMWoCF511h75ZtHNeZBj
Pp08bV9qZ6Ik6P8Q09qdmXNImxmcEoLrQ/6Lfpldjvj4Z42f6zNRtTQaS/gQY0mgbd5OSNAuE4ST
dTTYD5TFon1ZqGtI4CjPXHLDJ+qg1vP9S63AD+q/Or784B05lWAKm+3MnSH1mgha4ovpZN02/VWZ
B8W70IApt3Ecr0WJI0itssjXSYG1bBrlf3rpcVf/uYP09ZXAy84nktQkqFDj+a0ijwE50zgXgVcy
sNolX1ntAuuE9fwaP12LeiesdgiLXegVbHZfgLEm+krudbVp0HBHVzHX6wD7PSSXYRW50fq9px+Y
xNUNRjvC1v+ACYSjH8iuS/2JnY+985f+W6kb3eH4FBkwoK8UmklLjPmiJkr5hmdaBVGr7yuQO0Bn
s/cdoFWHIPqqj1KNtLEqH2ahjDzfHSpLWRFneLiXWFFintQOBbkOVpoR1mMP4/yOSn+9Ckw26+OT
Xdjh0tdHooTc75PPVqNu4d2kwZVgH9ATmZygTqE3Cy55x8pXlAD4V1KhdZZAi0WKLRLMSCFeL3YY
nqi/Hyj1/gRgdqMHB0GivWIcum3TVD6fNFE34BIqteTDDCdM9Tn3q2ssaHJqF9Q68IawH7sndSn/
AEHF43Dr8ipZd2fevYoY90mqDOK6614YjNNlaixSNOmRxGMd9w5+hKzbZVyZufWn01t8dSSkIRrp
gqGlG0ubHULOe5EXfE0TzbDGQW2+lw2CozB93sXBPCSD8RH21iVn5sXO4F+/KbePX0+uVHo4bq/L
OA6/NL3EFA70CsWkcWdljq9jBkbOZaw+fqwJvsp+2hZdz3X6++bMHEG8A49XqC4WL/mkCrstGIP3
EcsKZ9LV7YmDjaYQilnaqLkBNvS+u85leRbRLO5IMp0mz1AN+u8AXebSQRALFGDncv2+7anaanpL
E0lTJrihAOBpN0ihlDnEUBwGG+pfLhud3OfoJROrMnfDy24ysDgEIse86xm1zYL36ULLV8I4lobj
7GcrW4T3CDzThBadUIJBsTVAQ9zLTHj03iV9W1uRUwzKjYtPoZY+wwzbMByjmNZFk5irUuPMt9p4
OyX7eJDpmdih46qlsBw1soEU89xuomm3HsT93NxRzgFxalW7bqWdk+ufM5W1K+9B9UFQOVcUbfUp
FjBrjKBgMrggRcSJvZrqD2Ux3Ik1JG72yV2hnUdzMErHA6H7rnw7otb5423bTLImE3IDi/zaoGh5
Do4Q1R0zGJM83C/mG08KeGzy0/4kRs3+178wUE9ODN04Xlx43Ty/QQCQM9hL4Cbq1OuH7tYGT8pF
ODjrCWBtyodr4bW5FmFQsyoPboOX2aVx8Wc14GAsnm4TwtjU6fZZfD3Fz35tznXEwJ184q2K8qib
lAMseXh40qnV85xRmnu/L/ZCTWS12c9GzlZWahBIga0OFuXdt1joXJxu913Tu85oWIJaSYxzktFh
ScbBUZQ5QuFHTmxC6DRRk06RfcBnDLNKpc3cAFTvm0QDZh1v1zekINI9fJ7LI0cgsvSnfIWJE3Uw
naICjcbkoxBa0q+kHLMGXyvN1V8M5NvwNNBQGQrc8b0dCiIYfVIIgBxoy6An//t80V1H7onqXkfc
8BK+Dmpnm2GGBWoT7BL25P/I9fnB2hGGdK3TV++CeZeBOVgx+eRsTOarzBzkmHeIampUz6kCvIgP
SkLCGoWBv6xdtFzpVmzGs/U/Noz57HTW3kzB80Mjq5LjRy54RVl110TWnR8hGSas558QMbUczkz3
/wXq/7YmahDFxWe6qP3FWa6vJynnXzbniqrrk9qtAQYohNnyjL9BGQIdxnqb1fHUAx8Ko5voURI6
HLQOH0AkPABw7DV7iMe/f2K2UOfw8KQ7s52y/O2usgnA0XFoYUXd51C8dUS9JMcCij3KUUd0GdiJ
Wtvz0qltlZxgMQrys3QvcW0HE/myp2BSU/3HEvFfiOo5uf/52rhPvw+800pzQIp0i2EMh1AShI8w
dVRiEqwPFVdLRC/Y54Db0eckJ5ijFpUVGAvlzh6Cpaz91EieQ8QiFbHxIhUgZ1H58PzbnOgd04JR
G53yUOHfXJHc1Mjqh8x0/rD5i9QUx6lgN5U1dACLhfK+oEwLSXxS+ZlKIRrO0Gskkp7bByGkKb4U
nTopthy5Gde6HA0mhtijNnhQ9VH1WlymYCec1ori6Y9FJBAqTyDdJoBl/rQImtAn31L463NelLb0
Ai6QBLNgV45KxgWMGCVfPuCwNByQcvWtvDjoMnC5jVuAOHZUIjUyMSAlWElYZY5KmJV64yJQRk1s
lu11Nf6TSfRicSJfifJCx+LA27ReMrR0488RwJChYI4VY53Y8r+WDj+bys6szu+kryasdtnh8+gd
DZe8t/DkZ+n+1gxn+o5STc060QKy/mgLTpFr3A33h0aYon/2AK8lMEBLK6fA4lmnqkC1W6IsRuQY
dDFSa8ZIJ4X8MIkgX9NaCdac//+6g7OEMgazYLTK05mK7aDvf33yYrAAoUkjcgzd/v91pQtHw27T
4QunOvLWvZgNEGjV4dXXi1mjkcUjxs5G8xCzkHnGKEJo3vyxmJ353hULK3v6A51hv+JCaGhxq4Tz
i+jNStG8M7bkmu3aN4LiIHm1Dafo/l5gN9bJ5Laa/kindvHOJVx+uJEOHcYfJd72XU123ggcToGr
sXbjSiguSfhcu78gXStuPVM6VsRdXYbcj00mRQrJ4tWM+qkC5jM8makTmjK3ubabB8RCGsvawfF9
OwY9RqO7RlkfuWG1wLkxuZ06LwuSuyJOm+tDYMvn00i9d2QtokZNxs787fNmUVBCDGeJQOR53EVi
esAWqQJSujpws3A0r5DWewuqoh5/xegO5v9SZRg3nLPGsI4oATrj5BitUQrdkiwi3gSVvoFOPdtw
UkU1GVOXVDSzOzHmUuCGXMW3h+bLyACiWZDcaxrS5O4F/4+1mNlAgLoUTiTJXlbgk7jvlYsiCbLa
zNXxCSF13X3uVJxMf8RPwJfPb7GCFc86DLsrj7SIphXl2kxyHcP7Y5i/iAsCvlhrYjt0rM3wQdhj
sUjt/FNZUxSUsOrjk9s2wQqNYoLgE1I8h+KElZWkdaXkllOqLflRM2mFgreZZQGWrWsel7Uz4Rft
xr6wCefjD8USLQ3TDBVxkC0vvEX6ugDzEVlMRhQU1N4jJZ3JMB8YztEhHRZXjiKYKmP/N6htO8py
m4gP4NzOWQeSAScBN3gZedFJdnUtG3EVvy93/B9SDf4roDeoz/drwyfxw5jbdp3Uvk/bdcZluIs3
QpYnAlZhxf+PkUTLDSqlEmi5i8DBDy6OM2I46mej8llfX0QtsT44yIst5amcd61DgVgIIJSSJXqu
lXQf96ZCIirjckCOG15xycAhHSYZRLz+7DyDEEH7On+0EBV9/xLTv4+aR3gPxlYJB6g/7wxEZugm
JcQwGVussXeq4PIHQbklFbLbjcBy8gNbo125GSn7qxUEg2r/zTabMbu5kTa1jh8m7jIjjm6cMRjV
3wdS6nHCM94k+osFVm8cFtSuAFRZGRxyU9KWnWO2iYSNKUGhg4NLFCoBKGqECTQmzDTWHQUGQRSV
xS3b5Y5iUkrODITvB0AoDuUrzTNJkUSywiEJS9uPh7L2ecotx5apcrvfvzr02Bvxzb+8ZYX2orLW
3UQJsW9HSSK60wZxapE6ZejelsN2UFbgvaiKFHilnpkGOqDhDDAm41b9SGaP7ZqaqRkFJQ4IX3t2
0PoPa4ypxmGJ60nEKVNxweTVm4JLzNSU77bJEYRwsSf9wBWy7qHtsZnKwsNxgAl0PhOyROwr2EMu
fassJAKN2UwB2qZZMChd9DtPgSXVLAgmBNqwUmHsX2XRdCiqOAmN8dxxzO/AyWqmpuI9yFY0q4SY
K0Vv9+MhqyZBMN2v62+ZWxjye+KEGUx8wXkTL1kylF0eb2lt3fD+HKgsqmZydF0JEXXCNaKfqG12
GQA9Rcd3rctufwjbzepbiOq4OlY4/aMFdqZIl7Lv6Hw2U2rtKGu/oOyAgr5nIrEAIyjaAOEUHAWT
32lr6Ovdx8DwKwEO5hH5o7qcdGvJ1kEd89ztRmhC+X19Aue3wcsWTgOe2ratlrJQSZZBFO5RT5Dd
oljTnt7AN23pikEv+bXWszT9SLAcoF19M0S7MHpEZcGlMvN0NQZHZzbNNmCLqEqnJWRBMc5EDqv3
y3vYXGU7ishHIBYHHeNrYDcKEZDPa1pSzu0JaEJQToHOhkbWnaGhGvHHJazS365tfLBXGR3LaY3r
hU/AR5uUIwM/Df5jq1I5Y1fua3gY4G7a5LfLg7SjNBJpqXAHV4PCULp4HEOzwBV482EBB5+JWB+Z
hc4K81iPSEnZ9hbwNlkrOgZJVwr/lPHdEOtSWBPALegUe7sF7w7BvtQSz1BvUud7jPqYHKQ9K4+4
r8e5eH0+C6y1sYSZqdelDMYcbEgrR/2+BjbU3A1PQO66A3tSozQjvVXu8AzFwVpbo8aq9wSh21YK
qMya3IwdIdDzy/5LTrNHXZcHQF9TOLR60zZlSnlxTSgcV9HQDKWgaZ5XHKueMfe81+mcBXbOIcBb
XcXAMhIqFzYhVCCNqwB+bE7VFEfQxoHgC8CU8oZeO38Bk986JbD/biisTkK1NQgDcRAdnA2iAYxj
Rtxgx1oJxj1LkTboj3ESh0rFHr8hWHL74wzLBx2r/d/pRxQjFsqt8/T3RORi/K0HtDpR4HauvXwE
tti2KAepn2V7gUbsdEh3lVDdzre3b4SU0HmaTWjbIzfNJVS0F2TWnAxvDsuyDGpgeXsfibHYEtIZ
VWOMtb2XL3GQ0E7G/h6b53xaxL3VR/3f5AcLE0CQ0iiwP7Qc3QObj2gGuboQF9MKAKMo9vhLsgSi
amCs13UhVcxGzVprVS5wzN1DNns+2IlNdup2bbTZLzFC+UjeeI1Jq4aFa+QMZna537DJ9CVpYxLr
rkOw+qJ5sgEzcEWJucW7rZXYfTUUuBUSir5Dy2myfJpKc3AvSf6qlepGl90mJsOZFD9R43nydeQS
IqXnh/2Usk00kAlzhtbpbuqNbhNvQVo6buN0oRNR/9SXaI+uYo5Z3hhIvhlEw2JOVzBhMmJEy7vz
dAWGGikPSzAzu0qYjhm0ZBiY5DQ6YffXp+cf3tD2KO3/WKIZ2kD44i+Jn0sL/Nfs5ckl7WXpjnbT
h2gC2myZ7H/gK+q1Dh6lD5EwrZlf3cTfhhGt7y8PzO771nMgqP3kU3qq7hcZ6eQFm26kaD1I7FnB
CPA+LvppT6AzpajKocr8E4Au4tMJ/7drcrU7fxS4ZiI35L1NxQRjSjjNpqMvfDIPcV+C5Y4UdDg2
S+qTNquGughlMmc6ByfrlrPImWC/2MHpmX0gQVr3chRkR9lLyAqUlcxnIUUY8qTpmwq4Qjd7VXTI
4XUzz2CbtQLJmyMKmRk0EtB3en9X9dVV1zYIq93I37WIRMJ4JLSgghc0ytOS9omrwfM/c/505jdw
iRv8vFJLpoepfrUdVsff5pmC8Pad3nMS5T72g1Ua0ljnTi+6Iv1o5qyGO1/0pgFZdR+EIffUQLna
qgpXOTBQY11m49Ms4JXg3gN9IBvCa9rfsv2zerSpVcLVW4y/sfiqqB75+jLPnsrxnO9byvSHQ3xz
HhGySLDWd/ZKoeLqhFJEBbsWLHqPyzCEGn0hh83slzB5Vt45xI0jMEcoEH79lMCeIkb1aqevOEre
ezS8TWDQ6wqp5tQV20fVOjlON87gUX+d7AQns6JPcmJ995hy5LC916wsKy/ye5TiNwa8dAEPeMc4
kEJJHNzwlG5o/otQU/Kuvi3JFPMdTeIABdu9RvI9Xgy+4xhjoV3QiukF6ct1f1dr0E+6vJzSmpjV
jKhoDmkMCJ09KesKOxxAK7kcK3SvmhmjaXzn/OZ15tvclKpZ3sqY7vMBpvuJlgQlKgalFvyCzuq7
z5zTCynu7+pa9XOOgzwWctM+gbuqOAh3NQplkSXtJESuRYvY1yZsCGyGTSH1XkVrB/zg2KxywxZb
dOdRG2tnyYXNfmopCvVLycdEmeOP3zx1zwGaGQECRc/2AauuN7ZzE+JPuTK/8bdZ5aU3PSkeJFEx
FK70FOxFcsTgpmUBno8w8gIoomAtNijZADILM0sa28EPA6Cs4tTSbGLQe0O21R3/0bMwCjsCMicg
eDVp3A07r18c8V4AdhDaRp42XQvdTBYvPtWB2B4a2UC3C3gNc4UjYMOTkI6GMKihni1p0JzvzLq/
IYp0ZYDl0yThzgZ+HZ/e/DjcYiU95ch8ewovuzLkS1w5ShT3nmT5Gmi7tiBECCOPMrvxLzC0FZ5f
w4Ax01IPiEKKOPU7qk7rivQQu0rsAn3Knjp4ATZlHLOlYSUgUnirNRh4Bj4sYQs1nJno7xayHpc1
hsw95D9vA7QgRwRqi15L5FVGJI6wNRXOJTS9aXY3SRcSG6DwitnRaccmLeqK/ej7ONVjEsuVzAse
JDR39hl9xb4Mo3mOE9nZIwBN8BiSAipE95sgHY037coY3v5XItR3tjbg6aGILZO0Cq04FZVmkDna
ZtwiElRqmp+o5EuUv1KRCXBfjDMTjbqwbqUX4gUBKFH9H1hIDBE32HF7aLox8bMWRvQHDjHdov/f
0taazv9bswmC/ou8EYXoW7RwscLHHYUsZLzdfA3yPKb0F6fl2EbeA1XMhHN+ZjYeOVrQcE9ABmfl
EwCq8jkYbXEjwyWwp5td06HK8ljERBn3WzY86wcgRRK0AzX6TC6v4ipF+G9BFBqwDu9bCNPWo+J/
spotENuaZF9/oX3x9mj8iCFRwL6lh8WKEYp04PzRvpMYUHLPpKi34qMWK/zbDXIwFNymQnKCusK9
cmJ/eRyxCc1XqGRNErz2XsQBBgfXlGY98h0dmrZyocXULry/mnbI/eMRYAwtLUt6VoX1G7nYLHM7
Naafkdzj4kDYtdVsMp+Ay3wajyTeA3w+xkSFC4PwRsTcFYHTG5rHmtfDGF/dcjn/tW44HrbWKI77
yAA06skaj4qRBt/Af2AJdcU3jFhzFVGX3gYIMbJD8PgEx8UAIjv3lsjE/CfMeMTSyAFk6jlakVtG
i4Tb8n1DASe2/Q6Xf0EzVdXRR677luGyFoFqmxR8SrAlfCumCqLVX9J1NFVLKa5YJ9mxwompSe+X
4/hwh8Rdh80qyJDd4yI+haPvA2IqBmSM4wJdq/kHms5kopG2M3QhQX+wR+tRN/cOQ31bcQ3zI09c
FhSd0lWjiwN8FbriRhT8pBG6ihYK+cFoB4PGlASTqTaHEDD3LGxCsFyIK5rc/raXYEfvCMzV/TfG
t3Q/G1/ZAAkxv1li++HrCJab6dn183iYxWyeGBIKChPW5+SgKuusAW2IELkz4qnL4dzQk/t18MYD
XdbCCKBou52vh5m/qTqUxqDZqVnWavmX9z4m/JDdwtfILcr6gU/7M4DXGE8jkzaILHKZ8+Xmqmqw
fonpQIekCgG9jWvIChvwk19Qnx4nkKNFCkPGnSPQWUwHrgSm0SEbxYCcrVUTi+A3jmsDKi5URXGT
KeznzkUtILh2YQ6wPMROaX38OFqCamcJENffmKeOQLdEn2KKSAW0dIqvY0/4jo4JjKV0x2eynXxh
cNxJVH9rqNLGgDFcbLpPsOgt6/afOAnWDA9VQqy4Kb4FccTRWFYIrtKzC63hlmIDy0qXmsfVALx8
criBXfP8+iCpSour+Vq3B35wwd0oL26sFaGx+1dUd70B7hDjtLYIJgOWnnG8d8EF59+IYWzol8eM
HNFut774EwkLxETj+6fTv8e+NAAdeTqg0MvOa/SZtjk82uSjW7okDhNpv/Dk003faUMPg2xt+2sA
XH4jjzVgpjT82mOb/CbWjYAPT8DOh0R+hnTLnuZDr6Q+9JO226hpc+XoLwLlc1j+AV66qC719jUH
4mwZqj9FLCTHK/Cl8QWLPKAso4UjOjB3UQRVL2LbdD9Lf+bZZr9stTTfUFQECA2pmYj4YayTGYgZ
O3ePYdACIieEwPSS1OVsHjsDE3VYwAgZVoDeED531zTY6JiZOhgYJYpHsrnzho+Ad8ihWnEZqOu6
hwABfL1TcFFclrY5Lu0gPwop3FAfOVwKlBHX6p1CZUI1cCuZO9+sGOISCQSLA3VWVa9f9iEExdvm
ZBWO4sRx1MDWDoUtXHlZaBWKS7pFDp27ZG1On2YkjKIOdBy3Yqq0shWwv7kVZdnk7wKk0bhvzoVe
DiglWZPNVnk6pU6HpVZyYfncrfRkz+xVr2KFa1dlPC7Yh4esdKgK8iG3xE+WT7nKvRnmnLavugB5
1NPaeITg7GUILIkxA4uG0qSabcOzZv5IGURvFsql6AxlqSnvLxzVCdEVVMWiuVQuDNi555NYZfqb
vFWXC/4SaFpZlC5YlG/oxcAeFhA7/TLH8aVTDSWiF0wui3iEvwxPMKnCDL5NQItUZVh2cu8zWorG
6bw2NqJjTA3PoHiAdFahubhFVS7lDpdUiyJ0zVwbRMgSTIwQyXm6eAB/S8EDdoSZW6QjTYTqu3jq
I9pfTXn8yvu21hc4tdudgdQlSALQ5q3FgxLpykvgTMBNJh/mk6bwY82J+2h2BgWGOiicgi/nOVEo
UYR+D1Aqd0Q/DNMllg49Rj1YlABwFbt71+8qqqHiCIrWZeTFZC5kAoaaXeiFvjXtnceppBScPOGZ
CAcyxLN9j3+ZrRUZzAeRYSILVh+BE11IcH58kzJ3/fgmw2TwER53FzHTjNQ1naeE/3FDrQ8PP4CO
97pwwnWBjcnDn7ITDtlcGsBYQ71LJGeXyjOszY3g2nTk/g+iFgyr8ey0sI0iWN4+CGckAx9qRJvu
7XdUIzgH/RU7f1XwHG9sMCng5Wj3p+/UIEXmjdUNkURK1Oe7+KR/RGzOOfiwlGXCH90UJLRiOwUr
Ko3usScwKZG2SC1IT+CKcGDL/AW4C106TEPJfZGi4tlPwtkzUMLO/uNcE3KiRxrifnPDbn1K+u9k
92R6HSLxDE/Kni4W+h0loK4Zz7EvMUHXGSg4xPBi5At/s4dy6BV4fWCZRon4IVWV/Zlhy6SmFJB6
7xR6Xy7YVpANbLy+Q/weT0wZqiAhfvqqRyNkn842UJ8lIzt7IIo75RJ0h1QrVwnIceeiJJJh5EUI
Qrl3J3aeTJcJfEIZ/gkEAbcQ0Fg3ujGiZEWT8V1u5w64n4OF8VF/G82VTK+ivgZYrXJVuiwE+UPk
vVuOw7wKP9OcpP/WjdI7Gj9kMIsugC+QvI2NnaGGap5bdrsP7G89HX4iabj2Km2K+3l2w41HfPEB
Y+srq+gnvqeOaNLeW0yHno/knV1BSuwRBtCaE1PylNvIKYrDc4uZmcVb7IMvx5NEj4l9zUZOclQZ
SCcYpWMnrZbnNEjqJuiS6hcgAVdogM2M8am0EWbqxGwxGHL78rkwz4cyXJc820Y90EjY7M3EVkWN
9iv7PqWF39N4rgoJX7Mess06GYc2YOyGDvn4ux976xns/Bs3TrdeTxtaO7nVN20asRtrLNFWjM1o
JzNAwoY6/VYhnQ8KEsci1dSleb88bhpDw9+HsQHkVdnXpifmIlEPbc1z2xxTedj1zkDD4ESJvzIe
NBYjwwSfCkjHzIRZQKif/7/UYWKGya92zkRa2qYqaL5LK93Hii3+vpbdwov0S36VQQcKcoUgdBpu
5xA83NwFht5lVjaHkD0mtDp4dsnIPX9LmxslpW7ZxpGxeShtNxSER6hpO/eFjo/MYPSbRLAamnHt
ZclBQOto8lwnKzrVtTyMcepHFfgW3QIF2YTtqcwGpwktyJ5aafRhZxFattKbepn6h7AOvYMAn90N
2a9vvbywCo3mcg83gLjP3VujOp3HUi791xt0S+oLB5hKnVSA2Rdm3+vjarmEUZVEWJvirPtCZZSA
kaQXz9s5n9NvnZlO/Dur/kRcWi3H2KlmeVaMs7+9r+2vdgzCKru3apYmw2q0bNl7H5yzd04c0VrZ
eOuV05MNx6vhSdlVPjthu9dlZdG0JqeaXENE787p74i0UvrQjk5VOR3nmcey8IQ3sm1Xt6vlCqoM
ZobnElq30834cjeMyzt+Zt7ZIiFnm02WRzXPGp6PKrBCclrii+lzsaHnxVUwiHfte4AJbd9f7OzT
l6OzF1U1vFZ5dTAlmOgnvG/J6V3Hi8cvePSj7KnkwJTNRXoZ2lEB2J60ZdTDNrA2stzZe9j/LtwJ
KOVeusa9VFDQtMfUzyH8qUps3UP0MIiq+1jg0vFkGpcItzL1DWBYM7TU/vhyvsOpOydRRTOzednJ
U3x3C0D35OfJaa9QbGZ8RRHLPSbJzaKCRZOlJkU68ZoDSttUhwKWiAcBSZ4o0A1lyeRJzHI73omj
taxaXG1Gu/d/MARzyA6f7iL4JDfY3NE3E0OjwRNnj4f8TM/hpVs0uH+tf1MF4ESD84RbTb8wBfGD
Ofz9upHTau9Gtt05Ol8se0/g0X/5kzwo9syQmuNWIkahon2IdOEIPUUii3PEEU5PhB34jX7Rals3
S0kNHltksLMC9wGKUKY10HaThwK+1V1PFpQgDoCCuxzino9uLgnDEIfJMrMypX95tioOum+4IA3g
jphhR+rY9w3m1hovKghcUxNcT8CrGIvGN3YUOddDeG2kyrqBS5QXCGVg0lghrB4nqqc6Z5xDRHlr
euUCSmf9VjqvNIi1tEKHccdUJf/tvE0/9zHZNtxQwDlT4uUgea+NYMtxzKDpTnrvBpJa1yBngmq8
EcX/uHp0HzIcyMepXQ4kS8xezqaw+pE5eaaL7uT+3o/AfSApXzMEHIPBiiXB3xAMURPNUtRFTgve
01roO3z13zW7S34EH34ZmedlXCzEI+OFEeRG9PQfryCAvaKkIL4npAZfQ3ufnpngjHj443cylzdD
XLNUHtf61u782Petd8bc8BTzossa5hQzSoh7fnVHxlL63lbabYWmtjCE9q8nb82I0sbw2/7Gjw5K
12hBWvXgNIQMKRDdgAbbHvkBe1JkwfUVXODnsmWtlMj/tUTn263pjoDuN+Ad9UMG4NH24F9bSwj4
t9MNZZ/ZbFT5vjaxSe7Mxf4np05zGOr8cvydNeyKaFljvsOtvAhjbCsHoleGQOlbt5wtyxMTLeRv
PQVhKBUvzwIRzK0ajCbkqhfgwSsjKfQrRhe/rZoZ5gW53x7G2UHwj0RxECldC8HGrtOUnIuCP5mC
eht9xqwt0u1+S4wCrkG1x8ul3tRkP9stPlYKL/wECrSRhgPtFkh/OFFB7aOGOVJCRPSdyNPj6DmQ
kEXzLgKsAFStqw2Re6DDs0XN1b+3yZ2gGXY8cYBOqbvt+ueBdG38VMI3GPq/OFl0i4EvVDVwsBmj
Q57JaZgrVOm5avLMx67Y0i8A9SEi2xG3+fjY3m80mIxWwXTMshy+DeGAYVMF14n51Bicl0oOKnbN
wf9ACle3cRGInmj/V2c8ZrLbTWkiZN38r+6/HjYtBQRw/SC9wnBBXXEWx5FXjj8Z3XDqO25f1mLt
mg9es7SfypUyAw8Kuieacgl8ZLcUvAEcCtvKkD8miD9Z8Y4RP3KdpF179+U2ggjlTSQWjuAQybbE
KTfr99Z6HFnHjdJsuI2BOwJ1ruNx75MMU7EdEQCKtVSYvD3QJoo5VwtCcEhhxvcXtdsQirthWJOS
O2uZmgqAW3q+dm4PkdFrDJMzTcb8RkiQFP17XFGZL5+OSoc/K3VROT4ZlIaW0dQfhzkBiJ6fPVEe
d9KCyYI87iw0sfcCfdHDzwP19ZVM2u6NbD54dSHTFdFCX2GxNE32MSek2jV/ozAJqEUjtkr0dzNt
41Zwl0NCIcfgewOrvfH1qN3xEBM9cpUTHMlGt/pjm9OSQp57p51Y07oCV9WO5bjv/aW6Vl3k1i1L
A375p7EStuPWKy0ZeKoqS4Pjz4xskJB1pYb1b+Es9WRyOJi95tniD2Lq3Huux9WS88ZQPvoyv7q4
fqroTJPsZrEmliJZG9mTH62ZNblWMVr2xM5CFi97mCDsgAjY7y0zOiJNuwSxHZlGO9WFFA6ercL/
pwWaKLYAVmo82XMI/QZTUzWVlAsDCCIkPsdUWeNKTEVQ2PobtzcJoQlnzwC+XSW8LPHsxnnfnWc/
tjVup9RbaBPIkY49d9kKp6AcVz8Djb8t/T4bHTIPQERdSuKscosonlNYN0HepcKblhBoGLHA2ghG
+WqkhbXz0TSYgb8MmGYx0rEmRx0nWxrU0/MEl1SjZJ7JEdhqOx+ofRn4UNOAyUlJhgwOVN66npGX
aafdWs/oTR0RH5/Diq/y9a6PzOJV4Z/CUT6Q+PZZLSpxm9nnAcEgCNcVwRKs2uiVMI8CObctbmOq
QY96ssKkrpskxjRijkFyN/gF6E96oSWXSQMPP4F/WfvLNS0yW0WRvHFUh/YqjjB8YjAz+hQd0i29
yGOUQyHVdS/gWXF6Gw/47qKX3eA+Bzn9uLc0bKI78RUS96dO88nuqma1zJvrXIO9vQLRPffdYVtG
+QEH6T+5e8RXUEqr05HtBJTRdHWJCZZxwH1oNlccfurFsNVmIZlXWZHdk0dfiVbd85XqoY5By2LM
1+ThXgpgR+ZrF5PhXVntWT7QKJYSLlSLwgaXXMWVrfgBBbYriLqRbduUdGwLZQrh2Zu6rTyykSAN
3XQD2Z6pzn5Sdz94di+KXerqrYlWFExriekhTglFbyRjAWAZlrk29WMQJdTrtRuTuzflh7/2oMDU
rTddwXqo92IcoInaE/ATz4Y64ut3WyKZIqLagHO968Sug0fmHGX55eHHWsSJ0XZvWGHnqmw3NSYm
3c9NpPPp4jh/p3kTtE42QfzmI48ybyZfiG2EiVtjBOwVZKKJWDwO+3BSNWpDezX0+llCarsbDra+
llsI5U4tnUfMdOYmn5k5BlGDhYde1sJgBeXcK8LWGp3G4Q0lNhgU14IQm1BEEQdQj3ERv23PnLbc
oNJvzLgfG2erI465UCfZAhXiJO/oOS+Vb8gnTGIlsfKXWTOq1kPmJug9FZRjHK58gQLOXRd0zPZC
JDiQkuMvz07gXER3bEjX378Y7CWqRanIbSEb6D+PaS8hNYr2q+XSRcdskbosb/JdkheD6sLAl1W/
c1mGdAgeNsEvINYTOkZMf5C8UdDWj/r/cyH2PXwstmVMOv+EELy+mxd0z3Xl1S2JxwaUczQ/n9uV
BrLReQwAWIVXVEv8xrlTBmkJWnCGzhVXwGqHWshvuYq+PVm5lufLLkqZvyO3AUmBq3S9NZFlc3UK
Naa9X326KXMR8ZAqVCS1D94wdhmDJOM6vWN8APU1S2cNwYDzKDSc6iZPxWs9vhuk/3zEQx+krn/E
cGmru542XWWGVVbvYcBch5m8jvQll21SlWwqyfsN9dObKpZ+hJkyOUGFVtDLkZOhjw+etdWg2Ox0
VhBqZZTQUcS5bmiSPmTzSn0oB3+N8rpZ7jjWpIO5lcmzJve11Lpi+/5byk/XVtfcp5qemLNDkoYl
Kxh2eMuugdi6uEjbSgggM3NTVsLY0OCmqDmwgEW2dZCrBi62SFtEGxKnMyofJz6GVCYQYghyvxXQ
16Hq2lXz845KHSNVVd2Io0ysQayj/ZvH6opWkkM/teB8GMeAMor6DVe2UuYuJQaFNHAEokZfrvqn
KeZqTeqZ0kjb2z0dm2iLLOkWLWzZUCCmwCkXpm21r9Y5leo/GcwmDKhDXwLVPzxJH3Emo4f0KIes
NpfxPPzmVJz5s25c8xEMcIQV8yJ+87ued271BCr/jFu4iFiFoHo+cioO0VZo9GIGrHWniWzJWtap
GDthLZJtcs9y+QNm6umPMcp5sqRLOS2IO54qv9wKOx/pUsZG/6PtuvLTjhRvyj7JNt9iYrQzKFo9
pHvScVV5BUwgZje5bfHYJyTyi5p2JnS7e6Gp1EuWDLa1ICIUVlKTfOZqT2GhqB1cKTgl3ioUE66r
LL4DybEJyIRcgADnH01Yp625KXQOmWFzMYa7oLoTNlCDOMgfk8lCFq5xGRaeTqcmSkLhYramqr+m
wiEO32hUZoormaoFgq/B9u/NhkTklgbnwI17Z5r4m/u8mp8YQGmBh28RGFQXqAyl/MpdQ/Ctvzl0
srHA84DhmM5fulILtUMxMwO55vyweBHCHfyE1clJdKXz64/CQNvC51mBAdJBWW2P2trI2MOasE+s
AhJIkxCKbi9Jh+zd1DfRJuv1c4JIF7JWraLipe0YWYYh7RkxjrOq6zsUSjuln1xp46tQTIg80FjZ
7q5y4cYNK2LJ9AMXL0EeNV5G7FuoJS/NoaOA4YyL7Cc4m9mIOmpF0EE3WBJcyIuaMDJjEz65RK4g
4n+lAnDZAudk6HnrSMKfa3O9gFbYLHeX9kp5yZmDlZj/AsbIc4H5MR2DzbB+XR+R8pWFX4kQwKTg
p8tS+1vUmluei8SXkD2oBuiJiEIl9kFL4jbL2FPiAFAAMSyz1TW5u+kzKDUcVCKcWG4Ix9laMAUX
P1qvuDt2IHRivPmmdFqlm3Hh2KER4XYOMGIMYMg23YsEc+uNMtDU0ekdDhPw+nTdDTcDet3joF6J
mOcGXgvAZa8Mpw+frC3eIPGDv2mOYFasEIIc21qGzpFtFbYtoDUy7EmNHgHkugO9aZjOP+KEaHiG
5D/98nBC8EiY3ooyQVL3fGyOtGoBkJ16LXHJzzG7b7mTWY+HQjLO7JPFQR2zooW35M1sJLFWdmrn
QkL0P8/81rTG/XWVcQcZlN9l1OxzhVE48uZS9fl/mgZvMqKfz3TUCZZSkQ0UcpPdzV0iY566wkUr
H01EeHkEZe2hGi6ghpFH2jYw/NFYZ5JMKWMzOhxrJ5OWAllKWFEf0sDeRj4Ve2VuqPE/8V5ny5kk
boVfdVzICiBniqa34WuyV+htfyg7QF9U6gCHwgf51qxXnzOzHlvvY569uD2gyuyDgidUQS+FR1Xg
gIeXlU65s1k5CxaOypfXfF++fjLOM7C2X53J0ixg2mLmu614pe1lLN0zGl9zh2usVvWuDkHkpZ2v
Or9LYPZvhz5Wed71ZYgdXChT20/EiINlZTVYFxZZ3smM0uAUtReo81WqYG9mw9+lgFCzXS09r9iw
LWo08/ZpwN+SwVO1T2AAU+JhBddiv9Qb3It0GIMrOEuYpvlSV0mJV71bcKTp56aWKD0BAHdIBUqo
xZbwJsxrQ4eJj8mZ8tDVRKKUN6Cc7u+Fy/hkMvdO+GO6WkjKPfwsSSJTDsHvxQbxgtUHZnH6p4aL
mEn5o6oLJRsQv+Xvp7JNv/3pL6R8OC16SCSmAoea4OhsOxlPV1yLP9wwUcz9hnclE2hzsVctJNHt
qx3efDT/0M8S3oBDpgXMAYoi7g9ydPW/iAI6PaRU2sSbO6N/ZeQWnPG20+OwZN6kEWo1Zbjs2fyU
+mPAHJgaIHjS9+0x3kvI2aM7uEavXr+V9lMMbqmKerjOM0GqKvw+t2uHrWGwBcsJuuEuipI0WM/l
sv2MvY6bCEjm95ldPsvqgK7LtFUf/yrE1HiOBcAV1NoZm1iqNYkXVwp3POn6ElK9ofODe1DyF0/3
K0gWMb1pf+XF9CKdEl9vpJD4ZPmlz4Y/33oCpP0PYipyTthBw7Rip71CPnV5EbCq4SUv52Ghcz6G
CWznrNDdAdRJc6FYzqzUcDgIYaCaAughkH5ruXhehokBf3GTeukulF5amdUbCBjeqxtJXAEriwo0
nEBj0JWmxakqcaGGG2gWdiyf9JCrw1+KpCGtTVJdUYEkjjUDszatt9KdSzvLXLzEB7GkgAxI1JxI
zVWFVwi130QXedwOkRj5R4ciI49WCopjWe32MGwi25iCrdL0boK/gc8gy0FjttqgxT2Rk6bpPJx1
Aa3UTo4ufgaWwT7YaV1F1/2kEO+cAMlc0yt02jOE6LYnQqcvfNrnd5GhrID1nQFWbu7bnnnwbBkQ
k2E53zNlR6oFJHfUkTOVacwr687RIw0DHmVExr/AqQskLACNDRjBgYcfAMkehBlwYOrVR17+94hI
yP6tGJ0wu97mKSzdwx7aAtecooUh9MGvTMsz8mei8i+QejLcMQn1RIpSd6MAa9nSCnHBhE0UrXsL
rRFv2nxv4vbKOvp8OqmfH8UVQ+J/VYF1UFt9iMZ3rdLBZ72ahPaocN9fWACgaVG21k5GdEqpNCz9
c2IDuPSZORBzAjzzbjXpFwFqyG3PBo/XMWwNlzuiRt9ehcL5iqiNeqqRHXdJUJrMWK3P0Ho3AJN+
LP2DYq1Y2sDt6m5LaDMZK++UcHFbw0CBmGirPfKWJc1k+pRIL+0nr01kDvK5FP19HpgKpIAfttIc
4Pb0Add6kTSjUuRGwzZwaGmfLz7i1XwwUB/FwbZlph1egV+4P3lalfUoQZxssUJrSSEp4mddxxsi
9XPf/4CrlrmwcUBNZlz1B+HC9/92hGnLrhSwwv+tsis/ClZS08NgE0dhklxbqVooHosZV4CbDMIl
f2vPGwG7xInZ34gLG1NHBWOYGxq1WbxILR04Db4vDmRK9NYPOUVSkGoCtDUCRubEs23hWCQGUIid
L8ruoQfwcYAeEbKiQQGYybHTrGQZdOuQyiZAg9La3l5wXWPxlFJfl8rnTY9LtHvgj13mxkU9qNDu
8U8yMq1m+4xC1z7TvriMNZ9TIAtbynqr+yPBiTpSdTcOTKwlVZCDsQkCnlPDeyJkTAnZLWTh/7Pd
Cq3XTIhvx7B56zoZonB/kL4cvZs/i7r3eAmd8ZhjtsvrSQqzWNSTosW8Z0w/P21bXGdMTU6NTQH2
A8WKda3o0cXGuOawcpTerihVVTSE+UiyhkSYiXOtLzGISPb62sVh/cxQnqXRYEYQM1/oXKf1SArU
GmUi3eBmIowIEG6sJThjHpygK+hxoEtcMGAa4DSLhIt+QJdorsuJyhv+JSNQHgmB8h22449SHUw6
6MaGQ/luhQWISg+v1RioxEWKLAaD3KX52ayfWP5vcA5TR4SlM5nYM1M87xlU9f5xj9LboUCa7fz/
I71nHQE4WGMAmM0t6CqQB23DoY8YPydONO2B7cmyoZC/7SoTe4SqikrlBVaFKpilLzdHZ5KiIPRR
hdc2h8Ogr3tZHtIinYALrwDqzMnRz5PAlxpVvcsCVCnZOVzqTqaWRVoDY3kxk94RM/rJKbN7xHfR
uI1CtOowe+Jg7eVP6zQvzborFMcesUywvyUYA26utWG4CapyP3dn05wFma1Xc1je6cMrSQsL8act
kaVpkeYZzzjHkIv7jrLFEDGYAwhrV1OPZTod0z2weQ+N39lBC6JMGbaZ/QdaQAcnrr6gYcdPXBmP
4Ek3lIhYbAwnAwwvh+kRkdlJKFZ4/aUlu9Ix2h1Jco5gpLnbRWXnNyDjE5E6TuhxOfLG8vCsNWvo
gDt/rGmeOJc78MWmuGmy/ihl+JDjwEyCSTeltgjMUg0PnH0Ejl/psB0qZWUCTNg0VnRadfu0tS+i
0TJyPz1tq2uvgBMUHFEY2ZqRXJrddvCHf4U5aXxHaxpb4e1AEB2aExsY99CDz3+awUUKwv0NKL1Z
4EntFFZfcmc7U5Ck+5hhObP0Q23TnnHvkf1ZpC/yw/Vv3YqBGRkn4rTc9XJeptN+kcFi0XugK8Dm
kUGl4CfUedfRZ7rTBx/tiVQ2mz7jTpm6JmHXQYBENj6sDS//IURq4SRzqKhTpqlUATImw44u2eHv
5SHF84mjDZQcbFBAWKrsuNuvKxPbK1ecNq4NkkYZO1M4q+YB3G31xmHsI2I7kPngep86pGrQqMUZ
8++vdDZ23JnvNZ6QL7kt6oMUh3Ym+WFZNFzP5U2Ks48ahLkNas5TgXKe6dS7ExsLwfJge4Ga6nUU
SlpzkNrXOX5xvqBtO1XEcdR0WzWz0xxgNdb5WB5GfgMHFDk96nbv/S6vOmcIaeG/Zprnv80Qn+XF
tPaXTF1NiC5he4C4g/hUvMqAJ7EkDtqddgP9gOoa++QK/hImz5hs0pPMjOiA0wC/HLhhe4TNy/FS
QWq90X/CGsaatBfrjA5/F2VgdxZ0B7nvGcZLkYoeQzlXakH7jISyUPQ1gThqcjZlVEEljZeFBNL0
jQ2F4a6xTV440NMwrizyXJ1vhceG0LqM5IGDECL6S7IP27AcauVOwWVrChuJUlIjgZg2gmgl4dpC
tYItiQGJmLcpC9v3AYC6nx77eu0LKrX8k3fYbjkyrO16wPTSHDRg5HlC/4GozPuaFqBLawvT1Hza
LwxTN+sB0wOJBujp6VpHNngwskertlNHb4rMSClD+T72iGWOsYhV/kSe9Jxclq4sK56+8YqKe6Rk
HtCf9QP6lo/RHB6dYgp1i+TJR4MJk+oQkG8HjYhEKpObHDbCGwL3FBWmpKqNdf+PH7VG/n0Ybvno
+XKc6RxRKci3EhqtsOBrddq47mPpYRsV4abAEAvDQfPGEclNckUWg8K8cVNmY8PYVfNAizs7/APy
li+BzRHh0UIfgN0micuGT/eLUU2bLSPaCms6B7tcAm3Uqry7s8DbnVIkwq+tBX9Zq9OYgXHrM2md
k/MoOkhgYa6LCfBIQKot4QER5oAWv0mwtLM+OELK1vwnuDtKuii7Rd19uCExUOjCG/gHnIIBb0r3
eTnyvYg35uI2alM5Y0D0ebwPsJTK2RZfCHmprEnfF8VAHyyFH0LwNJ/VYfOodKwS6oyz9YMfbq1A
ULBwvMB3HqusSlMOb3fiAIgBjCsB7CI5KsDbXYKZY/8xmx91LJ1RWVyP7t7BNDQNACtvOJGmmZmN
Q/qYPqVMisfF1ZqwkfQ0UK18P2Ku3EA71oLdtAcymWIQmHr5jqFYZnr5pdgHOpdUiP8gzKotPKQO
X6W2j5RSErZLdejjY3rrBSuYEw6VOJ3gtXefDQeSqxJaEEB2vnbEJS1E/T6IUXfzqSjj6WF+YGnP
SOcGzzo56alDt7940Hf2fQh0vuakNX0xvzyYy/+Nz5w/C5MuYsbyhlrBar9BabJMFVa/odxZyTnN
ONtMGs/KPDVxS0u9yiazNMMng046lBhVcIIALuYMeV8+Nvmaw8sX735QBIO44JmrrmT1SjhdOwzw
3TIQTONwTfFZNeQB6PVA4/R9isRdF4j9K28/KKdKpmzkdyysjmTyhgiUhDuEBxS6ogZR3tkRAcg7
4D7jrX+dos5vPYFMmYM6EQizM6NQhcufb1A07pspTcfdfID6CtegOI+L9WKIJHyFgWqfIxTtJDyX
fk4iE++my1TfmgHOvDuU2nuFf8kDT6uoJW0hy8fHjBnM0oIz7exdCvbDhnO4LSzAuGifNlWfYLxo
xO0RJxlC/bFczsCvcW+fIxjgkZF6FMs6dw0cLzf6yZFM9PTCRyo+6VwChDreQYiN2Z8J7HHpJVO/
uIZGij1bfIcbIJwXsJE/E+fkgx5JBTWJ3x7BmjTWscueKdQH8mNizAS18LnFNVXDZjeP+/iWbBN/
+vphFBJbUsAvioLA/1m9rnW6qFclDV0p+W22TUzzuXn9S1nDjNGFRkUdyHeb/YthDaJz1o1vYtdw
1yuVOZVzWGQk5ZVl2fuZsMxFH/9Kujrred9nmrBkVXx9uOJf/ISHxyuzt/1WJHe2sbnbxTPlP1nK
7qvQFXM0IlhFG/qHCzM2G5fd+bSvv5FYckk0H/GTWv5FiuiYL259vo13XGEeCIvupw2hPlzBMJIF
dY6WRoSet7rrx7QDU+xP4NNSC7M4p6mkFQBHAmnGAvuwMciSnxPe2oAeXo+UCGfVKPTKwVCt737A
hC15b4avKIwolhBIJa05QnCweBDV8jO6vvq9mokjK4wINHtZVRWsx2M9bbhVoHQx7PL1elRv3Gxp
gFAKwO7kIy4feqJpWMzbVnDqBdemkZ3YtnknUgLRfN8cVWprGPB2dckKR2sfO7smwAWaGVDOOETV
HiJrzHJI68nSef8iNI9Sx7AH7ImMc08w316USeOHcDfWtoUO2JWBPJUwaUrgIGJ+MSyIcl3cSibE
Z88Z7ZmjOFJiehwif/U75kAZjnEV37vLX5G+51VZsPVRn77stLvLyJmJwCldXGMsKZ91KkYmiEC2
cybRNo59UWIsuHgFdSbWFxnqcWK/DZrUra/9r6/78wJRFP4qO/aYhK2ngcysuBSDw7Xy0VecNjQx
+wP7ahTxR6xIkeHRVsJNiG790Fc4Sjiq751zp6oiA+6ZBjvtsW3SLG2HEeW6PjP/CKxrczBUwGsa
M7qNJEoIdiR9Q3bOjRBoiuRHVHupAeVE4PxPMQE+pEj5g8TXD4tDxRcMhJSnWx2a76UR9snd08tf
5LbRDnh1RHk3XdSlujbjUj2EE9dU0I0L8SSOPRcQJex2mp3G4ScYctHlwBbhD4Y/K4RFpofKalJ2
PcFqOuT2fKql9jxNlV0YC9nxyzSR6o3gm1F/QZKRbYvLfTuaq7S8ep3U86/Yq865+29WSNgy56bY
9LJVJroIrg8d89iSu3RfiY/n5My1UGiEqqn6GWfeBtk5bNFTrLfuz6HSNIAUIDQMf6MfOjXAVzVf
mWqBcQRLFu7qWnf4Pisjab1ElbZ5WpFaEKxqqCmqMgO8AyADJ082vybgcUgOcn0RNxOOVbckksa6
+6UibXZiVHhr3cIGHvzRL408k4UdKo/KkEJHiGTWPLoVPlD7A+VkFqGQuzc0fBxxAN2OHSU3+LJ7
FNRdqoMxhUNaeJV9EeTWgF+rRACCdpK9iL9LcWmjgnQej/SJUzDzmB3eNVqf3bI8SEOSvxX5Be5O
oxf+W4Vnea6/UjSIDB/rI8ErqptadbCZWMAikLwjZKm+Rd4xeLzTd2t9PS2Z+IwSSCsv0y1CeccH
LHYZaYOrwL9QzEOKS+fm5BWeCcWDVfZcd0/EZ3NuIB0zGZSsV37NONt5izzgrtIptry5nI6jxwEG
dVBrRK7mQZDxdKJUwxjoIjPWb4sdw3Wha4ClIB6nxBowmOy8fHVtHEFNyESL1No80XHcuEiQmR32
c5NMasVvQqtML7YlOgPgLsnpl97+NkXn2eyf8Kks1srhdm08J/LkBYpRhBM3OltcvsLHki+kyjRm
MB8B6+J/z7G2KRlyiTPTnrk+1oIlV3cYY5iNHe3qtmgaxkscU1q6f/YssZlbeSvLYru2akGpEzN/
86nGIu0M4fi+MlTETn2cFWx6v14ZmprseTAhUvV0GEzyP5EAiD1Qe1frLjsscDeG0KgF5fdrwv/v
omuttN6I208IW68nvPfIcGSPz+vpYt/ZDmTu7MFbuPEsRosU644WHFGGRzYWor8ZuJFFL8Oo5Y1+
dUmz6Ckf915OsiKntfLVkhuRy7xftpBEGqQ/Yc0G9IRhQlMxg5CfEiST96MMBHsoEbbLHhqUtRpX
1gKXOZr9EBSlgRmB9Jx+sP5jv7tX8/1F9BELtFrVwwBBNt/ngQWu8zmcEz+VO41l2bhXw3gS0mAw
Sja+g2cX8KY/D/UpfR9MN++atFaO5r3bypSx0LunNxjPioEn/zrDjZlN1sy3TS6OCdBG3cEMjW2S
DAkOg8yu4d511hWB6NKT/ZbNLlA0lGtlQyj26iA/A0Qa7CbZOZm3A1Nr4CB4xC+CKk95CU7++/KS
ui27JXI4RkM8Z61i/SYeJlQTYBRtATUGOVZi6i5sy1C9IB0EbIwQ/2ZAQLzeOOkaeHfsutA/hIcH
yVrvxnyA3mfxiFYgyDzUDUnoEg6rQzOIHhtOfYp3P4M/9zuvw3G5XVKsIL0Oj5RI/E+Rm1wzsZbx
vdzn9FsAP/7pRCwLEODyXTjlTQ8K4E7foDKtOQ0CIwxuyGOw1KNBUA/liQxB3gytv3m2kd5Blk9k
Y5dseZ7R2OeJ8KdQ7rkhPLkDiM3qU38aVabJAXm2qQyBCwK04NbV4kLKeVthozCJ1cFagYdHHT20
ib/mW4FgCBOKWH80ju/6Z5OvAaNgia0/U6BuUMDuA7e/whpPfsnVcMfkEG/K4nLVnI5Jqy7fXHJ3
2mOW9xRnxYzwCo9Y1XIVl1/+nJbE1PqIMz9ntmfyK6ua8dUtzdQXI+snHhqQhCEU/j9qAQllfB+3
xX0pdklJySbjNbxms3v0se2ngDywoKxtCAWeSoL9cV4IEYTnBvuj1XwjhnaKVWIY+7QBng+w2WQk
H8q1gOIxkBdgHw5K2Bf7QnEa/zQ5JuVy3E6aTC0dJEl7HyVzabq66NGSuJq3T70NXnOnTwO6mD/4
T1Xnj2yUB4okUn5mjnUtWQ59Lct3ecs3b27xrRIZuog4U2iw84VW8+ktHUdjDqZfD1+R97efXlQg
3deip62q3CFZbnUsFg6Py45hWeMYcYxgvg0n7SXFh4WvqIXt5fqoyfctOiBEr/iN0TVAt6grwyE9
U9KAnJTTOp15jRHnoIml/N6uinQnKJxp5MXLZ8Duqy47KF+QXV8nKucKx6/nLoY/FDDO8UlR6j9/
DiDbf8LIJr8oGetNK94HqZLjp3yzJYRmCu61te31IFY9Rgw8abz6f0anL1mV5QmTXlUCTgpFc9zs
W1F1MvSlMYJs0qb1djgnYkv72cDpdj+Y1cLdA5WTK37FXr1Yi8mWaN2pAsOxsp86cFAuacccaJFt
/jNcXZPAV7xNscdtSnV2MD5uzvdW2ZtnRMZqiM33MC0xIs2iU6sK2FRyymoihb3z454n2lrRbL0W
QZV9b2eNnMLEk6PWx7Btiir4BEDZUpKIQnjor6zYn6bX3jL73QjHgvCZGotnHiNHqkgk1NDh5/uV
NAWxK0v0G0c2JnkD/mA6S4O1xAEZVJ618XX2gmUlwgVAAXCbX9zDBx4OeR/JRKNytoLP/1VthkaX
Ik/HXBIYNs+jS2CadWeEkUpQUrF4tuXVWYhgQ5cemvopae1gsFgyHi+nlHAG/pA4gUmNK/4iaZcb
dctHgx+B5P1ghQVUXNfLReNGo+Mphc5AA8czBzkZSG/DyXl34dYKEfFhuAclo37thTM4VK1nsuWa
ALzFOXscBXDBZdFmEzg3AEvp0+Kq27mbb0pgAEy/Hl73phkpQzKvbD13DFBN5OYJqYvYmAuD47xW
5ttMwWzajt6ZWgFri3PnBK+jQq5Aua8bh3r5FTEpRrlmuT+ZNSucxFCHj3QvYzV3VMNZ8QjxRN8H
PLh2UCj/STBi1qZ/CXjgom1iNxFPSfrCsBxoMCYyLFKm3+N0pZAiZ38enDu357y5nGQLtzyNX45F
mNgzRZxatPYJy0oyOTpX678tacyORp7MfJQK54mMtIurjljoUc5zE05bRwnXu5OhQwfkTKJMNoA8
1LAspIK1rHGpWedVt9d8NyWtWtx7wfLAX8x7fD8+ERpEbHGUIkMhevnVTi/VRilYI8VY6G2k/zWw
Ox8eu0yhn9a36TgDpEn8EWUcdHXs7VSv24mYq5tiABOxdMVymZJgT2/XxIDipaSy9HoBSjucSyMX
eEdEd4tNUzrepBpHfeuUpNazRyYR/1uBhkVf0o+8b7AZ1R8Zjp6kreB6mvW/OFFtP+yKoybNVGJU
MRHUZ9obeYo/Sd6tW8Ti+ix4L2iFY/f/ddnVW2voNWi8MMHiRuc/A6/MsrFEbIdvEnviM9WTLGM5
7e0E6cGhSHk/1osNQQ69DeR2E6I58zx6DDwg0T8QNNzA3MjrMbyZ+mXPGvjA6/KbWvIwfM8E+4qq
JxNu4ruIc3UgIW+asg9g0gJ/sivXFVYvDWBN4ELHjyb7zQPLRDHjyOhG+iRIp7oIuExoZShO6asV
VDLMjUJJ6mwORIMCr8dBBiQJKj5L1JNIZA4iArIBvD1ZbIYA2bkgRGmJbk8/a3DaUleidt3a3MzI
X9jxDuRO+qwtaApoa3dpP4r5M7er/a4uJILGsfxfRe/tKwZQXCIgg/zw2virhXPCHs2120YMZ63u
3eUs6UVKPLvBcIJWj40OuRuC0FEwao8beTDCXNYs2MGvIheXN615eq87fkS3dnSk5RSg8QXMEpuy
lepIREyjypfIk0zeFZM0wOg3euQzzPjXP17wXSOa7IlOfenWvJR76kv8+2+V3VetRyAWc3RQt5Sc
EMdV4gNfFXCINtP5ZmAk65pO91BLI1WjUmgiGU6rivWesey4Fo1SLisw6pZ+Rwk1TUnX7iYXNk8g
FA0Fo8379Kfy8BO8U5jGO2HKN1QOY8+0Kj02Fp06PhkJcG0yEYojOUPcpIArGQsj2ILpz5hY69y3
7qEblAk/iBva/LxTg+h1E9kut+HgpjpCVRST8HnxDj/gmPpz3OD/I8DyWf4NTAXWYPl+eY0opbiP
qqE8AI92GJCF+9PTqMMtcp+x6Ppw0dVDWO5mHuZMq6F+Ehtl9XXbGctZjgEHfSWYbpHK4r52UDDA
/etLcPsAEVnFonHTaHLPdjYCpTDYi8LrE1RrjqpLRj4yF80WUWgQ1o+rtRc/1KrkEApR/e0G93Z8
ztgoIi4GjdEpsHw+Tbw+q3TURsnrJ+vem3V0HvI6cWxZDGaS8QF0li34b7D+BjOdlbTYPrS8AzbU
9JL1hI0XBkiZVjETffbSoWmuZt/dvwi6DGYqHSnIzC13SUNl2qu+w6NPnodzY2MMP20VRLt1qvmJ
/ZfHdJwomjH0lRJFWLHLRSHa5ooPwJx20kW+JiZ2IddmB4DU8dVdt2qGRHzg4/OJx9uV5BaUCOJ5
DB7+UJtuKssFve9HfSIWDKf8l8WdxwLjopxWCwcIL7iwRKvNjX4CK6tkd7E5wiMRdEELvcgzB0pj
xZ6eF9BMrkKMUgdHqy1GAR/mkWhfFxizsfxQJ74WYCbIAERkE1fb8Z3WXSw3lYh4t9hJs/4MiMfl
Ayjg2+sOrWYv5ZdT9867TT1rcfnNCHmSd58CDmNtdOs/9QtGKusr3RiZLSeBkO7ZJnRubQm1IBqE
1EkkUJqoXGa7Xn47rGGSfL37PKnmwSCJyS1leL3sQs/CEj9vgdEqoX1/oVXfY2tO8/8l3HCvHWu1
6irGR0Oq5hPFvv4JrdxoUahOJ+kEwDvnj5VUqE3YwYI1apIQ/ksWi4IAlxNjETKjtBSMCVjhOSAC
YgI77TF+uv/cz9j1aDqFWUlrFTVchU+WAZW7bhW9jLphCLiSWNxj4xi3S3qQmuZIxCNGjLELKa9m
YS5graPN1ENkiPwRVhAFNAzWvrh2r0Lis/1xU3IMlHMspXRyZh49CoOhgXjEzJYBwZcwV1Y8dHLI
YiHg8xRl1ZNfrV+TQ5nx27esD1wkWcoU3BgfXEqCa6yDL+laVv/SudLRbKjzaC2FOK09OSuKLmxD
y0v3bjjS/MavEL4HCDr2KZv8qcpYRgPYRUc5MuzZqIbdqiCjD9Ty1LXUfs1WJT2A0GjRjOMIyO6R
8UBLVAXN1nY64cR+ylmSfka1MoGdusQMs0dfHuQDuQUPWd+jrOEd58JiAyv+co9y/UR/CyyC1P6Q
zorgF0rs49TU0lyUBOPxDmYj1wCjEe8IJM6YpiD3pfCys4HPvC9nkLuUoAKVpF1/w0hjWhifi5zL
i2760xzhHp5XOTyvydIdQlmbbeg9oSaww53+DPABVDodQb50KxI+ruyW1V+GLfQ8FquUsxNLCY7J
VLfQjf/bn0B0J6zM3oS+BJ2rKvIBx7+iKidXS1Nywch4zrEwfmps3UoSQdxxbJIA0YcYCIdFIGdG
idCrNrR2fNgSOMlI2s8hc4nYKecD57kpMaIneyppD/uZoBr8nGkOKFxs6/ls2lKr4UI4y6mDlqWD
F9OzL+SXX2fbRz9KcXiLNASgBA29nw/n0PFmZ0jbgDu3Dj/xBaVN3McB4C+7+iaPL0ofYQwHy3Qn
615/LFinrmOBq9rlgp+afgIDY+ZkyinO103H8iD8JYlZqOfvYG3jZ0h/dZaLc3sW+tX2Y1juiHFo
tpbn/W/fhY4JZU2AJky01GGFDHPTy5ecPcTsf3Lxoax8w8yzzZi1/LndCHRAorA/lRvYGL3rxohF
DDcQcAqLYCdcuglhOU67OY4zCdRByu+9xwIsvOQCQzRRqt+HTg1lSM4tz/2rhNX5AVbXzsNkmPkx
eqH0+EeNUm82aHDtZ2uWOkXpKxzvf4/XGJmlQVyEYGY+kHSJn6FDbqHMhMuFv6bnsQ+jTwF2XL9P
HOa0gUYwJEhpGlUU5hYBQgw/BmJHVLB33RrLewv0qmqOgGuzrPQNoPRewHds6Pz0Ht0e/yO5HeEf
KX6AFfNnKqPuOtekeXmqxZKjHciMFkwiBOVkMfXx/tG8dT1AzQ06jwr134kswitfsQMpx5CZesD5
rkQeesykbnK9XvicAgicPs0bpWWPpvF1ZmIEBZuQAcxbFiACftsgufGiGEP5TMusW+aW87jgmy8+
EjuRYfWkFASY46j0dkHHZvj/qDMGMGAIwZWA9WXep1sX66dyv0MuqsIoCMwaeXoktAvIJFta35GN
KNtK7d7akKXAJ+8tkD/8puRrhFVMm+4jr0prQY4bpAOolPKr6I9k0HDk01Fmzs4MBkmGp7eqsy0S
gAsCnUiIDOy4ue3pWgmgoAUu9Tqqm7fEsf+PHqUXS4aZQhzS5gQ77nCnfrXYRdXCRfR3XdVElG7g
M0vyTq2xF+KW2KYp9hr2P2A7/mSeBrEHhT7JaZRD7epnBewEN1toeHafMxsbK1xm2UpdJFftOGep
Ao6YissXuqOcC6In41IcsVMNK6CiOHr0MnWGSO7ZHN7m01HxFX5mptD2Od237sPBzGDM1XZT3ewD
kKxwZCZ1mi+8MC2t8sz24VEPAmLtzZifvG53JZh29egKyDFVlHrRZ7lmUl4vqKCR0FMzF3vnwhUp
3asc/ZSDYH9zxpE5lGtVsdMkqfo+F3V4MR9ctz+q3LCbcjLhg24eJ4cvXHyalmHIvXr8wPVZJM7i
TLXeuiGuR8wE4/T+NKBPXdIvBUKlu5wd0w+xt22w68MOP+3vz6s4W5KQMpO7fjaybbgVRCeLynhU
Vz6curg4Exv6PDQ07Jirv4EqdebwSry9i3RUJ8Iq+GKy0GyjHsUcpTy3X1LT35GIenGXfDN4ruNd
M8BFnevtKn2BQ4cdrddLAwFJFSMFJMbgFWGZjiPkkDgk4FGTFeddzAJU0AkcheClvyQ841zPxckC
9zHy4en+vFNKsxtfqgsm8hA1pzWrUo5ec6ZtUnJfiNIPe8oudwGN98MXgbfp6peGTv2Qm9vQmftD
llCOWMjWzEnxHLADL9j7K0lLVq60RLQblgoEsif0DEOncdABVET9x+I+LDy9ah/YKKpt6178C+rS
4+4hHLdpe4T7qYjK/waCo95go4IRqFXVt1FK04TXM0oSGw3n8faFQ8nxXd1gLECX62mas0t1VY3E
ZahxZTuTQHxmT7hOZNXzlampEc9Bsifyc310HpCghnXnWSfmh8BH/BEuLEjqEs7nL5WA1hXWq8p2
Xyb1dkn9SYuRMzyiyimRsIrpioFcutVUB+wcsUk586fqIe8ko71O12K6uXNmnPeuB8uqBuiWb5n9
vitOeFONEiYpJJA0xnE1fJ6e6yW4enI3t+63XeWsSjm1+xqZFGRbfFP6SLl93w7cX50lcN3fyvrT
GSnvN/KRt1R6+iH5b3+8yYmB8WmjBbGVJwzeTiIk0XCd+3hewDhvrpc1u8ra9G+pmIjLcLUWFsYF
LBuQS2abMLXshzWf1enknWN/rXCN9O64622IKWwEVCt24/CZgV2rrXkkCJkFnD2H81Pn5ZkdvnVl
+F3xKdY9PQ74pdnIGyPiBnH+QFPJY6/nJmb6na6eVH5kocTctWUm8npTVajEbBhFj1eUGENQVS6o
Dq8UsNAyrTjzwnKon05raC9AJv9N1xDO46qvOwGu2YsE98CRPdLPpurlbMMBI1IHvcB47VCt0xDE
nz+JY1RIJVfxae2gQ9JJXKuORpFg0MiieuOt1R65RDQmbA3V4hKGrxaFmM2KH8ro4Z3OclG5WUV8
46REfmTYZ1x747tz+hGelFIlwXmc/WSO9vFE9yCw5hj76UixJs6Xf18ickcex4k1sMw4Qc23026E
GFKsunDfWi7/Cz39/0bN2XZ0qjjlGnPA3xtRQetell35VnUWEF4ZmB/iALw6FenfyL7YTIP3r0ik
d7Hx19u4c9ha0mwYR2rqX44G8Bg0DSa+3wpPvANJuIe+mft/7a5nswMRAE3i3PNSE6K6G4gty01l
rWIHavJ8Ua12uZ7zNro0g8Bp93O3owMngK/cqoNTM5A8Kmg9fLmEnXp7pXRzUxhKConWC9M7nOaN
n5rebRKx8u78+yl6mqqyDLhDLUqckSKxpcCMzOUfTiyibJ7eyAdDM9I9m7kjow6xFd1wbD99tqVc
il5SRIaLRMCEKFgizQgFMcZmxyHWDZxos+pgFjX1bGjmgvKvyym4gMSpu7GSZmX1I/Hpd6ZGw1Kw
xJ6rNvLb2ONSNfHhtwQ94gJIsiEBYqx50Hg4iYJYNMXa2et0UjfvJeThkdRx99FkS/FSW5yvmT8o
lIIevs3b8ZrXiBctMqX2Wa4gYggZnE32VKYBJuddArXrYODCqrPV+HSi5k/AQnRBhuMN24QVxu/M
SH5ONm6vE1qRu1LSeR1WesKqzCM8WtO3Ihe2mnCnVnRCvOewgQ48QlNPfzH74RLcBUNy91zoslom
1yrXGuLCUkWXETAblXWjDA2bX9Fsc2SGB5rSeBrj6aMzuWG31NuVErYrYoNItQFkXnUZMmFZjNvw
ysU9IG74W82Qcj4JATnGBt1cXvFA8z9iSMYo4rZzNRu1BaC3EFSaFa3iJffIF/zQoBEm1ESxA9yl
rvRoVIesOSG1fGdpD3dsf/CR5c1s6xqlZfYIvd/HPRN2LfaSIasLuaiRa4/jIlFDR+ICtLWfZWVr
LNkTjYgGWigcXFgoItqMQSnQ5xiMElthXh/f/mfLjGsLu3QDP/y8wpR1m+B09QStT0HkGeTtvIuV
OW4vtf0KZtXPa0y1tKEqJTSvz3vmLe32PqKTy7U9Y32LoPiaTDjKIm9/OEFKm1vK9ux3A19j4QjY
d2KiuyOvzbW9R75eREcnaOBuFpTvb9W9CwCQaspaQr3nM0vr5QkYVZdPrNP4ngmHt/dUVKz2DtBF
4CL0zBMJahnVJE5g5kC6FfZHVJYkBCFcuhqzwtgfNEMoPB3Gzu5Q6zblbmOA0y5HfrJZfscNTnle
QsMMw1Vor/eEVSkw6oq5+O42xyc4yazTvG1zqiLupw60HWp2Znye6e4K7HYfvjGGtx5EcTEPD7Wu
o+LiXF+lDjF2KPLhLu33N84y5Kdxz43cISXWXepTuzYjbjDzAYvb8uRV0HkHqivoCLS80iKz2fJ6
ygCnvCelu5cD3hXHnN0AG2IzjcYF7JzdIljBJgDYSBvbAwZRJ+HCLl2ST9nI6liGY1emoCe3b2Ar
nFJlKStJGOoZ94RpB4HDrOS3i/h6lx71tg838t7WdLyr3GwbAEWHR5BKPIs1b42EcKpi/2oayrvE
8W3/CSJdyyPGwMRNJ/3sTa58FMni2Hz/MQSyfeuNJVM68FstsMibASgRzwgQI4MT3O9fHueIRnQq
K/nPw5OC89BWTX1Y1hTARt2N65kPHLFCRuLde6LAqO9wjbUs8stvgw/Rbqh5DsFT/dHgazpx66SG
hgKPfHqwwN7L4x2NOGA0TGlQ8KPvGb2wZEgwuMKEM4mnjadk3Yyeqi7UaKWFLOzkapZEFN5WNoKm
/9/AWe2JI8cu4N0qj/UwET/iQCsNGhZ+4E0cFIJ6bKYjILqRbYVfQ2x40jiCHkjECmPKoBrB6DID
2X9vVaWStRdX2xjudw4RDmGciSHH0X1HCHuPn+JThJr+gEEU5wwPupHLzxPhSoDrVv/I/fkmPDVa
W81zqxsgtOVtwYkHYJle8R07+fRdlLDIBnfS0/Vv6QmrVGHr0+Y7R/kPoV1XdD8+bbU3RXq6jDLB
2s88LhAgzrgNKRc0rL4rtAQj0T7zwnO81qg/Njay11zSVwPdZ39f6MnegpXb4cfydfmAzHFNXkTA
51h0VKUh0+Gn4ODWQ+nkcwjuvEqoI1RbWypSvlDG5srb5LR5+NEUyNS0lyZ6qSYdhDc6FbkkmT7Q
9ScVJ9HwoKJQ4uniujMow+g888a5H6hy90xZtxXr1Shi0d85nziDH8UstNO0cjGlVDWs7DUm2p86
8UNAz2L6yfrPwKxLbgvYXyiq6MrUkmMdR65d/QtJMdLDF3Phm+blTPIRvGGfh6m/jl7I5fw3SLP5
3oROefTrEQGYnG4NIBiCTBgeOJkP9SBMRnMLiGCZoTvZHGQsDGKJd+6tucDF+i0ooHdEfy3bdbbQ
8S+ofpMJ25w2noZ3JLI9urDq5GLzdsrJqNrkQkXWWJ4Cy9qc+cEJcZa0qvvsYlhewnQ5PVEXlMCy
KetGqBvpRyD4Rvm4RAe/kChPdqNm728cAoyn7FH3RwIML1bmWuDUWOMEF3VGIH37m371iy0D0B4F
PsGWHcTLhednAtimrI7+BPWmVuCSw+ov6WZAcSG62dinUHWS4zuHsX4xnJ0AX7Ooji0XhThEdHXf
0uQJVxrFvwhpF2RL3oHz/dmOoTVvU3eUuYbn1BhaWTn3/sghsenWrgROzjUBT4cpBcht06zVuWS9
1JZr2d1fS0vb7NQ4c1vtm61JkoeYi0rzLnnCsfHEPzZBXaI5rIGxCdUN8pOz1Vo6r3/P6ZuMxBzf
8liaFDNmQ+EAQrjc4b+5sSRKU9kgU5Bh+mSGSBpuQyONQ/gKVZubBbotTRFlNhZOD9T9dyiCOKj9
jXg7NI1A5l0MUcHn0cMMcBPenSm/yDvz9DmwxG3Df4ydkEncwNh5Uw7iXLTkphFPrbOUuTvAnE3/
0rj2d5FS0NEb2AEQ+LDJ5b4k9fZSM/PCMk9GfXUiNqPtsvX+qVxObmMXrgn9RKLH2MbnvyP5s9bg
6LN2X4qM6ZQE3KApfwxEJLBxScHoacr3fTXeKWDanL0gf4YmZS2sF49QTrT4GGj8e2f5AN57cC6z
hOru822UzDHR5OjbmaLTRcfiIK/p2X1X8oYyC0zqD/PDCKPWighhaYthon/yG1yzM6xYu45gDqwa
5zu98GDZ41LbyOJlQ4JE9g53/oQxAnmsOR5xTv/6tMHUBtm52EMDBiCsIGvpomzbcnx2LHaozgnE
iHb6rEaz+hnIuuLphxQFKu3+E8cHAtBXgl/N3Ko0XbflhDt1kpv/MGdse/A+zpTQrfvNRBC5hnhg
93MbbeUL7WVqAeVimyJBtkeBNDSO/ljCUwMLGNmFYcZl233K6d61+91vUubzo1KRPMvQLhPkhADc
3JER60r4y3IaJp5d+Xgd/gtPO8sm0yENqyCZGdm2OYBa59ncjOkllcDderSTO8OEQ2d2foCtQGSd
XUIhcxDMV9O9dQpa/WXGoEgQLUgsXftWapApjYykkCtr7CeHf3f4tzi+JKLIxkSr5gno2aXGPYMV
AyCIUB5uNSBJRGm2zLRuk4WKU00V+ujuErWgAO5qBdmstZii3NiuhCv0Vi9NVof5W+cKFKEvc6pu
v98XbNo9q0n0GiSUaqpq82BWXOSP7lOcDyUmRLKMI/zd7J/Bt80gEXli7Bm7awzzLUnA6Xra7MrR
z6LwdLcoOvBvnIPSqde1BW9efHUrC+soolalTnKKZaXU5ZS9DaJz5rlYVSz4qFzVfmV80cP8KGnq
XO1Hmv2QXyVhVwhGplJrdpC5MFzLX1yxOsrh0aPFwAsVFDYdIyFbdV160LedrZFjEOk4iJKind60
yoFSqRHUe+xLNSaLzXfmmcnHFUpcndlf2VG7oevUE+g4+Qt/IvhommzmRPixwLpCIYV2hxhsn02q
Jk7zZAkZsfA9PI9eEwFrj+IBehhNtDGP5Copj2DX7o6hQfmLT2j2QdGLR1ccSnjZy8Y65LRDHRSi
uwVYmC/m30EOZmOBQCHfSWNr0T2iR8PBp7oob3QlHAgX3jsLxpYLurHYReJ/2l5/dwCBM/9SLMme
Ct/gZGJYwgl8cvmnPNv8DgkKFERjqsed3go9MQx4jVC94Z8p4FTTIPrzi1pOj54L3Uf6jqeTW5qb
vm8JLvcSyseOtjKoI113YvWJCrJ5Xq7Rs4qXvhtix8oLsHltBAuT6LkaINQ34QNqcn1E8UVbCEEC
6mMltTJoAPnIgWXjLPFNyWROu6BMLA/r9VRkkKtZK3kglzdp4Mt0iDF/ZDlr2oSvfhTq3OjuDQzm
QEwRVdyaeSHNT3ptZCC3QcGY3WDIc4XeymOo+V3m/YIZrXqeuHlkam1nm8QOMGQlJnMIB/f7xSap
WXmcqDfuKbMn2Gq/YOxX8bi4AOKG/0gh1CMW/IIFaSqiDq40KQc6jpL41PsmBxho7ShHpLhjzq3o
IBgxkkDHanpA64wC+VEBiQdRtL411oE5UywTdOpI27mYgS3jdXgujKZL4RIZcS9MJoVAiDr27hf/
gvrYanWs+EhBqsoJ/xLz0LCdzSS4LtwQBGOjfmBu0tIATSE2ifegSXgNKRUGixE17+/p1bJO444S
Uegyq/ZOfy7MOUvqwiBCZJaBNeEzwv7ejCpFMVHc0OLe5JZ3GHO5QhzDJ6fOzGlts3TyLMYHs065
4UidZAKrOiRXbuAUN7qVLWmsnipacgv+lYLcExk60Eat15oLW/13jip8e+ah1JdPkyvFugU1+X76
1c8p4IAE6Kw8yr4s0av6KwTyGM7ELcde88uuFw27ol8iifl+QmBVrBAeoK0tWF+MS1nC1jy9m6F5
hh6orJKSwpF4Fg5J8xq53qwVkfUNARcOgyrIHnsfhw5Fh72igyyrQzYeeEnKETyPrC++R92pQrDx
eeN03HUe2DgdDkboqbHrL/lGfLyJbKom91gZKVXIm6BTCm9FtH9Yjde4m+LmotPeZxmIQCb+haSo
GiOXbgaWXc9XVlM9KlUZm7Pj8vC5rvwvy0NyVSB8ephOQhgGz4A8V4gIoXjWnH9lDJoWdGRS2A5E
DYbRIhSi0F1Ocwk2ze17cs7tMjyB7O2bVPqi3wOnxwUkMuH+yBZ82SMwrJBrxp5k7mOjMMRsdrtK
9lgwhiEtOSXWj3GxhZmB4A51/8CSGGLKdFSosLwgwi+Dh7uIhUIrrphiz7xLr3VUrkFfC2n5F5qm
nUtpyeUlwRNrw78g7yCNfyj8F4gSE6+TDFb53639MGwUjf8agSr9j7kCEsA9o3txrgwD2k+cYlzB
PKEt5eb3f+SpiHRwFee0cC1nDz3WhHuyXye0NZWWha0yE9Bc+pwYMrs/06r1wcPvpj03HmSklpqk
y9I2cW1fOEncKzGtCpRP0ciz+GKcSk9shCh/fbYqasaX5k9qClRAZ1j1tRq7K4PTKQMg8BhZJNVV
PxWfbwwKibP/wny2WuvHE6eL4V2dogkA04WTnJZZe/xEAJiNnwdwIi3jwxgh+9yY5/By6Fey8kMr
9M+lIt9bHjijpN3vIAPbvnBbI5yfl580Cv71q4qO8ZvnLPWCVw+zX1MlEbHAzZk8Z8khd6JOte7T
/TcIAJgTPN4wspMKbiW+MA8LXOx5NHQmIOAnPZ+dR/GxqoTj2XTWI7h+D/f1uGK/RgDAp7zJwTkW
OWbxN1xAbc7UGILEqC0m/l+DmXBfll2HmjkTywmpJiuDpQufPnhgtdDxy6Mdx9J5WML/eHPi7xGP
TbGgTIZ0qLgT2j0ZIgeRxZBaztiP8PFENAbM97BYRyMRGuz3mozGwdunMn//OLCdIgsStCTCFsiq
gdUmYCj8+TuElfCwTM7D72yTIe/u6hoz2TsaXiWfYz3p6ExLRm/LV2y/rRmNYrNlEdEanv4yA1sQ
lnf3dzw8itbPdJjoH+F7m8Xn6K9DnkgW7pJn7mapz/sUR1EcLAU/JAHuUdUvycP0e6f1iOezgxlJ
zvGI+FW7mK70UD+x+YZ4+fdX/o6uyL9k0THS1GUcyVQYRM/4uCVzeCocYE5R7UVJzC9/D3q7XTVh
raK0z5DA3YzwP6yDPjUmN/uqb/m4/hLnyIrTC03RNthdXkVDpenE06yHUl5nL1YF2m+NTjSDx8jL
NwJ7vutoN1fmdKsMoxE3qTvgT+h/H3uh+PpuPvlgF0UbRLKUC1+RwbkFAMIPtbgKheKiQpaTCxiv
A3bNx1e+Fivt7nr8yCPS5VAOIacUHTaX+SuCQpYMPqy5ZPqR/H2Q334kn7prJ3O3MRYaKENCThDq
CS3Q6b3X6ySSQgzOBrIczNBuNr6L9qVh3XumA51ELoTkSd5MeMwZPqa/nRoOfpVY1MA1nf0dYQrw
VW4XYFlB2eunXujLIbgb/xRTSTuUwLBD3f+4F56QABViyR+zX/xDoP/EwgJMFrIMKkYDANoQBa3Y
I5YhHepJW/HZ2HggKh4MSFmpvsH1GQYPYDPuhi2zK4OuXF5fV77M36jp6Xyb51azl9nFcIwDhKr0
lIWSISwhGgFrjGyE7pFbpGZjdm5BTN/DB1qJPyh5gWoebu0aYrn9AcR9XfizrgJwDZe7PP3ewW6w
nGzs/WK3tQvvssmiBSiSCsg5FM5AFW4Wr3nkTA/hAEmz+GAw7y9x2OG1+tdT5uXSVlvdiRqf5ZqN
BDReDtvzGuDN/4TkVwb3Bb0qan5dTKZ+JNZXD+wViDgJ6CGeeQUkV21ZqxRIWfRt4gym8MXXg+LU
OZhROk2KKaMGq1noeG1lCx48xejSidMrfwxuPhDf6JII/BtVYJFsiolnTG/WzNB6lpoKgysVjZRn
9EYOY9XU3hST1xC8jDL9AlHzyAhcy9lXZz8HgM/EswuZd2Pp6pxxuO2B8vcMUQdGoKfDyaOQ13hR
xMjjLdwvs7Y1nc+IwyWjjl2MCc8R9PjLhVCMX6lOzKfPBxXwc8QUib22Z4UmQCuIXU0GJ1VKTBeM
YyzxPvyC6xAJuiPs0SIxeSXibx12zYmnEBPQEOvty2Wmv1xNP/7ocIgt2UItnuSxPlpPfTjkazKU
BF6HbE7YEM5is5zFTWxxy53cPkntOfXsjTV0/Wu7CgrIiuNbhMfkSJsFH55nRt1RgrPGP1+wUdD1
bAoMwSE20tKYzY7K7IN0q9RwKli1qXLwSHdafbzbDyJsd6T0hH9lZlIWNJV3ph/0MoCMkkJru5Ym
N1d8ukxPyC00xIfiiiHYr9dA8XU9IjhWXzhjE2Zi4c45OLhxYNGwLujHmAccFDsSPixIFmAM7RDq
OdaVzQZbA8n8P3b7YCtWqg9bHqOubWvfCuiIj7/9pr7hxe8u/L8rUhYmExwWtIHyPc5sKHQFcVSC
oXoydUI9f/EJDCqQKWdw8oG79XUPehbGINXBXTLqolvaSmra1TAlDqH1J4lAURoVmN7r1mYsbzRd
Z83u4OgLkRC4QJBHYbIj2coJtnvkY2zSCmPzxiv27AyZ8eho9Jheqxfaa5MKuTZJxCU2gDT3GqD0
wDAe0N5kRpgvvsdQGi+N0cQkwqYUJIhoyrYBGfteTl0kxPa7rkwiiv+UFZp8Il7HszCV+hLlkM9m
plyjbDy47CvgpDRR5Cl5dL8V9xBqkS3thX+LYZ/C8RUlKSWKOC/zBPJmfU67I47tILU702MWoClJ
5QZCkGU5lKXp0corngICW6bqi1L4YQOlfzPzIzdrTvTMoxNEhF8dTeoqltFJgVjx16avmOp9liFW
01umz/tuVddsatP7ugyhlutqpDx05Pfa2kYZizAivqq8HgPD3B++lvWL+rVNhdfGn3bSmJt0o8gR
kuh6A/VxzhONXCPlyKuXxowZhtLmkPuuvrFKoiKGvYKQOqDJ17LlU5Aqg5qymJNyehazPO5G06/W
u2d3OBOUq29pIOn1yts5nGG/tyRVMK4lp/WEWG9nKEhvs4yzaKqXKbe5f6T+vSxRRUQ1iWGZNH5d
68cgzFHFz7+WVbs3OlcFGZZmqBhL7Fj0jXlOFiK4necRK+nB4vtXr2CiiDXyrzhDuaMkZ3bIDLR8
TAfHNUYqfO87T9YoiztVIuH19EGlKBbwG73fEk9Nd4ZploF9qwOBsLkvaWTPvuEbiC3otsGrcLFp
Gcp1KYpiEpZTzNeOsKOZUU2tIZkH57MmxayryLMwcS3YbKE4jiulBhHkqXdKzxuqIDaCFvqMOIyC
duiU8LAlSBfMFyC3IHRCySzZj1e93ml7zNrSYpcgAigStVT0LlDJSUKxkN8JU0GvemlEBAC9nJC+
WOtRaElsOVx4uH5ZT7EzEUHDg1RYKAulX5E8+dyMBS2g2Q7OjijAekWFC8c8XCTVgHHix3Gj6Q4N
e+locV0HsQ7NGBpk3sgW7EG9NkRruA4StMUSRkVhTDJIEl+lQx29th9mpO29rugsIyTvrJtGuRJ1
NSqExzxM/hb9VIwLfVf+XLwDpDY+qylNBjjegQySHRuJImZZyZhyPaTS5TwpY/Fwp8uNDMuEwKOr
+b4gg20B3Q2FDKallP/j14kO2IaiHWIjuXaciak9xtTUqMuVkQfp7mGR4JYDC8KLrWYKVGmi8LMc
DwLuVGDomV+ggE5cz4Q111jlMwrEGrCIFLFsMOyO7e97g3GTBn8hR3NshanQxvl48j2UEtMRQAQo
zblBAPg37Q3lFIIVwgVWqySYM2eoveXP4A9S5XyznD5+aydWMMWhNhlEXbH+dyIM6+T4pW8jX6Ue
LMg2N6XmoZvfqXe5nCfCHo9taElWX99OocbHbzADMl+lBjo11nyW7Lx5g9/Ro9Ko4PDLmtzI0OXt
lx5gYjsV7F7EJiJhPlFdakImlazz257qeQ40DqYMMwvNhU9BspGbLVpSn5ctnw7FzfS+yaIycyNd
6hecnwX3vn8ZEmey1oa96T0MPxLI3XwRfQj2j/9Lgl6xhLO2UAkQW60Rpv5ZWeA9+AiETLRbYwaQ
GkTcXXYo4gL9Ets1B7k1OiibiGTP3qYP+HRY0QLlLm+hWGMgW7OvUWBim6GIAkYS83IL8rP6pEsc
NirlwgbDo1l+s/PLL2eSraM2AO6sgBF9jarwIuHN2antPK5nXpJGDsy4ORm2N/krX+FynPP1aKIe
2zx7mI4uEDBBt3Zx6VuzJwS/SbTlUJOmt6mujmJZWbwPvKKMaoWTy0QYeRGfpoKHLllNiZkQscSz
AcEwgTDcTZoEq+CdFrC2DMMbNkM5v2VqxFAcUKR6mY4yIaYtGJ0WLN/hRHTWNvQ+RVWCsmdVaPbj
JrxV2n3JtmOv23NOxeQZhqxZVfImOZYIAQdTcoR60LpqFNsKWyVGUU7YCBkfrDFl4PYoEEnIoQr4
dScPU0K/IRzbKNjbuqdCdvLtghBmV9MobodEzfD1yc4rtH1/A40Ygs343tNYg17Vcfkofxkf3YJ8
Stnlfy/47wbTIp10YuerYV0oggsMFN3fBNT1yEGHzQuVGlfkBJGHQ/U9zWG3LLObXhTu/zVaICTv
B4eUh/q9TAmzQrwUQ7AkI1r+D6KxT9NvVoDuhblCUy1zVrfrSyFN6xtvpODmi68zKtj87csWN95P
wl5n12A2J9DlHc8Tmkt5OI+xRtFbG/i06qJo1t0G5ApSBc3OfoUZGsCt/NC1DE3qzlKqP0TnZVNc
1SnO3+me4MZFkDJerY3o0ajCx8b8uI+8fIdkWcPfKRZP3BJoIiGU3POV7HJVGpCvkSug+drAmnvO
VmFQ9yTdl/mXv+6mrLwIPH5CrU7t+i6w7RAZUTHJoZo8wgY3CZ2+osvBH/7mUeP2kyfStnkY4/vJ
LkCFAwSDdjH3qemyj2PMUT+BKSe+jHgTLKznq17ktBLzr2B8tHeVJSsLV7uawLJzyJCRWAfPkKRI
w0g4FnA8Ah+xa5/at/Doleg+RkBH+wqR3rFPiiBG1ZkDssC3Qxj7uDsBUDqmjM4oR4wCI8JdqjvR
nf+VK66U6TcXmYwFPrwY8+SeUIaEpV7tv7/Ay5SxG0U8SRJwhr7TDeLgfLGLOKobft93aQYun6AY
2/8ByIOsMRlLhPqkfGuD3nSR4nqwJ35rMoPzULX0zs34hzcUt3AJiJN4qh1XcpMUi2B2vtrdrsdV
ibyWa1l3XLWAGmSNxLKEseID5o5MNT01Gr1LU1hdHIVvAyiwA3eN6oL2tsM4SDBy+WDJxuh60KcG
dCsqdbhHhm1I6uIXbZnaV6fGcnBX0VJQRixRrME5hygfNnu8TKUcuFb7cSW5eXScicgraM9sTwK6
G0jfEe0+GdyXK2DMSGvV61yTK2khk18PBHaUDjt/11FAt6PSPYz7Kfx8Mbh/OtKQusQi9MVWF3X3
QYW334eP+7g9qHsT2xdkvpcfH5DJmrkDodf4Q6ld1cXJLcE+WZrJpOcXxn4bdHaLy0kBSKMIYO6j
3skQbJN6Nw/Z6NLP0WfTjzFvqoON++4tk5eKBn/uSGUZvLzaQmCWFSG1Me410DVjPgwFL5+kldm+
88YM334sNq93DuNHvl4NDitDf301EyujUcfbnLUga1H7HEjoEwL6+H4KoMpQw+UrQG/CCAqQsaaR
mMFcmx8NqGNK5cZCDs63MChuy0Qc9T7aJ1GQIyVbRg2TGki8RjytFRHumCGiOgAXo/B4xBtzCzvt
slJ7KcCId8/VIMAkmAWQC/8+lOewbofzThvMGOHDl8vDMlRSRK1rxYRBgrRSkMT3IbQgtQTsYN2a
31RTslmFS0EqD7GszE52Vu4QV7wBrINTYbIZGlgp9UXt+VHvONum+WSy66lVm2HJrTQFc1GvsoYv
k0sM9nybzgh3msBf+M+9lsrEiB8gIpXs2/4XfnuW9HEjM6w9FJb2BpeTrDxJujfmGnvVUj0xd373
Ia2kyXICgh7y/5jkI/H9reToL2bOGSlUqbeH8kNRgmxiRbdpTXMnWCpZmxTZbq61osIiViPjFTgR
Xa2VyfwiuJHk3pqvgFMpiNEEqkxsPTBzUimZCl+5PzKISXNVP0/q7Fu2J+PFJcFBIcS/H/80/4Sf
hV3XvtSVB39z4iNBOejqIJOuOTqWMro/EQ5BD6q6WjTffDuMp24OdZH7rwAoERg+GnjLOCF8H4xP
MKRqie5AF6goVwQjiPLGAiW4R6zZyo8XLNDtMmsO4TqRCq9ViMh7Z1tdrvkeRWw7HCaBZcFcXsp6
+i4SJYhWz6w4cCFl7/mxebsgAaAxi+ZqPR4B0qYp+V1W0r46hFgEMTdqRHwV4RNTdXaZ5CsfHJGt
z1/8hD0Z+i7i5RfVsluLI5aYx3eV+k6XYT2rrH83brpXrdnTcVM8ucozx/oVSNyqU+CuoVJ5SKi4
gEBvHPRuuHsG9VoaqvHPiSpGfY+hePY+f5CTLlt8t70G4rG/uXhKqtNaH4SV96YWM0d+DJnNcqby
Es4FyAHr4HuxufkihcI3b+TaTN2AQLejoRGOpdd75oX0Or4SYrxAWRIKH3hajU5leHMs6HJhUPkG
AroDogSwoVed7VHNZtCtssa2ullpl3Zt+ASvNnnnJ7CfMth1tYJFYYcZ941H24WsV13bjc3wie1r
TJ/53Cyytyt8SuJj2OXZ9NZQpzoPDjE5A3l8zgxw7rOP8Z/Q2GPtKFGVJVfNOkXWk4QY7htCosS1
YKo3rSB5FTlx5GMt0Ef54mfiYJt2pgeaVduvNE3olSowcnYVaYjDiahxLo9mbzxuum9JET79kYYS
yYMMF8GBIsVyHX7jRkf8gH9A33BsJjC6XYH+78/MSlXhiVc2qaEF5F+wdSSIbfSv9PhP1pkQxVsR
hzYhGH9W99VknbECat/gbPQxtzdirjWOljjfq8cn//aF6WmTZdcz2qg3YVRCL+Cn1w/QrLipVCch
We9DGbs5bdzEziLFOW+ntjh5/iKAZpgJs/jSmBJmbeR7sh2un3DejlZaAy9aerQQ4BrJ+ceXrQaS
XOoFrHYd0XsBujGNqcaDPwcbRNL62Wbr7n+CsWZ84P0TR4TTi2IU0eGtxF2Tp4xiU00Ls46XZBVG
gr0s9RUwjbIpjoONeEjPDUuV0/G/9haI6AofCuK5GNTwWTy87xgjdaeKYH62yLfsu4Girmit/IZf
rPDpn2ncPK8l+llyrKK4sClW7dQWFF43/2Zx9eC8L8viRyOneJVHmMgvdll9uNX0CuTx66zsL3DB
qhu0OGnrD2rK1G8kSw9rkLpAfVlCzjpobfPm2DtNlJLrbneT82pIDy723mayVW5niXTySC6viGu/
B2MLVE4ovuZP5+UTKBD5fOufR3sJqFjaEfn10Q5hkAO5P8usfz0OCT2fRQC0N1rH5DUjbO1RigOa
sH6dT0OKP9caLkmTEMasLK1HgMCpG0f3kKBpX52dk5bGvVz02tebj+aGx8J9zLqotWab3mOYIRHp
PWXkQiQzjHHbWoPYRrIAo+qLqEQ76da+frqRFp48cCC+hhRaWeqzEkMWIJeTYbjH9VRsWOKZ9IK4
L5VqwxYzD089M83p193rqhyD7K3Fg9XrDyRg8Vx/IbFV+i+F0RZsKwy6w2jWZwlFGBLOLZQjTBIo
IENY0eb633GyLpWLzfzrHAfyK8ZvowtFTWwACJ9RwTldeNrXNgTIHd81jV0FUYOCtRjVRxzEFZUR
FXdgjooRhGagQWtkbKqMuKaBPkZYD+oEoVjgNEUVeIjzzj0yd0cKwhVMu4zsTU3dR3PBOg7MWGvu
z2o/q+qerDlYPDOVmJ9p9z2DGw9iVVb4omeFK6trcqY9/SnAHhk1oS2lnuioO7hg6bUvvdXe4XSA
Ca+O4482jW30WTGtsGIXftFvXCDqVX+gVSedLH/ZnL1abcZlopsU5u64wvpfiV/uu+ibno5E02n1
B8ax38hzwyM0QE2NOimTVKkZ13EukdOKD/BBV68bviSzkCZUguDCr51W5Qu2mxPE17QPKZsy0WHN
pEgiylGP4opx5LeFh/towxaQKNWeReWPm9ewPUKnAttlRFLFOyhkAZqTLmHp7k+j+sKynmFBfIfs
zUyFw1hYuRSQkfMI7DvAvNDLcAX2LBXPvjAHZhGnoKrvDt2Mz/Gzcp0+ywKOU9qUhxsFUGoVDRU+
IAG9OO5H5y6SYcNbwt6pusKRMBzdjV7L3YpiR+eHVCeFd3BQGwRhO5US9V+iVDpbY0i/hjQ09iuz
l/w362tkxP/KqyJdl9SSRdVcaWDas0XeWgBCIK8axj5n9+cQPJjYeMR9+vUuwg53gGrA6iRKpEpy
cg0qu2sfGoTqPBCJx3BUbUeiNetg1SkMHIi97q+U2+1oGcjKSNCAM3n7/4c2TLfvK9Ed4Dz6r43a
hqBZj9lHch/ZYT4F7BkRC/FYm4wfyj27jlN+BW95oYsFcLrFmO8F4DH3Yg05UTVA8VZSNvrsHR4O
FUaoEn/QZ8SlFtRiHwjvw8GAp0X5NqTuMADloK26fIJQ9IxBSAZvxD42tx2FLZfDXlnxsYH6j3V6
tLEQ34Ay1V1pkVFWN4DKjLJTQTcH+NGEBE+uhTiqwLorrE3EIUyTCi3em12uC++VOhKqnQcaF+YV
Vg6PF/U3k2BP/Yk2/tAaYpSqCVYhW0v/5uAfa7SdoUzNW2CPMdCStXHi3oYx9nX5m2PaMb5Nmlch
szPByVANIfjFCkmwt0VL83t7Ge9xSXYMMpA2zKBZsYxc95ymcUEXZnDztlm+yIjPVd6t0aP1NVPB
OfmFxIE7zISnjelzTjuIxvQyckqy+SFXMNykug7pAyL/IBto1THksupsBkBrswaDY0NjUHP9DDUJ
7WrdMVkw/T73XAVkzfBxPwbiaD6qXYX6ytAHuXOJqCTMmKLXFWf0PvF3JTo8ErslBW8/tiY1xzHp
qAD+cIGBy4tYAGRjNwnvNhnQuGP1AZDw82itHwR6Wc+LHirXe+ITH34yxdQQIr+vGltLDeFfEcvn
ZiX58XwXgcCmj8VhnMHojue/BJ3Jt/GN8BBkZ7qC9OTW7bJ6/Ybz+OthIeq6kWviay5kcX1amQxx
cFzy1AATL/5SIoqDb+1405mqMOGi+NsuQci305vrzhfAwUmWzzvk6Wb6DFXlReWymSkX4khsvzD1
JolPjTFs/eNJSiwPexd0dc029mRgibdZ2zlv+2zKMgCjcQ3zDiXG9WP3QQvlXqzc4TqbdlqK47GV
JuwJmwXFqdRVr5tuKHDLiK73Z0+ITx2ThntbhFJQfBSgtr+0PeB+nddqywWBiae4ihZD94xyaePo
2VGs5VyeupOHS6U/DvlYkfA0WgJr3Q9yZT+5k3+ofTvOBXdK8Hl5rx0+UDYYs/4gj8feWcdPVJno
Xx4yVdKVnL4nkW024ZHBaCXGLHTH53zBmoBOlLh7T4FKeAMup/vE0WfMFx6APigT+nIexMIk6rRv
c0+OqsfWv9Uwkr0fd59qJi0hsM3M8azLNa9mdgYz01Dj9rS201gkHLzMDHiIvK446tqLGGP+AXG2
nr4fx6IJSr43kJ9d7DsPTU56d/Hl8+4xJlkKHgy1jp86xV2xxuAxJxTuKuJ4K+8/PZOVO88se7WU
7mQo8udF6xN+vNITlSEEtTnLrJqf5PQT2I0n5d+Nsm1PhV9VHPWfzvmWltsmg/xznH5vfi55kUT2
tqmJnjtagLoDeD3imWVSAQKfQqsmsxsrcYl1UVC8/nfW3+F4x4K6fNgZR+wvbK+ARVVRWjWwTLiQ
xmI3vTUaqvxSCe+MNLHno9m0rjivRQfCsQIF6TeXJx0kpqt1N+KVKHwge+cJRY3j4WUJe0QNEU61
k3Dl5Ar4qPj4kFHePcMfLXA2IHtVzzuUt8ki0pNY5pT9PG1ChT8yLyPG/dQdfvgbjLK/il3Avfq8
rlIHbIdhZCyLKdar7ZkKY/orp4Albg3eRHFTMCVmiSs4peCTHjWkXfQBEmkB/3w+isgXh7y4yLMF
UMLEdV3Zd6Q9V1+TcHs2VIYYTwfTxGac4UAzZmQdOu6sRCe00bu9FIXrqF2BJrhIPhmTAtjY2ndY
0TgVEgExY6cOqLFfkIYdz8M2DxR+CuwYlR2xX99gf/AYJgeNT/tZqjCQ2gC5C2IIMU41XdzDNEV5
89khgQSq8jkmm5+0z8fSimLGIJWBrU6rBE3x/bd7b8htykxaSplE6eHxsBTvq34fHOrg+ZwjGbi/
dMqooSeDLvzDrwzgiSEbpwKUPFRcOYJCrahxjia3Wv48oxglpmbOLHFcZTiQnM70YcTj3mhfgxsz
ATaDo1Tg2sm0A52YcgufTHu6Upllwr4I/lUsjT1DHDSJFoxqnB90BYSNxR93Fbyl43s1p/5TCZK/
GR7i6ezU2+CLhjZpO6HXwFQnuvl4u2p4KHMw8SA77TyKPf+ys64XqXMXYmB8EeD08dByQqMQjdke
yKy9ACRPOPtmwBLaFY1NjrqW/WJ4frxITF5rHD6SKtKt7da6sOA9g6AmejlD14kjSglGCYeuOq+m
G7fgA5/a1Vco6iUGk5HTm7JJsydnJHKXRCJYi8dt6HkMnCT0eN1IiMDvZEgifZm7aJLxIqRzIRYn
MkJPhDRnfMiKbeYjzxrx5p+UGgL/ZrvbcGiBYAZemNR4vUehhYxd/0SwdC7SXu9mqKFGFzjq5IdV
Q6EkDtERRYMSfgne+kHhK08lY2DciRzQmiTsvkfdstvI8MwkE8zncj50UssG4QML5jVpSoYY9TpM
noDOLwHGx5tfHUW01OD11VIpL6z9x0OebdXeNFUoL2ensCQffmhaCbwqJvvyUd7/qRqC6NouG5E8
iJ52JCBSE32eOaFBda4524ldF6BbCJ0JJlA3d04hiIZvCRU8eLpMU0w5GYZnypq5HH/VjjsGo3tB
K2j9wxUFKPxrgs5Jf0j1EpQd1st8kEZJ19uF1qtkAalImIAz/3N7yND/F1GIpCm+41tXyVBgEkJk
P/1RB30buzyGanG3akw21gXNmZwS7f8N0p5AH6tAom+nxua+RheshbBf3XWBjfw2JUuBtIrs0N+K
Wryl6tT1MtR5y+yfeE3NyVZFiptgCacrG1BbXmhY5zsknGtkqzzKDHK8c0RIRxLxJjvKaZe6gKez
+t7m9r5UVPolVghdBdIPuxQ+o5pL2E75Uem+cJ5c/JXB+W070lbL3pAtoVcERMgL0rmGAvcIFzSx
yhV2DeOwr6HzOegToKTgPUaSveiiPL6mdxhqoZdy8jEFMLZVF8ITVuZL8i5FDF7hEejwGvl7l/BQ
oo14nnCb1RHAh8kQOpYg4Z636YKY85oiIIPqw0dHyEuiu47KNj5seN8iqQkiQyuJNNUIkLnKFD8L
IE1+MyNXUiFUfYX5MXKn5Io98Vu+H42XOQxSy2uwv4RiTqP8NP6vB6m4utFTD09Qiza4h4yCvJPh
0W1670rBqls2ibocdckNl7+4jmCx/n/oLpNomvxOFnPxinwBILuiAyhwz5/cIhKnOPRIRATcIrg/
OVGdkm5qmg38HiU3V1hIuY6xDD2XdMigRY0iGB/9HehpWCMYaq8D7L5tfw9nRI7Ei3JOhFA4ipFz
U+tkvtAEGA3tM4FywkhokipLV2uqVi2w2uqj4LlyBe5ghA37ymrvOciZluNfngMAHhCAhA1Cppkf
QVMfYimhIYAmVFczlLtEXVfV7cOLRxB7kuNPZN4RY0J66wY9JigcGuYRKb4rBAb2FyMzubdN/5vW
owjNfA6AuMMlioCAK3Y4IQO8S/US3LZs6xCwltLrMn9Ax2+XxUGXhgZ/Q05P3qnQ+TeIOmbJAcvD
w+NrfxYKq9sXkbDPhDAcCKUMpFCAUWdI2y9gan81NTviDcNaWjdiB2p5wkVTcLfGxcBkeFROsAa1
HgXiS3sQ3tbUA4A2aAvrIcjHqPO6Qk3T17QCDs/FCLfzwfHEmM5b+ngxqUiCUIndTvHKRQ0ashwI
JIBiwrTTJ9+uLKlfEqEJal4zH9iCMra+EDdDP/tuPn2sj8dRo47oCTvURuA5US11taNgthPl3n6t
exWSYux3LioSQm+u4oIoXJmrKWZ5ubZxU86VTwjbcSVFiD76Y2m2iOjC/6Xze6uZrqMU+nCY05Br
MbZ2MqLsK1Rbbf3N81hotQ/n6osbtA5ahk8WlKRT1M91Vpt+uKPLCmviMdGg+bR9fhdEt2AQ/WCx
TnqRfxYCnSjuBywBerFWXbQ/2M8lYLfFHqBmz1zBMZgU1UfIZcu5o/Pz5wDBnjVfi+m7MxQcXPhk
oLXs9JWDELAYm1Yg1sBjL6lQYi8/YRB95bYI5pwn2xe73sF5ZDkoTyJN4VHrGpWNEa8S+SafDdtB
Mud8fqaxCndAbLf8by9WeUNc+JUzCTE0uqs34B5ekxs2lkrzLnMQC1hXzuJY2iTebrsMUHLSrhcM
Ai7/6umiHO9R0HQZw+TjSpYDQhzdjCzP0VS7DgNV5D3kx7qTkq21+V4J/As3BQYUfXH5eScHSqfd
JXzOCbg4Coh8PtHqIMeU4QDMyLDeGkU0+77qforoovZSWzEAUBZ1RcapdAd4Xc9jFspUYAFAJSKS
IdcrYX1kF05mgfinuPiI1w8aOqpTmtkfqXmwBkyj+w2PTDVAIE3N8maQdEmGD35F9qpAH/YxogIK
ZJ8WhawD0fXKge6rKy4ek5S+qi3fijrVurV6ICpwl2r9/LdbwQjbyxFAjGqBFMKPNSlSRFEceenI
W9uP+piN9hmtreHPYuYZoKuUFcOGMvsHJrfKI82f3YYpxJ4tsLHWuYzFbiHBkPNJHtv1hNfX6d0X
wBJeqEx/n4Lu7qL1MmhEqrI0Hj2jZwfgBOoANUBihAKtknTPZxTyTQQlNyv1ArA2EXZIqdfnU2/3
K3Ve14ONn8HLdZQtW+yzvqHH3/C7SmmIsVlPl5EHmdC6NPQ0vXvJAz5uzHjb7SNQT0En7gccMJW/
4x2OgAVMMEyTms1MxGEDdbghfGvD0NiB1jWam3YZqPYeg4AoRq0Z+m4+gZDUBSkinVL2jI1lfZzA
aXNPvYO1nt8Zctp5qSw5dwky9MUPoKtdu4LRMIlJL5wB+ZIyybEJZ8hm0p7CfKJjPugHSvjv+sf3
lyze6mLWxL54sfz/4vcxz5f+n7+VqBb6XSWIk/O0bjMtawzQ+a4VyH6aaqhdE3QyCEXVZRjLPGa3
OEFAOQ53WVnBFjAen2egjyLue6Z2O5zlpkT1IEGcbsVn91fMM98lZGIqtRwj8vc+ifH1BHQ1ftmm
LRpQ3PorZciHox0jRhCF0SSh6xK33o6JpTQgN9zk6c5yPwRJAzULLS2w+MG4tKNeACEzEv2On6Qu
mpnTm7ZZ9Wg1hdsPpzD10+iooxTSVBRuC6GVdytouA3k14kMv7BWGJ4Zye7c/DIC7faW7LQOd0qK
6M6D14etergE2QfrIbT50yT9VnBD498v4bAg4Zt7+Pp7tNkiakvc0iJIt+uqHbMY+f/jxtAuMCFC
SZwbXdJGimXDsZYd7U+sg1WMsZqKc7RctKCTFL8OfOq+7eFj6Lt4roSVe1xUn6ZCWcqeiCguOAQk
WnqjRiIWKqAUAI9XCVBqtOK6J5RtgTwpyW5aTCdMHOu5Uesob8fSnswKVoUKbjh1NA0/9WKSi+rw
32xvnITDcYb5y7MqqGLMqgEWobS/XGtVzxgE4LJ6hIcLAaSaTnmaPXmOyhXSbVfyUEjhyj4l+r9i
RjuySGWAIbinB8NS1RvJffufFVTJae1j60qUebGkjWVyOzTdK9H8Gg56rC8JeISLKPgOjgu39Kjt
Mx6Ti2BTOHyqhwUjqVcb9Q6Iz/B1q5txU2mf+z8G3A/OtXYs98xbzNVaWGOvX/Kurmn1CdkmolGD
HdYLsQiULtTdFOl5RW+76qjFTBlIuDM6P3fV00ALyAXDPHU/6iOjlkptwiRC5LW8o9s5Me1KR8LB
ePKaUWolLAyfaJv1KGwlaJ0oAh4BEiilKpHj2EngzmxbmzpQPyt7wkLDqHL1Gi1O0sLn4u3kPDV7
8Zfb++D/bzd/XeXFa1mvkXwdRE+pO9m+/S9JjKeViolLdXxfq27Es26JWVv3NOjhP2uf5ukj9L6X
uPwGcGpCNk8+8BmD/Epq3o02xa1D2QQrr0RdKheS8/ItjDLNOvjc3FMG8Ubdzcjliy3ft2uOHTo6
mDwFbjCDV0x8GKdvtHROGoCnFMUcNFtSthwSvlPaNNlfFrY0zw2KRmHSYKtIhX9dndDv3pcqm1CS
6VzzoQtvLk0MIYARa53EHzmjORrXnqASfdc01WCcjACMPp2p3veFSIgRE4Sf77rkL8IeMXLr4bvW
S2fJBooGDYOfkzva3e8kFCg1SNxOoG/IFmXBmVjUIMr/3GSmcrA9qwLuXpByarqb6I+76QZkH6dq
b0EW0lF120eYJ57ooBPKUNy1wAKGI4Asmx7ZGBhuNZdmCQzHRDzmqKLDL/5YLRM/uWtok+5i60xm
dBSTs5QeCofG0wPF3OXEYLFipxraM1NyVVk4AwQiE6144tvjzvT/FQ7GEFHJW8IQyQCIJfNC3KfG
HNrxWrF0pz17q29KoB+3SJSJRxP1zAlaxTEQqbUDQtn39wYxZMZBr2l8FV8edVmH5jIef0u19ifq
JAI8OlZA4gqLd3qj5Xaqjkm5JvblLFqaNO8MdMjB92nhzKfVZvmH3x9MYASbXNB8GatZ67bK358j
wWayxQ6orRVz7BeKTJKIHQJsVLJ2SKvWkJlLa4GZVWsw6Bl2Dr2Y+1QogK2h2lBpt3in7PZQwMry
g6D8Hi4lraVtPCB9pjonQwmmh8bEnOddqWWInjy3owzaUKeYMyLaE50hvpjcoPunrWPBMwsd3CYo
hr5GnH83xPWDM1xnEOTefMdolgRt5iZO7Gvg4qh7Sq0kwvIpig1czSecBEdOdyOeMuDTfcUUcduu
fHTR8Ps9jaeptcqk8+ph323MEnpgezz/nIqXHcgfGQG3xSiB4pk+4da2s/f2c11kPKlrR9GMN0g4
3voyidqK013zrK+A64NI7brKLSaSl1p6SuZ+F8Meyae1uwL+fVn675lvHFQK/0GW/DwE//NTEqLw
9u99kjScUwwLSxZiGK/3PIkT2YjIW3biLLkC9awknQKJztOc9Jll2ZTnFNGnjHDPmvtJacGHmlZg
Rb2+xOVq/JQahgdxBd5ONMZm27SCcOL5Rwdti126ICiizyyxWfhF4ikso8sFrarUfxaKYSkVFSeE
x+VmK+IDv3T+107cr/6HFKlofBHaFOyDXyAfvgqN17frkymNV7+5dtU0BIccZuq6faaJ+2Qf92w2
AiwM0BgsRGkQoB0OvHzsOBJ8TQ6XCP91Tww9JUHEHS1dt41X2m6AUZ0HSWFB4/QhRVMTO5GAKQwW
Kf3s9sLuuYADooEXedeT2NeysvFlkCBWjtbeaWuQoNjDwhXAkO5s9EkA7bBZ50ql+a3Vl3mRR49A
Q0zmYnA08zvGtBb4Fv4ioCY1ljGkwV837eCA7OURmG50LLgrp7grW3BagUMmfbG1C6LhoKoax9vJ
/jKLAIOBke+Y60Hr8RKNUqYDa4tTyCkBydGEyLYGoQVqVYWvKTiHcXk7ngZwFxpn33ypiNg/A95z
CpvkIGYv8rTsJ/9EaPoqen1DH3CJNkSLxjZMBsMEh6F11JZFwceC9L5vsg7VIWWh8wCQNk1FfYxN
337KoYTrFTeW2xaUlbOf1k4/ekeLaoVWtT5ny5h8PwELYa3jY3grqc+5VHSDFHJVtyV+BeFW0QC5
BHFQt+dBRI7hrZzfS7yMXmDZEU4WvajZ2rwFevNzCQT0F7WNSHfjszaGTzQLq0FtQfBBQxpYCLNh
4efktyDzhU2eHX1POYAf+gwiAT63d94sL3d0NSvOYzE7TXrsM5Z58Ae2kAcWWFV2pB4aaqpveLm+
0ucD36YaZhuE1LpywltOzX1kKCzzYcyCnvZglG5sO5U3whHM+kQphqhroxdzEf0Z/oqC5aeKTOHO
Yk+rLRH1DywBUy3AZ7wzoDXHDhaTd6ECmaNzQ+QF+jNfUEJq2/sX9+njHWuYlkRkwXqxRroMblUV
34Cl6SI4Q06qUr+dS+8qZSrznQltR5qb4iDEBPUzmLU/h43QX/jO9+/96UviYFbemXDN0kdGTV4K
p/czaayQjyh5Fz9EHY5TBWz28Pdp/Qwc8BkqPVbtN+uV7m0FVErDS02+CvQRUGdRkSxaEbfdszby
AjVs939Xwk4pvdzEcFkLsN2meF7mlqeULV3geXxKkrzhL08PqDapr9fejn+x/ezBFn5nO5l2tDDa
SuDmv4+cFgeFrkPDVvGaX/ucvI7xulbUVvNl//zIe9orpbtFFHcdP1vzupBqkyLat8JnyGki5OIc
B/cf5zXdEUJn9uqF9CO9fluMKGouKL6JxkXfwbIOUX9GJWRfyphVNbH3IDhb7F8Q4Y5rylmVER2F
EjJvlIcIYIVcuFcMsn/jTnTsQtFyXmOWHieXwmZIi/fh6KW5Ki9dBUqnFYyPJ4o5IQjdXjD9HhP2
8RjCrGdhgXgI88sj2zIqVAFcpHljlOTkekOeNuBddklimFEpevWwMZdffzsignynSreo1sa3DKOq
1aG65ErDA11RclyKoF2rJI3iEe74gl/YmwxjODTndYM45MHWoXVFZJa5MiLwbg1pmlQzwIKXqySn
bZN7u31y7HpAzo5iLetXChbaqX9jLVpr073pC6RrJfhBKbGp4+9CqvnL2DpNw75Op5uUX1lsnTS5
UdcVXocfyvfiORB+SdZ8Vwf5dVbLFu1806UeZKGgZYI7mTx4hsWd1L4BGZ76eUq+sIcw/tPJMNh0
sbFyCFlmBV/a9MiK5PgX6Om3ddLWxTSnM5rILrXYuiEDq/Wvb7D0BdPTxkReJwXUrwK0Sht3ewGb
r2FQSbOnIwPp8Ra8okbZ9Lw6u+obe8CgJJogf9JBtF/Cka2pJtxrBQ0VSA8FZ9kSvfbfJuVI+Ld8
23CJ32vJpRV+u/kdg2eTcWzULTW485HEvIt7K39/8IecLEMaaAtzVN78Wnz/oCJCPjd+l+P3iVAJ
HI45BWcIC0S1Tznir3ED2G4czYCCJ8Tnpul27JWTCF+Us4HfDPBlXSQg4n+4lK8Z1D4xE6vf41y5
Envq8R7vEfXlmuENKpdZk+tDdu2Xsxy3ISQw88TMubSGsKgwgA4mB7rWqn1JA6qy+6xawzwHX1ow
dReGyeibg91fCil0VsDtl2eoC5MLTMWIqYgBlu/B7OExGQckcTCLhtkXu5i9hnjxmTqJ2QR3CNMf
TNRD2Zqjao6jEF78ulDA40aUr7D2p+KHfnkJnuIi+5vIMpvpSMpZdoC+UDai9LEKeQNXhyFNjtPQ
MJzjdFRpceZgWkAW8phsxc8N6QDYBk4cW5K9+aAXROn8N1pRLjh5eU+Wj58oNHn/lZIUh+W9oORP
nIUp/6dz7fHmklc5UwzKt3hyBv2HL9x021CYctrLk87BxdKpfnUTrSNCFO3BQtOsPn5MhIIpm8fd
l7z+IP3zxkc1bm1wnpHmWFp3NHqiUYcn9sArk7m/LYWR0ndNFodl8LSiw2VNvBtfh1ERapWgRvMq
DIE734aIPVcFdz00uWRPF0GsKIK5hiHU5t8YzLZ+MGkxH+vUaZAfC2wvaafwKR6WucwOIU4DFVA2
x+HfDOlOuQskgnkGUWr8CCLuj4PvqFudgzp64CFeomOEqwPr1jT3tvsao4OyDljnkBSNugBiSw38
53P5YGoKBijNHIDYfCDEd2+TCg62zWQLrO061XaNos3YPYVxjLiLuBTqYEPcYSQp4zTQiLt/1ETe
MND4d7B+4twraimxoBlNY+zd2Ld9Euq9OhslxuWux0xGUBN4QC8W4UOJ7vn+pO+baBnQ6kLR8C7n
XJGKFXLit2vNWNMZjyf29Nr7JCPZ9URiEkTrt73nDSVDR1K3UbAMwHugW0h1b9BkZQKv0IxqLnhC
o965dyGrnK8l9U/oshqDB7bEznKl3dlYLLGemf4FlYNSTzXB5hTauEhXJgIrhIKEGVRt4mxblsIU
ZK58js8BV4fruzuKi9Zjt8U689Ho4iy1CcTu5yOOUARtns8hqWVzqMiV4B5S7X7Rnb1+gzS+GgeZ
FVlG8Am+jtO5BsXbhbEE5EfCcUynvhqlHGfnIe5jePfqktsnMGN65dk25fe5KIWuR90Ep2u4OAFs
u0Hlxw9BRPPaFvEnUFjZTwFnJQUp8RzmK9eDJyG2IfGcsZ0PSWTYtOFS2gaY5XFeguPGZ7bETjA4
r6ukAVQUiR99S/P2SfWBaiaQFBz/Y2Of4Qd1/OqUn35CsGRa4NWGX17TZGP7fmVj8jriRyYpsyOF
8sHJYGPBIxYL6jieSKu7lDL4dvg84PyDUrn87FuRiHt//ZcMOE18dWrjtqKOH2rOD9aQ1M2ShfJx
bcLLKNpuiZcbFKcts66k4T9MO1u+zco92lMHy/2c8QjFtaZDPn9WYHk2EmKY6QODSRas0pcbvZ/f
rRFT8cUZIKw8+oO48q85OkG45s0CkZ5PiPvbYA8cwenIIMOiLZjQ6nUjbBJ0IJKhEt9rQxixUV5R
ljxTHMndlJA3q/K8Ie+N4g8g5X4gw/sb9TQi4ImpRyVoUVSmmfGYFMMb1Ff9ClBsjsYUmratIxIE
XMdtt5AxFBG3Zy7RDwywghiOnemXmNh0BVje/aBdtPs3J3ANn7DDU7Zg+lS0zZxBEKWDbBBxk5fl
eCdz8QR/0sdCrjUyu/RAPbXfpuhn+sQXUna9a3kRlIlGJt7nPaufKWfPRtYf17kO18hcVRIWjiXp
Ncnqd837cCxM3RrcJkBz6GeINeeZOO3fSAkiHKWPBcO9WHiAtL08ny63k0Zn9rsFRf3OGvpDZUBD
0/jRMhL+oP/9o0EQdsZuKNySX9XgrEruD9Vmt5Rz+7uALh6Ib81JLZWyns3XXS/jJisBvD8JuHja
h49nV+iLTQ3Vd/0eOOxwZ1Hopru7LHLcF/75m9oU0jC0zg7ii6uuRhotaCas5rCXWI6erp/D+OgX
Jfx0vkYevJfT+8pkOLAA+SzDGytYi7MYt+8jum5o5PwGkc+6nf2KNXOYYCBTHCqHky2Z8dX04t67
xrAbwek+i/WN0j9GxSxhGoAmlFpqio2eBGvOb+vMj+yAoFx6UUfOT5ikLLeemKWGMoQmE+phk+3u
5OUraWeDbJL+dzfACbBEa48LxqMV8VkpkonLcFuOZq2FnJfjePgWxdwqFY8IaH3C9iqgRGhuS03s
ryYBz/Jr0Ao4IE0ABWuhdn+Fbh91b12YIRQnitqqStbrUc+q9DTbicfsMte77d5qfyjYzgTANTUU
Y+i00vi5E8tvZDXgFqmytQbwEfXZEvNRtyINptDfOQj2uB7WQv+GyzEoFJTtcj/s+YyCD9u7c6ZM
Kj30dNgsv4ZiKToCEvm4PB2ZNAiE6Y5GpU5JsDkQVge9KUqiFhTGqwiaQ4Wp1lp/UdVKJeXoW5uo
Oyp/YyLGmCpI2NtbAn1XTgsazT0G9o3ZT7FJIndfXOt59VNJzabub5Cb9wAEZH4Hc7jD1Ak1USFn
WLvUJgLPc9dHa87lwFwGKWzmOWRtitYKmWCXAqNSDUffTlu0BhqfanCb75r+dP8HN/LwkwWEpELl
WsrVETQB0Sld1fyr6uDn/tWJlZ2qfDCOTvFm+DuD+VuZwF6m71FBeA7pZzVFIcYD6zR3yb0YffiJ
k3wwFYl+QePVH9/MdOZsPYkso1w010E9CJh2JZI/bvgoxPjUgrfvYyMR/oJwlSoroyLpHCh5VtZy
14TZ0EvvDTaWkVMz5CvUorKAuQ658JpXQIAfQ/JyHsrW47ZseEWeia51+g3Bsp79Hs3CNHaWws5J
aJxxNaEjcZnqZ8xcqaBptGfGRSF5Ks+LNU9l2njREGxvArjgLvlKz/slvjrF0BGOtOgnT2gPiO2w
xDgoFmnX8Cn5LtBbxJwQYJgbvgYNLiiNS2dQPyw2g+sX5+yeWdPbtZURiI5SdjNz8ielrfPw0CBW
BFk3XArhGYeebWSIFhYIDDjHUxsuzd9yTEe/imwtYlftt5dc8OgK78MXOjkwvh0f0UHkt2POH9p5
C4e8EuX+fST1gu8VCbulam2JI5BwIOV0NjzoSwmS6bn72vHF2glshhtx9m6Odrw064cu2RMtd4dt
MPI6NqoK/CkjwRONEUXKxdlXzBHVaAWZqrPnq7ltNXd1dGlieRnLWmwyE+dcUghYPVKr5dw2jRMz
IGo2HFH3VGdwqq1xpJ5h310hmWW+9mZHszLQjKttNycMCLcA63gXnfGri0m8qa+v0E5quA40aRwh
eBjEkenpXamSpUrhzEBeQBrBA5IRW6L5ehV0ER95onHj6kvr/XwRNm7iaSLZ4+B6cORnNWIJc+fX
XddnxOdkuQzjzAR8U7Lr+MI2QYUR2TZx9Xb1hqChA2b86KxeQiT+g1IOKr7kGq7HHEC/e6ld4tRU
KZe33XUHnbtlOsQDHWSilUNFOWlJ4YvxUdQ7VfY/ajB526RA2gw5zgPtPzwNXNIVntYvWi2Jn8Fx
EJHTe7XFp+SNg+zjE4mlzwwvGlLtMAh9p8ocddnN+KotCJXkmrn+tfjo6zRlPhAOHmGKhVUslmyH
FdAf3CC/BCgeye+a8O823HwZhKzdPGuNEkPMbKbrbIQjc/0HbPwnJ341VqdTmpGw9q2w6ThxSdBB
Pqakxdbdbyty/9sUqI5rWRMyL+baoNl3it5HgX8MzPCEPsqdwj4x2AEdVTTaUWJIKusKQ6sVlpDm
Nog6MMkUxZTtVpw90BzQ4B3VRRAFmi+ZuWKkVw6/cj27CYcJkJS0p3/8CrLk6Ok+06kkOYi1HFwP
6DEbCau6eUyWgor7qVr8uvtazB6NkPj50CGut7eKgwvUdJvjvaTxgXfMKVWGY2oqjYZJTrLxJ0ur
KDjoC/1DtDF8rkumdsTgVzSk3OJ1NznS8db6wCOq1yCKGg+cxeGkbm1dZ6hJhV/7PnA+WtWHh7fT
wTOoaEo/TKyKK5c1FkJJbHij12UG2Bfc/uBfIOz6/C5caG9Yog23vE0jFQJOEnRI+5EuEyGlwEJ1
asUrntjka9O1byYqUmaC58fk4rxLivWNr1Jhp1o1lGlhWxJY3jrYHCn9+4Yc9zgblsll6Bsk1tHf
MXAXuaS1uwrdGsc3EIi+jmO9+JHbs2nKMwwR7CynmgiB8v3cQQ2Md+GDzGr6lyU+shFWAuOjybUL
uWc63XXCAEzAHAyD73ai5YCeielCIzaNJf1vKHCvP7Fz5cV2AZXACo/X4x/96GE/DSMb2FrGj7wi
z8Xl4UoU35Rvqmk9J5vE4EESz7P8wKor8rsmfboLPeo9WXJ0XadnC5m2H4j6ZDLRTr9k3aW3VEUQ
YeKLLrywuf09ZC7TIhaNdWO6iE2gHxj7OYqx4EHl601nGi7obWrjrouN+kgY4B/GVc8sbbXq5rHA
ImiiCnq/CXwJcjToECvv5FpFhPgDl22KfRu6wkPlA3VtUPFefwnWud/Jg09BbbeNyfxgjOgGEAUe
dyc/khxECvvboUFA2x1SpJEjaPl+FBaRYag95vG1Zd/Wgn+2KdLToAlf4lmZnxf0XU9zncM6y7sP
+i/NfUbAezIW4BzbXQMx4olWX8HkhDhXTXJC3bupmtZ5ihJpFObWGJCVsAsi/HS7dgUXXnfr0Ayl
Xk2W8JXsIJOz1DxPMSy7roIGCnD+yD0pq98cUx9o9o+ZKG4axUjbsIDNYpyh78ugNklz6E1uIQpz
m3VEDylJhDYuCcZQh7xUmxK0hNSVUCUHVUKBzkHevgUdIkbUSiT6rwYvDji1Zv64wBG6Kafo/oYH
hZx4hJkmr91VX3nnQoelEU8WsG+UUr+DIRUDkkgDO+rC43TpZj4lJ8IuBiThSKmuWSaNUkA2h8Bj
5sihmn2ZQRtETtKMdrziVNDFpXYAR2bnAsB8U91XZVfkjuawxdAU4ngxpnyjPXULlWRtoDbltNnh
79KVRgaEI7DXHOdzB0OpWH/ghwDoAGltPTxQCul+jVJ7v2HcAV5sZm6EUizxhKqMVKudf3Dp8Mdd
Cez/enRBvYvwrrN1929nvJcJ+LwCGJSK118kenvciP8tThH/beA219AE0nFmuXUeJYQyqhtAwJ6e
ZfHqH0KzUddgZ0fLq5r13pPZJq7PWmnuCPfCSHy2M+4xX1OnsVGK64wy+dv8idvrSqfH301q0Gy0
gbVYNVOAy28JamMw2LQuZ4PQR0QT0LS1efDqFOkFycbcyIro/0MT8t03xAuFBWdTMGuAH7HevcGn
WzHquqCntKMyAmc4S4o/icvrdANH4EqvhYuMHO189gg4685mb4BLixPYW4Lp//j3FMoGpbQ52UuO
4yU59iR/lYBpskNiZMSocCWHc0mKwjrV69QtvVA9ujVngiFrzX48fDDqHS4gYE5tUzsVDdlFDhdv
m1OSNGW29vYn7l09n6sw3XNlyyZ/PWZ3QdZy5060BWX9X9yNGEK9JABexd5lWqA1pQIldiO+S2dg
wxKmPOu3aGYgdkDTSXf5Y1ey8zheH8fEt5g5WL8UNZ9Mxt8CWMXpCXPO234qvsQ4obie2fVRamdQ
9p/SIGsoCzSVnfxN8LLPnArtDVuFb1eqol1USTAfSwjdC1yloTVKXRmAFiUIztON0x4o9ELGHBDe
+5/amO0IdCViK+0wmuAXbzRqW9CCB32dc/O+NFFfolf7GF/ZirhA1B4GWAgiWhpu6o9/qSUlm/W+
t0pNFw0FRyaTBGPV0KKjyeMKWnPV6lU+cMz2RnlSnYnS9h7JKe6cv+Pghdp2zD4x4Bo6FTD2e8Kx
1O1VclBEpYX5rbaTPVH/3IdywruBgaAWxngUMPU0HOjFEp7uJUqRnihSdXv579qKcB7qgnHG7Hvn
sLf3qu2ryJXQc9Snw0oxhwf3T/Ur3vcd7LHHe/gdm0srD0V9/AHO4IvpTgBDiaTXIeoQ0pzUkIlq
KMpkBz6ej2fsXxuH+LuvWmkEKblLLohoUfTB6QTBHKxFL1poZtcM1Pw3rptQenAzfBmB3SOUyUBo
ZxMJeRl257HrDQBx2JnT5HPHmdqxKiaQEf0tsar3VlcLsbWnyciWSeO7ksSLDpZ1Ss2gjiFGu0GJ
MfbLXsOpC78QFUVNe1MckGetCzhv/CNMYPUftTCOuf7nxQOc/mP0EfqbB5cDaQGc/kSYxhjtuFHz
tE9PU6LI0uNgguCswHSBEODhHYrXLBn65E41GZnBw982+NU8A4s+iIDzktE7/7nurPLpvpkb7EUE
KUE37cQJBwd9jfv1bJ5GeTa/Rp2fwNkyRN9sbiFRGq9E+hS/oat8vHdsl2rpaEPefYOaKN4GQ9Hu
ktRWc/dnXcXVfnEp6NrLwN0aUpK+rw32X8F9veuIXqErEvmq4v8P9afenEUM48o3w6lDMyFnl7Ry
tXMi50RdU6T9B5/hJmGDzQrt0mQYlMDgQj+gt6Cq7YUlU408BAXojaY6P9FY5PuFXUsle2ta3EkR
v38F3tcXSnYmusdBhYratv2SPCuH+sKQbyLrWJm9r32z5f4F4WPPNpB52wRtd2OBZdHwKgGGLVjW
nR3MiU7WjaR185C2t7DVO+32hwSEpaR1WUBfdBoEpxi6HkeT2+MmuLcniuq0qGAkc+Jo2owdg4ZA
yiWN7y//GbYrLBW9sCffUGXxVrs2BImOajmWBlLHFgzv03E5aGAp2FSyA5suzsYaRknBnGvPf2gb
0J/fxujX3Ucb4qCmfjJ9PWjjweNd6OWms5zwswLHKTemdIi0w/bcGXYMQ5391Gm+8R77RGlMho1P
lPypW6qXbIX+Q96tJWw/ABhXALE8IxNtqUBtKocPTdUOlc+7mLF/eczr1c6LEGQNgZTtwsEy1qdb
fniSmDw5Kby756OqE2J/xF8rfKtu/gsvd48we9R6LuU/96vAr3Fok+bj6zTIzO6TgVtjfgGMk5be
wbYPEaKOiEMPKbRefvDm3IX6JkzhWIAAA1yqGYAnCwJKo5LkSMIPre4J2aGqOIxibqi3VNbx80XV
Op9oys5MIYaQrsuUKitdOTHUItEVNTraol/YRPdKpR1ZSq0ZoyhDl403EaUyMxsgYAvohIluPxGy
W+KcVxuOK41qPwqz3wVFIgOA0Zwyhx2nnawjha9GnP0BWG4OFyMhuJYsWynwDedDDZBMy6jHjVy/
1ZBeYbFW5C37QEyoiLJuHvEczokWfZ+MnoK29AgURCTTEGeFWyJh8HMfw2li1Ffb9wpEeM85NsU8
l0dPFXXL199N8biiT1K6qnN5N83nDua56hAADuqY7L+skXo1WOhQrtzUISwwhg7LbUjeLa04sdhk
6DE77z+1sz0fFF2UcENDL/DvHAmKxaewFu7XckRgT0NDmjEVd0dLL2JZHDll52nT5lFLaFOItrl6
BW/FsuqwgQxtKmyekkqo3mVCeKq9lD+CgG+Wpnb+vlC15XcB4kfcLgPlHHfzlyf3ie3wtx/zn4s1
/RGw4QYb1wIwbudM7pSVVdMsrc0ERgiBWT4Q734yHCwLfXojlOW5RaouoXYhbUzbmOulGKG72NRv
uNowu4X9IJ4J/c+AzLgydDVJgHl9R4NljNDPpBHz24jQP0FtnEKgUivl814UjuQ5rYuQR5GdqCGs
tmB1i8CgdD/zzPFt0NQ4kiX1jjBpBOpHsFXSZiW/Tk8jRHhd//sWCBqKTcCfUgvtmvtjyAxOvWhZ
8VEbWpBtsPNgfBGCPAa2kYq6+dffIP1bAUY/kLkFP8Cit499OehHmjJtXjssB7nz/LV4CQPeyqKG
4pZtVE6+mc15Rrwtkbb2iYoyQVpo5PEMnJlzcI0hmo32NI+af4XM3H5jgvnhk1Fiw5wFmU2C5SPD
VK9kLW7l8blAPKbgPp2Dwnpu6fnWyqVmxW/+vOibKRNMnlQ0tnAADvMCSBURscte5PkWAwnxA8k3
tFNOdeXyjNX3gGMderswhjj9+mg373KwR9RwMrZb3NXzrPNhCkkUiTuRHONuRl2v99IyegMAWy+p
VF8H3/KNBBTQzvQJANwaC9VNWr604JLO2usHIkLAhVuY/xLmQ3sMi6RzuibmsWu7wJ01uxWl8yuA
o9g3OB3nhbHc4LFc98pdaMC6pkcJGtt48BITAFRBbr1l/kM/lEWG+rKXz6AVFkAaYGdM5VX5oWYY
TJZAQ+i5fpYh2PZLUe7qmRfzawJ/tJoKu1vV3ivQaIS16O0QqPyIGafMrt84YdGhEoIaBHWhmooB
B6g7rJEucx5kCz2YcgYWl+n9u5wX19QHQFptfR7RzHxM9UR5eqnY7zc6QSWfAFI6pk+gQ+FFKRB+
gR2FsrcYc5tJ8mpEyX0Wz3Nden+yw4QIMnCOgavYqMHfl3nm6c1mDZIo8vKHCsxMLoC34D+jysD5
xO0kMcDwC4rdylmzsI5Y0LYMibIg/qrNVQeNILVQlkjcbB6GL5INy35abM9Y4nEDOJvc23ixAaT4
MTyap6g6boFdtlg1jJwQM8viGJCHHPRBknbWkkNs12Dz2KR6RWtJze/Pm34bPQ1Rw+RyVDSu1C/T
slgYmfH50tzAGnwJ1cr/w/P29z1KuCeFaKK1kEvStHhQ2DyuMzDZS8ak+r0ebWicXV7zxwnSqwRs
W8Ls4D7zWypZI96yuLfXU6ohVsWzcLGkcQiMtJP09qaF4nRD5uFMfaQWG/JMO9K3ig4RJ2uI4wST
3X4axmGvfRcOljlqGsluZ0aqNk+nNZ43AbG3DkdUR1imyTdrpfGzddJlrSrpe4UnQ9zxQY9xTteS
pFxhP9EuEhLLGp6LZzBzqty9waedyYiEN16uxexijC8d8VavK4SGJRxhb52aCNLa3RtslZTyXo6L
h2y0eqaPsc27guCoMaf7OUz/B8gkG+RBzXMMmVoFhsf3OnoEoH+Z6q+mlTltyFfGOu4nPydm9XVp
CLdauzPBbIogLv63qcO3teBvZOPmrOWHgsAnc10UVDCpoutI3bNJ82e5tln9BeOi/GiwZCMg40Zk
bqI+Eze3wWMbeATzHYEQm1lux/Z/15YXwGuRT6ENJ2dYeXFGeDEarPhLmT2VeV3OVwaozUXwULB2
KRp8LLNt5QRh5L9k5dw1/xUVF0a76DQenTbqdI7ZYFEtBW1V5rKZO86TbHDfJT0w/eWm4HyWnbvA
tL+CQ7unO57zOVKkEDiTdeTojN2Y4d3wut+iv7WrhDCrNC+bKUPwc/ZIfyqEgi/qyL8HSYPyxtnm
jCq+Iu8j4QCH7NIZgJDrmyof81x7NmDPSILN9leIgTHD26a7qtuqhyWtXAs98r2DvAfqULwVAsz9
npaajEXnMlhXRGYkleEYJp7cdHo4khKtT6Z8T9d7mNkMBY/Alghe5J4iKhGimsqHm/PzuOpW7zyb
tLwsqKy+jP7QYmPQr4wqn0zr8ngIr8H1NmS/5zqQno66BOsloPo2aFfcP1ZTVg/kPSpTLUk3KCCm
iCH1jaUmeUX3lGn3Cp/0k95wnUWBKHELBxOrfUyA9YqljwmO+8Zi9LZBo6wCIsX27Ry4enpQRJaX
MKXvYeCLrpO1bYJgso7nRcWzJE9erVxael9lb1SCfxejusLVnJi91MeBuCL4eIkKLJfN4o5Gz9iH
ZWLKwOA/HkmBLClcIZaLnJUZG8fwOGfhBwvRV38gz8O3+Ew56VupQ2GCy2q0B8MdhFq041IgTR9T
gSPWVgj4FTQjstE70b84By8NR6uIOJvq6s1QLe3BWdcZjhmOG1XvyMSiz4DK6ACCKrK+8O+UIgl/
BIgEPJmvyPc7RHKtv0yXuQgujfKMYqDGXJRkbCeFnsBztZRRViObzHCO/SBD+2RJalIO0t/ylI9F
bfIGkTl5QPQtGE8ZeWdM0jzR5uPdeuFNFObg+I0iyyUmk+DLKE303X5V22U3HqApjh625w3nrWbA
Phw3Dwnnkkap1y0YvbliPLGlR/glg5vYXks3Dt5vclaw/msGHpiCFMWmpJvBMrbCrRY0A262vm1a
rVTTyMczsIEtU6flVOAmiQluWoa2Fgesoh2CFMsipZogKa5W3Nwa0HUv8VWwIgU6LwKCrNL1t+l1
qA7pj6cNq/ydqzyKCteZg0gJSjL3UqHUyCmw1aETGLrXK/7c4REIqalLI0+RFEc3ghJjBTeOF8EF
ttO03xlXuSqnXMuX/2dlmIFadc+Ya0wSb4qQe8wTz2AoNSl10VzJxPWGoytNpDt72AoyEJCIGWBG
8rVYZ4+uyHHN+p3bdYnGCc6hSoNgFEMMszb4qbytMGhqDLd0YNk4pvIJNikP+S9H3zH0DlJRrdLp
IHaVu/5PHR3VU91Xt4CVlMEErMtAEHavdOPesO1mM57nSEWgqj3INyTQprIw28rVuhdZLTAlsuQw
hnq+8LEEEQLPtmxE12SWWKW7u1nB3PjkLvhGZ+anCUqRkcuZlTm3BXCNISINHqcZ4Ff3xQ0Gd1y0
naoa7f/SYqya3pWtIq34L/e06Ka9kgo0q0DWDaRIPsedTNO8/26RAG4phKiTdEW4iBb5U/HRCZdX
PNy5WujgPwSap5cUAPQbkaafLMBctHrhP/0XyXD77lbPO2sUhMWONwlE076/bqH8BdVr6pGewYKl
Lie9j4UaBtnWfgAhktj5ffVhqEV3WB37bySt/4WAbABoEsmG0WetkH5uS5LKfqaFLShl5Q6/qNvY
51NCVE4a+PQI8qANNulE51w4GW/1RM7b/8DbqsTGjCc82/WZAt8CjHivNLeaUH0ahdJ4d+3Mg6CR
4ED7qPiu2w3faRcys/SmvJNRXksthRAfLNdbHH1SXai1D+Mq981oUgA0zIwd1ymIXAhVgjn60F37
eC8eVjfIwnZ8jVWAykA3TtjAoWBT8lyAJ9XnLCLJuRL4rCyLJV9rrqytTok0m+Ei/F6sRL/e+mYr
1QX6Z6RwIw25YIzGgcrqcFq8l8ltAqquvsD6tjmXE93x9OpOii3y5V7UnB53F10WUjN7eM5d1pxN
vDpNUSLL8K+l25ahAaPoKWEJXdrY2EuBHPZjFWqwPa/PvkXCYIIcgJfjasp29LpzZS15nlYZeJp0
V0MxK5yp5/IhnoNMpOX7rp4mDI7jw2O+nZpTH5NjuxrbKPN/Is8KFdIempWT4tvKbid7hs0lJr6c
TTJYudd2EHShnkx1THw8ffcfQkOf7c5Lr0g0v35L1GIFWXHNHsugS0MbXZbaSkup2HpnkDATfxqE
DRNmRiZPu+vl7AxLUM0Ikr5JmeclqSkFPHhce7Qe4noQO3yWJ1GBoEBo8tE8HrT6t6wyysbUWk6m
XxPuhSPmLVEC5BG4bH2yWpaNj40n0rlvW8GBzv/DOBv7qN4KXpINICUNLIJ4sVAVvDaSE/tvxRw9
F7cLufP6Zcz0Yxye5rXsZNhzgJaFZw8cz5Qq/Sxt/s++VKgoXz/G4HU/v5iurWJ62+QVPlkydSiF
GQUAkAaRjxxDU+zwsLmnljghGlTDb3kYc5RvWA9NPOeQy7AVzkpRrFUCFQywtmeDEy7+zAl05lr2
CruI4LYKViyg0S222y/Wt1X66pyu9+ZzSPwo5QNFrT6QjGRSYISLtTAnBfR0zwYcjPgKqQQytuty
q6usrAmKrVElnpA0kq2QgZ/PM+p+8m3hyqQjW/VLE/I1n+DWGjih4DYvDU6VvZdmx9PrF9Y6cYgq
rf1bNISRUGMCqdXOJ2E4NftV+7M5g8S41lzFoLPuICVyc0BJm+pP7gNuyeGee/6SGcDdpWFe79zO
CllJMaGCsEu7Fv2r7Da3Wa3X5+O9PatoFWkWUOOCLQp2zkC9hw8ZA64vMAvAC7VMNO3L+jM9FE7s
eRH6HpTfjHbjvEKzfk2/Nx4y99q6hHEi7Rfzy22qKJgyJ60u4lZiQ4i15vbUj3EWwDLayFcmSJAR
ejt2NXgLG4s/ZOfXeIL4okhZjG3rRAl6Y/P/h4wS4KFGFdCnQZyxn3r+LunDb7+qjVbKDBRKxzOc
kuuvohnwFmyZ/m9Z6dAF5unE7mr65Mu3nIubpkQriCRw5Dxy7bBS+YH8lFv2A+TeNrEHtPDyi2t8
Y11JJRart04drRiR1yKUQxYJ3bHQIRBU74rdd5wiLIwiLteQphgf4ZWpSeAz6ZFBmnZt8SggeAP6
98S268T95Tlurhk3LUsxl+Ivx1WEZboNXDH1a7Bhl5j7Fu25RcZ+te/6SWg6SFtawZY7CBpyTWfC
9emy0qGFinmd4LkPMF0Unw70HkOxIRdVYsrWe4jgryXwF8XsvRgRkZ1bkXIwrv/ajWGZRdWKksj9
etq0Fgg8ED8MvcMq/dRcbrDvXk9meoPUOyRbcDcr6Nrs0NGAmIbPQAeVB1LeFj+T3/mQje7nSZ1E
LJRASnH519w+5wHmAD/Dxbldlzc910SMZIO+KjCJXaRlmItQOSdddJLf2RVHdWlAoUt5rFTwG0Zt
AFjYZApQNaBGWpnbU3yPamYxGLXRFzZyidnXOypzjUZ6ove+vJ7xin1sfP0FEbajoBkEuHodLcjo
3WsZHQzY9gM6B+/+STe1Hy6Ne7NeFcwIcY8+foPZDf0s0sne7eWKxmL117AT1yEWjvpN02/tq8Rt
HbwkEESageNBAlaEcvv18gKfw3WfRIFM/6DXrZIC3ns8zAXltwd9ZW5HYFvPGFUzlpAHjTNB1T9X
8+KzVRl/DQZy4jF4rdqPcQoy5/NWe7PyZ8H/Wdy2/FJEXlazMYGEOTXPtrqYl8JGxy1UN2BTljRC
8cLB/M/gh87HICvA5F2e20ZY7tR4lX+8CwJVxjuVTgCKjGsAD6mk3Q8XKeGhZnkPPrFShWBtdB5w
lEep4SsEzp7taJfDisFo8q37QnGpI2GpvOTSWwP1cZ5eRY/NO61zazZ1WvUm4ha42xzyWhVp++io
Sx3/Dw3cYe1C0xBMXrXAHAdLXMALGBKxXndJs/UWKAniGpzbLzdGW6Y1tOGLL5a30zYIlOIaG8Le
BtP3wiW90vd+qjkzwwxeWq33ULZibP7+wsPQhgLCXRLkUpoQeHhBhC/OA1HpsOmoh+c/vlJPGKQA
obQSfGwJnobicYGewqrVh0rWKqS1ZoTnid0sUW/Ipq+WFyM8d1J+7kxttLL2/ACfEi49MUdf4+T8
zuvdf5C7AIeSVNwygfI2L0NFAm0gE+/1BUn+db17aRMo70Wv0yC/ajFh+O+KU36MgiN/8uGvH1xj
XQm3iULMS1p0RX8Jm9dT+VdY7qQXyuc7XzyLzKWAEmwf1P3DVN7ukfOC62Z8jF6odVWVbbkYvc7O
MgVidzNtNhCT+uQDiQwrQu7K3TdSOn6SP2LwPYLFCF/c+V1gvqizlWMoCLgssrhQpV56rwsbkk0O
YYso2o7G9HnjV4lNh9oEJYuo7IrRUbVXuNu6bV+uCWmECRfaRihDxHKxSCge9ro5AQZIxov2sJW+
782slmnDqPSC4nfO2tT0gzMj6r5XO6GyW94zNBepjJ7yIhx8/Rsa+Bw2vjeSg8oEXk0G21BcQe5t
vlJF898EucP7Xq+TT3C2veTnwXRVUAMX3vc+wXXeiHnvWOMikOD0o0F56AYZq40y0Zsrof3grmc8
z89d0bpSGi2Po8/SeTligQfIKx0anRYYie/lXl4wR+ZZMticYvpJp7A3LQbkNxRWVzCu6mvqOq0j
dTpIBdC7+vfuHodbXWk7GNqIkfav0iijlLazN/b8omgH6vfUMjT1xmLyh0CspZ9mn8DfDfBJ9bLY
SvhJgItKO9GjR2RPPzdetXJjENBt6RnYGquBk6BzQVr7kMXEe/jAfkFxaoIzi2X7kC+UwqCv0b4q
K6UqWc73hGTcwBoUBd1eYjC0sbCwyz9eds3kVhjxrj6VBUJY6Iq8dxh9fqJcwO4r8LIN76Zs7EL5
K8d0+gT5ykYya3Xz9dKyU1s+z5H0DhKD2s8aZ+XT3NyV/RP+vOuhjxjnCAbCzmCqXhD/agcnxPM3
hrVx9XQuB+IH8eD7zNl53V5usCR5ExL4ShfwlThsvhtYEZGAIZ343erFIKjdWltS6bY7RKm4tChR
cTCaa0CsmNzuV0z+p+juTdD4+pbjYJ45Y6yJfvCw2cRi2HT4WNzntyz3JRhltzPjhxghccOoB2EM
25HSCBhRrY5JrYBMLnBw4aWopJUwuGE6LjHIz/kyVvnddbUFiIB729WWYFcwaNnU9lUiXcHmuNxb
jgLzL0NSLztpzD7eo4bkSO2wfElgDiZKqU6RCkD+HXrBaF+JbU1GOJLpVPMcHoXSw4p/xY3tuFV3
xcj6yHTjqS6YTMNvQMp7PgPZbBb2x3NUNyZF3yHcCEWCUJMfSEZFpAOi5p9cMQxzUjUR5xD7dm7e
p48JQMe/nGmMFZFSa0IF56FGgwbn7iaUqa9VLHvxDuxYDzmphG8puoXffHc66vZ47IZkI3hYw1Ex
Q6UbtzeEymrAyaVBTRXAIGtKUJxXVN3HUpcT/wT+0OFa++ogMQvQJX+EOwQGpjrHVGiWJ9aWBiBr
YG9KJTTGb4hBtXPU2VOSJicZPlehL2y3Khjr5Fb9u2dwPrhuA7GFzrCnWN06AAVdyf1lA8BlnQoi
2aaQ4iEa6e+FqQyJC7fvb0jGGzsgi/TQyZA26C3QKAK+A/OwNpFksCsCwDAJwk5Tn5CThkaOnVku
L8naB375eo9hoSTJEg4LujE05OWFjAMLuW+/cq3Pw/0mVSGSU8LuMHYyROBZlWCCNTira6+uOBrj
24vcWoGhckqZVpVQQwiofFMaiLv7XPDM84XOLOTJ68Lfe654HNb3KjRNEiMZQr6QvBTkk6Oicm1u
mPDZFmI8MrSfRXywD+qrd349pD4C9VynDtRGWRNShN9qIuovPBk5qwVh51s1yfTEwqp2cAeN29as
bm2TaT0870Y4M1pmACN85ZrTzGR/EzJ5JR6IM1WU2bhqpPdfknOHWa3LbadC6LFlGOpBvY/qaUiy
87MDLW7f3fm6Dz662skc9BSvHNSG54o/vYxU6c+NA3G6+zg7byc6vdmmR0Aii+2ODte613etOrFS
nU+brRdfRop1QP+S9WGENJW8LuFL8xQbBwxx7TCDVpCeRQDjpw8jj/UJqt3bCvv4oEpjL4vno9ux
K1L4HNnCK6yiO+kWVQIZSHSQTaNb9cFywAIi71m9nei++8/qJ1zSbJaKADROMgkauQ2nwllrLwW0
H+RL6Rc/Fn+y/OsL7AgAqKs4eK0kX+eJzuaRiRjlJf08nlc5dTyWSo6QWgKvCvDQEF2AqhAoSkaH
EvlkM/1TgER9FUgyE4vnlTivDOgw5/KQZwbE5sxb1Agibae+xHqrzy5JXyQHvPu5oLXnomOY8zf+
QCTyOJXeeRCkffGE6n1pBje4fB8ybexXEWZkdh0NzRZ5+V6yNoVAzeJFFzbh7bAq6piFGkOrLK9b
40hzds11DCoQR3wfaah9WGiumSPBXD6OHxVP8oqpvQ7U0s9Y9TZgxfMzyWS5dWrDoQ+toAPkM0pV
w4K8IwKCbHoAYUAJGCvcqA2nc5scwnn+5ppR/uWP+Yyalt8XMW9Q0l1c6m5MdRcNSbwHpMDaPgG6
Tjt2GZvUiaM4sxHEieCESouNay0ozzvb5djL8FKQ80Ok2I7O/cgmi4a+Wz1CNvvV2aYBACGcJIHF
Uq8qnmH9QmtehgQSNtUB14gUN3EfTlri0+f0u3Y6IOWeWwFwHHkdIdHLAECDyAgAQvIW40CEGaSK
tpHur6VYwGRD2hCwMfY2+qaDzTkaRqSYD9/nCOhjoxU8X/27oAA6PhEaw069e50Boodu6o4D2UhG
lIJRebmtZFoq0IVd1aeBr8n+A+muUFT0Lm0WRkYiRMXt1AeJKxY2bzeBrkaGOHEpXmC7ZHSOTx3N
yic1QxzZjY9rr+AwClDUyaZEZTfXAdsDhEUv1Fxl31sWENb0/u3m9Cg8mP/8MO0sVO94tDSOQJoL
x3Yq68pQzblvcl1CmI1SCZLhTlaf/v+vkEOWL7OLBF3aG6yOUEKaIL31pU4lxAM0xxlUJs2e2fYa
t5SFxUKrU7CyYrvssFIUexfW4ratXyYIH8QoqFLqYZnQgJ91rESz7r7EJiJwZBDTBAGjojYySpB+
0dXCuzdB+lz1MYp4VJdUs6PrT7i0auJKAcDv4oJfWZHfoA8X3fTzZzQi56NtKxWOZtfYzvZUvEM3
l9BxheyDmuglI86OLK6jHC28RgkM3H0WjxtrdcLiJycYqjwFxV6kxTaJBNWqlvNIr02y17m9tTjK
km5xBL1a4tsJU3LLI3LB/4nFVyv8q0vxncVrAzT9ncj8Sz5BZQ6i9Lma19n5iGT2xRG8gzzQQSCw
rcPwLL6hW4HF3uPLuR14Zv/HspRe8wgyd2oMJW2clRwIN4oQQYYff+ll78DTvms/R4vykR1C/sUS
PMJ519cbLp0qapvVPYG6MfI7WEmwsgctyCKWa/mwrr1fsFArNzbTb0SBFLAVfNmzWIYlyTM3Y6J4
GCI9V8a6RYUtGx4h+aimymfSn8TxUVMPSH56jI5BxOu+59xh4q19FOUj17iZiE4vzQtUGHkOlktJ
M2A+ROTGRJntG67rQjaCp8RQp+fPqX8fvtpIHNzyTgEJlzTnG4kVawAspTgB4xXiMDI1rL+ct3OI
DibfI0HVAsMwc0JpLMtLaXETlEN5stF6JRUHAYdhJIoxyUWx1iw/aDWdTuG1G0y5a4VSh2/J4yGQ
qU+RxLoZ/NCHTb/SF385o+pxWtQft41ZRx040NeWUov531wcOEw0uyIrCeMhHM+j4HAYwSZ8pH6d
4AhsyA7CXx02k1l5XKBTkurbYyIbCRU5m2BYoYcE3cG1fOzGJjmfB90FdTSMMuht55kTrmn0cUuA
i5PrzUKcnAdBi51xdA9oi2Vh0UGYjMiXynfuBMYelxNoFl10K2RJEotHj+YIUn+uiTLClS8QWChT
jbpGOIrdgVgGh2p6VVUfn4gt+rMyQLXy2uEqVEJQvVFc7V37a2+fE6QKdNPWfTcJ5k0bjHyCCqS1
Ti9DWFdJwudGvJkoxeHzN8R3TmCXHOn1tnNIrKTzOAOpJkYT48EoaS8CByHVcs8Cl0wpZqTX5Wcn
nHH8fEs69ON8mPjLPRzGZIhuLjHlXFmjqmCPj9Hrahm4knBsktbwd9wF4BvS36N594po0SHjKRup
jekXiRFyn+XN+FzOsR6iec2asDpWm3op7EAAnXgNMGN2LMLljMhQCjyVcG7WcZbakdyzh6oBtlQw
yWWFVqqHmeBqvFaIWzjcGvt/QpqBtEEpvaoiYwa08M7beGEkNXKKZyxBTjrb7jTrauE4ki8ujudY
ACzr0mN4Ws/1Jnw4altisgPXfqFjt3vi6xDtIE7zkloClz1Cxi06cqUw0xRwAZ4atETrhs8vGPzP
pVMO7i9aXCwNqaWicvByvnJJ5fKXRMd0tQjrwYlKp5ejs0IPCRKa1ABIL/wxFzbWIibN5Zoryi0U
Hl/xQpen5Lmd0Xln/g6sLYCmkmabQZIpyLOIJVs6jBJv2u5VoJHVkd1+qQrBCZCnoXC0m4LW0YFy
sbrBULUte4sNGr8+tuk07+4Lt7XBlu/YdODhGVvpGv4Kwzruvw3Cn2Ur4geYbMoOlidbJJ0jWNP3
upbb+M0qQFpj+Z5WCbDUYoLmATj91Neik+RRXQ99+ZcvtlYu8LLA9crpd7O5f6E3wfr4qoKIINol
oxHdk4AzxISAnnUNsvPPVcld2RzVaZEme9zlZrnN80T+Uz/fhkWBOOUzXuBEELM53WOHvGs6meT+
tN9vds8dm7jMztODRTBild008NMOj8PGtdtm1JwLDNKUqm9kE+UVIKFbOUve6vQm4t3Pv+YQvnPh
WW9ZgvaIlTVN3n8wz9Jhp2KcyNq8LVO+Z2aqZzPQ29kukY9lXzSwJFEVt4XDdRcOx/PhofBrizyK
e3eWNbnZhWmbWqkj51SGm4tPXyE/UT/ljvP2JkqFcCdVcylC28l03z6rGqH3JFVSDcQyflcpIU5f
nkMVrMkzmZMGUrdQo+gHKebuTjozxa4Mbdeyhh9XYRyjNPEBChDmMd1JcoFiRNmPMiS3SL8suLXU
Jz01APyKSI3N/05AgUIMLkJetmHJH7gVO4lq1z1xg3f6brK8wGdQp2dCz00mNafaXv+IDqmmq+wT
EphKIJT89AHYYMAQBLFRend/g6cqwZZ0rOQDwu6pGLmANVq9ktgk0v+eb57hgUFZdKivNQ/G4fEV
iCxXcEwOBXD4qvAwGOTK/UJfgPAt62rtcSyRTYWhApDsMHpH5bhIjOkX/i0Jt4MnD6f5MLnjGNBg
e6xdyghE75jsRTA1F76d0QXmfOvlBIgnW79rk2VvNi2EEToVa2T5KH+2Df1+FAvvET5SgC3jr7Zr
WYmPsoMd+SS7TLQ28XdYMyVWipC4vBbMeXpSH3cvJHaHBdJ8Ah7wNmdcgPUSuUm6/c1manlvYC5+
OA93+n107w9GmHMdaf1pCqtMjgPvJVa8TJibCjsTucjY5nyawcKasM9IA5Uffn41EIWYp1zotJSS
XxkeYb1qjXDjqp+Xfds/hrnlZB8ydxZjGUOfeOi+QgM76PuCvaog/YD67ze9tIIvDSIjYqwozSFx
3VQBPnLIOtQ33AnZJXT/PSK41eh8ohaUirdUmgx1E1O0hCeHiYGyUyH9O1ThAaHm9W8zVclmhWf0
BCB9/4dJisFpdpmyHdQhikCusZ4B0fl9wMy+af5Ku2mETuErjrzOP3GY/CbROjqKfIfWl5ELSM2V
jEO0tf1eK7KCugrD+RMzkOWT/UnQqEdfGy5dinXbE6KWOIJUzs8khN83m9eDs4hziWBM5WeZyvT3
c8a6Ng+3cCM6Xo4aEh1uwsV/N0Z1zbNnEbsGYD1vBWo1QYCTUXnyVZYBobHUujmGNbZ6GVs9ZLkw
w6pSL207Ly/+X5CyDQLynfzEczD/AIJQ4+cWdxvLa+YxR+PaOku3blnjn4YddWjLexqpvMWLx6h1
H2yKtBxfR0QF9iotpw9nEMICZx633jvSqyY9fAvtPyYppA0VfHFC1ys17P4XSDrGNkAgBJ1R+jhk
J9ab0bqOsJ4FFX0gmuZWufWwA1nmkNHyG+JvLV8q9WDqOLs/IaaB6+2cdQj/rH7oOgJpIdxqGUGg
rGLuFbHI6GVPxpPxWBhDczc/m0NFYrpRlfyiLTu7YqvOS0bb8zFdfzHemDUTc/C2WSErc7s416Tm
Lkav44PgmIzz1oy3S5YGcHYLkD3azSC7AQQvHHXCoQSnWQpE/C/OmJLOwMXk57ukhbKbY5XNS+lM
/W9P4Mm4ZqP+DEccv0ODuq5k5DxODP1HhmMNyWJJmulH0AMKxRiT05WIq8wUoW44GerKZsArGQ78
LGcQkqXukmIwjr4iEdFYXy8DIttikohKX8oN7rSt13vO1BGIvl3pwg54gLbMtpm6B0T/ivx6eC4p
Kk1xf6vBPPbhYRlLicnKU4nyBSRyWur1g1MWOyzzLcl6UEkiG7aviPN01yx8ORX5hZEoQllATJoA
ayDHpDskJSbo70GEfaKxVlBAvP5r+zieYMOWHZE3GVgNIdJR78TD+qLo8P/8a1TafUw8tC/lfW0s
Wa+G3TT8LtftTuVtTdidK1TeIMV+LTgY8Cp7x8nRpU7P5uriL9zmv9IHRrBfpkT7Fpi63foY8JA3
LWh7bC23+/s9JRDwNrOuDjNPDM8vk/+LphsFAchnSVrjOmA196EeLS4cdmCbMuKgYX9khqE/sZov
vOqO5vg+lQEfIJ6NA1UXrLG8xAwoTZr/Rpt1eV5S/55m5cqYHphFN9ruS1qZQxGQwdksGz/H3f+0
LS0hoOgbjtwkOvgkCnRbGsr+i40FnI7vQdV3XzfAjxBtBbujqGInhho4yFQqdRuqAhu1HcHKaoMV
Do5RX2qKlsLGT6qHxty6j9W9Ecvd/F+PYNvnoFq5vERwn++Yfjwpl3FaFE2RlVWat2NiyvIlAyAH
KucDRnIuXX7D4xMUYXDnU4NvYKsVdKyEXYwYbuwFjCIjpCmvgRmDYX/9z+pIRmfLYrfrnjOUPoo5
2w2sIM6mxJLBXk+am2hGYd87K0+djkfiffyUYFTymnGyTJaxaRv9uE2cGYEBOhmbw1jS2pt5vh9N
zcDnyMOuIxW3a7e+hSQ0eC3G4A7Yy8/8Ih9Xs4Wt7S49GmOCqZeXtlE9zA3nTy53RVFFOEcpA0/q
BQiNmoPxJMaolfp0HDoonGbh4LJ1MhGLieWlvNmYfPZNhRo60UosEEP7xMdaTbdRgQQkDKS+q2MB
lq9E+dUWLp6KcD2vrajBU3DC5vy1UHIApMUnGJ7eNe0KVkYFEr4DIxXzPvm/Y3m1zfNvjSGNqEfr
/leUbnhKJPLabmiVg/bqHdzT3r04pLobjrzan0/8Z3197Tf8M+5s3Lw5bxzOFbaNXtTKL/svS6hE
IXvT+ed9c1Juxgmko8ewToJLohG82+U4Bqn7gazILhqnqcB1Jfw4sXgc5v/Nlw3QTrdhRKeL56fp
cJbMsni+DIbxTt917ax+9XjMC1wJesr6/pzSUZ5DTvKK5TEDUmu5B3WmFDsG2OqeKjeuXUyxRCnr
vxyOEhj8PUbz1l54ZBdbaHOJpT+I2nzVVEuKYYYOPszCmNusYjLQGrDTIaWsFEL++qJ/9T0af0Rh
Vgc8cKpm2p7FMSYgclJogIMiCj5AL/rSujFwyfw54bymRDB0WYPYNmOqAjv0/wNL8hf3w66NRLJw
b73ni1INZV+lFBJCoTZ7a2W588dA04m3S2ZqrnEyR2hEMwqVSB3FjTrGHu5HBWzJjgD/UwEFceYn
RooLNrfSse6FAO1POAVTc7RYZ1Qi03SvLJgKN2yeMlJPyYOVmaZ3ragmmOtC2yQTUsU5OwIzvE6X
PXvuMM7Sk4x+RESZcfC8jt0+2MoIDifNpf3K5HXJ2okNdtRgi5wrY3O5Qsok8KPXme66xKAA9PTs
UwyFnY96Ufcs+lxjIlRn09yzR2APrpSAS0SKrgXKZ7lAu0Mj5iYyUYH/PFpkJb+CgkFRDudXUBvH
Q+SPyRsVhu0PM5i+KaRM+8q8CUIclMTwvZELJ+nFWDUASrcYFHOj7ScmQXJfMVOugBt4LZqbZDPe
cmegop2HRDqgfgKsFlaqKp6Kf46rQIgV2LoJEw004pMDXIKxWVP/yovPSF4ceBhGyscpm2Uwu1el
Alj2+dsFLxvWfsSjB72oFzuo9kb+qzT1OwYWgoKfvoB6BZ9Wr2oDvJD/VNY9hkfIEfIif05Tpgzz
468jOtK5qyoBrNOlVwykeYxWXw0fiwH2W+9SNFkRQ7b7IubTpQ/daa6UiOgLRH34cGhV6v9CZ5SU
4PTeHIhtkLHNaWDqizeHDx/ALmDmAC1ni1D7e+oRHM2HsEZxz6Vgw2W+vp8L3Zta59dk0K4JuX8M
xpsCBDUrZFC7ffV/9kCwMxWuGWhmEM8lVvrYWD1BNxq2uo6U19OZ5Gkswg+HPmLsLyDok9WO3T9t
AwFvQiDjUUa4sOP2gbBEIWGW3PpjA+rLMM/4nIkXHiz/jUIGvqUxRg+S32H2PWjV7fekQbytFtfz
Vc905B4Tlwzvr84+fOSfVf1+assAumDOK0arXyY63kJPj4pfyBZ8NhzIorGLTEZAtjVndNiCUsGp
VvyWdKKcKB6geT4MH9qp+DXNcKslg8VzlyefpVnjsaeqMtghkdaAs6cf4B+gOZ4LNKCVruotS583
0eVIbhJzyJFIpKYdZerDXxwplt/I93Cfj+68JXJJdhePB4bLtslf6LeTNnCMOhSj1Rvu42kp8sKa
MpHQw56poMtYIndtuvMFq2Z2j2logDVWDQW9s5232q0B7Bhc88QJer54pN+6WA3boSzHDyTNcT56
ge6732yr43l2PLPdHqndPQoO6AgoroGAgw8Inz+rmB2918h6hIJlo0yAKolYcq4LJWZsm1nXkWFa
kUmQS2n38SziC+yFUkINI05mGfK/8Xfuy3t6Su1o8eM17t5poV8Hn+Fj4pALfylGjt8GbUTI4qwu
rIbaHikROZsYxD9OpQgGB90Q8eFaBKnfD9NlAS961VgK4ob4M1sR45mYKJ7/OcJ8hjAlsEcvMnwn
xBUyPFkt5G8nIZx3ZWmpvOh6Y/7DhgPRgebqysgD5oSjMqxo3K9GgbQcMqz0vMRyXHZPIFynzbvF
pMdLfb0ViqslzxxIdoTQoiPjHk48Om/LhWKkFWn7YSIpdpygPoBimt8UBwh+6sXzEWKsd2hWkMcY
eIK0SQWUyKDkQNllLoRsF1WXdopqYqGA2gNEOcrb/3BIih5/oYurLIjPDIG6W3RsLta0GLZXwrKW
PU9j+ICMxooVCPLyZp5zKfkLM6EulimVx4Z+08qqwuaZsXnJO+emQi1gQAmBdWVSvBCB+915HhmX
/Tmuisst1l6thqajx6HkfzwYq2pcluQWyGCn2HghDkLw3PbzqdlONXYKAfDVsZMUjPnVeLWAM+y7
XSn0UXZE/+RdN1cUQoBZ+eIKekn70kin1JLUXDHPAHGxC6Fy96qd/BsimuhUZCRSpKmlQGqKGlbX
qlg1iU5bPngtzn0mcKVM51LjTVNVs0Z7iTpC0Ri5xupW2+eLmP5TNsH91jKPWsplwFkErrQa4LJG
LAcP7iqWBlQQbQo6lrqPDoWFRWzVkOHS3ZaP4liZdcJjiDCeH2UDtCYm/uInv7OesWa+c+ideB5d
WCvLlXm6duV9fhX9LPnbdszXlCY4g+mE+e3r2gNsNB7bo430IEUD6cg8ZK+TgX5j396gDevKRvdb
73lM4ZaDpnobmpU833e2GgGErZpeygVv0zo8qhppFsZEelj/n6Whd9Ig1PyEP7pGnRXONMkXbBmJ
4GhLZcFrIPZu2jOeD6QUpU8tGqE8pqih4I1kEy5UAsRpAxLOvNnlWXaRYsoZK8nZCfIzudm/EWk6
2x+xuRYOC55KxEbmWUZvEMOFIT+gFeWn40odRVmSLX4Cgzd1UvrhHcg73fpLYBi1F4JZ9/E/iuz1
LZ8xfR0yDOEzJ7A5lv/a4z9O+tyzayP2CX521L+GkDzk0im9t+UjXUo5WFlPp8WdESwqtDR2Hrmi
PORaJ25ipC84gYPHjYJUFnG/x7n14VAGH35Qtw/kHVyOcare9t36qdLB4Wt1LA6121L7GqRd19Mk
LnmL8dvqjAZ3AotIbUQg5Nkr6adSu+l9W2KdlLOMMDJeU/M0daoNOgCScnNFHKNCYwsCail7EUID
j6zghOF2CpBIJPg7rRs5jBYeQASzO5OTcl+IILddsNBWYFAiqEsjwilZMaCqk5GxOAfLbazFnucj
AHsABZQYbll50Pr23jQbKfFkCwpl2rCoG7hiNZf9wosl9In2CN+srGb3DsNrmkaQFBrdaasgmWlO
0wLitgEY/bFZy3BiQ4+o522C3Ega3ve70IQ/p+C6P62faUMlFErT5PLWF6OYLATxFAbg1Nm5blws
VV6AJcxG3bFQ5bexltm/xkpqnlsz0Ka9veFnT5j2r38J+DD5Hgt5WaDqcO/wYCIWQ3f2lgVcKCIu
RM8MZbvUtLz+u6Vy1Vzhq28ejwJNqdcPEUjPAqvGE00fVPJ0rhWgJlPavRc5O0Ya9GWc5JiOTyxP
iEbt3FlkAuQE+nhha/FpCnX6AZWbj6LqEbD3KaUEuWbQU7YB5eVAOkKKQ4fv4vifUtn+D2WOkl22
SDP2QgQ/auDElP64cPzwHqpsS0mMonJwB30j29jYVlfWv6Kj08NjHr6r7a2Iuzigud6xwgfU64ts
Lun7Y5I7A13EnSLIj0Wbhs5kI50dLxA+wpeC01WcDhdokW5t11st5WreG6ft+krm4NnEu1og+4hw
gjPV7NvozfzAhbpEHs/vGVYnmeRV4T1+Lrtd7o93W/DAL2qJcON7/YS0cIhfIyoivMHkT3EBsKv8
Cjwfvo/ipEci1WKt70eWfqF715Y7UWDuk3HLl+Qw8xW9xD2BCy0Wxqmx9gXgKMxbbALZoXmhxORR
1amXwEiLMl4+UtIrVOyTx3+oJ7J3oIoLI9Ae6FiPZY5ciGoJE7ToYh+87b6dnhoXDUQSU8FUlH+m
ZYk5+TshBw5sFaSM1PEhDT0ohb0t3yeidc4rDXMzx4rHaRIqLjIhFrvhTqemfs1ZtJrd9NWT+6Rs
vww5FzvIvQiUQJ7IeoUJPIPkcCz2bQEz/ghNWL06eKHuCVhWwPGRhvZMWc1++HWYgxwvjYSpjxs3
nIcLKRPhPPiWikmSLuq64HIoJ6+S/b/UuRlHH1gCEbjEh1Vle6EdIDUWQjR2IeVSGND0TUO+Q9RW
Wz488a84ToPSh3Zg9KGm8KyFgxZbVdduvGjUZMtRA6YHdp6G/eW42vMxYdqTnwggKT8T7HNqPl23
otWWEUALaeTPMPNwi49TWnhcodvkHRX5uMcsO6BBlhtUz6koOdBXzbUrs9+xkDmDMnKhuedugEJn
o50QgUSpAJLDMp46Q2O/ZaLYl+wVFqejHtDyancuB7tBQSvBGwMb4WS0hnPPZOugkRMB2g4qudxP
CCiNCXQr1U9msSY+xU8MK1SEvV3ca4LaXpCMzZVyTO1SvwBVYcSBCJljcRqc2AuWgCX9KU5KirQJ
PFYPqWWLyzfKmnSRezcZ9EDYxJDUHU6HVEJEMQcOVGEbpYaoSzRPuoGDZRulk9G9DTraxI+z93TA
XD6SpjFuZzAV5c02XupbbM9yZ1kSYEZNXMZ9l93uXB2xmSpfWHzYmKC9t9BTbYMLM3522VCAe8xF
kZnaL98DF4nxhGZe1U4P8SwybD87abiFL9fHVsv8nzf0xuLBUFof0aHrW/piwDfxTMqRxvqnU/kM
JVj8CVdk8wiEwJF9+rlkxmBId7LxbgqFb5EDwFyS1o+UGV7AJY3cnT5Go3DNOV/X4PJWF1pScnrI
+KRuqNdbD8oIv+NkYoj5kErV0KDgaGcgKh6bK3z/DzemNlXPLQRY3s+pcmQH/pW46dPLbeSUBJRa
AGKAoIxr9Ogjwma5EGKvdVcrBdeDtf6KNWrKH7w/mXO9orjDLOXJ04DgEf5OL1+4YvfYkBePt/5r
D4FZbseiMvG4cpXrdUv+j4PGdjB7FQMq2k4gRWYKnvNR7tYQT1OMWJBusWL0uuP/z8TvJl0cJyzb
q20O2WdsgYYdCf1nhF4HK+SHRDvVL4DKZ3obkGFeNVfB5WCQKabBZPsdIsUXQRDlIc1vz8ssSaBn
P7EZ61RNAwMOG6kWanW58n689aGYKdtZhLBAAoTwe3rPhJrFXI+QS+QeYdMXwNb+Fe0OIjt6HZMi
08KR0rhI/zVmaR8I2rQgIupa/svG0R2RQNxwyPE8zS4wZVwP2cfq22zwygi/Mo8hAS0SmAdagyrm
66xf8q/TERG8coxSsrZmljfR1+obmb/WOb8zYvCkYDBRXA/dcNTZMyqRGkZIRzZwJm5susCchUXF
3BsDpm9XpWhJ5TIdYXQS+TGXAfwWxnx7MYCM5s0CiGXa1mXJ8IRFxnBf34ZzGv1WyM+PnMrfVNiB
Wv08cNvLfHctt9zgxu8DU+4m0xRwqOVZI0kglxdYt3ny2/eL7GGIs4E0zE4qr/gSWWTCzI8mQhLg
pNQ/BUtDYXUupG3reuwZUp2tOHUvpdxelbqZTkznjGFs2o1dkmzEB7P6YJAvJH7s0NduiZsKv0t9
fb83ykcEvhtDZvx56Gl7nP21afsTtzOvlYi8rbveJfKcRNFoXB+qcsV5vmAgCffY5NqaC8nfyP74
JBOogsD+deN7/J1fhoqnCBJxouLwNm3AHxRnL8HKTVn4OtegRQKYxpl0yMw04JIEw0mfQ6kAa4oB
5NA6D4gRSvMyQBKhHYeFxi6iUQ4YvS6zanP1XG9Zcw9maUkFEpQf+mRDmGerqK29+gtvaqW1i73O
e90+lVw9baADQoiGqUK1yvjuyXAPElYOxYNTnlpDgMZeS5ygMg4Uo4jfyjuwmR8Vz1XoFLfMFgmu
MC6cYX9PbpfISoo5obrPWo7EnpdC5BZgEv32PJTofSPM1KNSX6vlwjhZkxNi52gs/lFWMyy6nQUw
OcE7Ts9skiOnB5BNNnN3dk+BFsPYEqHmV3aFkAeKaWrdelQH+myRAELFZXzA1HOGQeHN+RI2tdyF
VQ8hlOf1C5hOdD5f6dCAznpWVI0X0Kr10HTIg4eWvZThe520thYQdvtTJWnXgGN3CfivMAEjSfRe
lq1sbz2Z5sXOPW9ypayvDFRBO50uwl01rUDAVdPHky8N/vzXSb7N6snzKDp0bGzRFKrdb4BZ4Dyt
Ckel4dkmRTioeqoWSOacyfab6NYDAQauzg/T/YI5qloeHS/sGaqQX3oAS6MBTOtu5YZv4tYtf6L8
D2BDvwxwzy0bWW+vFqD40XFdmKDbD0gAQCn/HSGS3DXH2UGLqo7fWNqkJ8cv3v1R9QOu8cmxnGsQ
SE3tFVQSnc4rGmU7Gl+IqoE20V87B5B1Wgst2ZiZrQaXrwekqDJ/6e9KLosS7+mmewczLunB7e/d
uEDLZYpvu89Ftua3mSLp81naatKwp5TvGp1nRT5ICTc7aafmjqaGHNVryz04ZH66/u7n0I14mQQd
mBje4lkAhlM2nNXkCK5EQN5Qm0s78x7fSuEupsdUtYh3EfiGx6M3ZCzfCkVNr0fC8c0MBfZn/rvE
dfA7l45ih5Fnw3QJUNnWRyZKi4w5JK3xBbl/LNYi8JrGAgQRSYOc+6fuepNUuEplQ7KmNv186SIh
S5JBe7mzxeASQcZ4coYtO9ji5APhgVyvslLMsC5WmrGu1UaZFoiestAJ/4U2uSF1TvWosyTSMWGg
689U7CkK815626dPWwthuFpVEBDLZLtdUDmcZTlmnM9nhEqxN+AGiyIp7+48TKjD/MWIaz+GQGUs
QkuZij8wveaF0n0vgnfGtOe/QIRdWIPolccGnc8mHEFpn4Zni8AUANOI2SOqF01VnKXe8fdpAdJ+
3637DUAKMOOxp9doYt4frqNpaKA2hWHR58d9DYIv2T91zUkHweWvlLo2xdQ/wyaJ2RWgu1TB1Y7e
Rlcc3WQMxTP4rQWXH+6cjZf8ngcRS5ji3gSHCp6oUdxTtA78Brm5Bh/cjZRkhyu8aUfElDpoERN8
XSNW7zHaZouR+3TvSh04VNi8DB9UXMBLgk7c3etMEvAycmxLlUUHZPOJBBbO+3jl8UKBdGNCbwim
yyUJrLNE2ZMHasOfZ+LSpO4v6S5l1FNYwLu/6ZRxAHmR1cRQQvlkj1C6QlU1pTseB4J1IWEB+4mC
CaJrFY+Ny/gZlFZ7EqVveCWkH6tp5B+S9iRRqHnywn5hzI0wd+OAPRhMEYNvSn62voJxwXi+KyFd
IhMLJjaPAtp7cb/OE9BuZ+TdbvUHgwv67XPvW0pvBZ/SaDsa+QOzOu2E2neBzeFyc5yW1IZMwynM
T+syP4cC+DZ5ThesWJgQzv41UpY7/8dxbDn59Y3GbBVLsKg/PZFEOCP3pZS5ExTMtUqVsDJun8q6
UFqGmXqNoU2ED7FgZzSZVnPDbacIx6ZOftTioFjlZPzpFj7j4i/lQqnCXCmd5AFs11RBY2rH2Npw
VeuxR3y8MRvEoXnoXgpyy5zpRte7Rk5k8/s1GjZ4Itk3/mguSRJYIDEBBwgimztMFIX+ZcaD+O93
by3NXYCDMsZvTa6jp4aiROlLqu5YVaWgn47HW4U7zY8dS5aPW1wpdbFAB6zjZDgm5kAgqzjWKWCD
sWDwKfs+TDdztYO5ibKghTb0faUTun0oimEnmTlkHiXIlDuceTZdouSKcg0OvnTN+MA8/uFUrsQe
CU0n8OmmZKNjUfMFxPzLpAa/tfTGLVivHYjsHj1MkSuq02Kqa2PO8vazuAHUHo13tryIY99w2Kai
+C71DmsdcVZzMlqBNXZHJn88rChNqTTnvh10316cV1CeGhrSrCjN0tFuimvNQVteDSa8vsaWO6cq
ASSJIiJjQSCAv+4Gh/6N7cY+aoqPgHShBS6IYDSkQ3Ukpm9JpazibHKlRT6OGlrSS9OwI/R1EEbg
PrJhBjEYLFfU55uMO//Jz6lzBSXZFA+uviFl4paIwrS+bBFaUDJCzMOnUD1odRFxbPCIE7nN78eh
ypPxgTyaWFEawx5lLwWzncO8jwv30mB6pFQ9virgO2YBwbFQT27gVgXEhFvF6tej5Z1xhW4C3ZYc
eGaxvEEZqPdG/yC2PO4Qu3JGuohnXjH2LZvPssMCJenQV5R47rBQIADnIdMGbPrv71RwEdFViM9f
hm1mtQ96U0fp5eOaqGk4ao++rlgTtKsS7yK/jXs/t0PmmXl+3/4eJ14d/AtfMyejXBG93hvkVyY/
IETI1YDZ2GDKx18t61IsACsUjrHpvQRvZNx6+Y0mm9uWbM1X1yhlTZO66pVp/1NYkynh+RSl12Zq
WvBuTabq2tb0aD6hliWQ0ckdhxXo/FVFLXEe5IRwQd9tS0pvDl5g2CpujD23W7fpbMWylZQem0IV
MoObu/qTu3eJJdE9e3PeIfy9QHe4lnVd4oTxkTZTLIEQi3GhIsgcMuTzpnybrt9MVNrEhhq3UR0E
xxReNRFj9EUD0NcwXxTcqNlg3rcP2Fcq9vX5WiP8ymijknFUHUk6eFklu75u1afLICp/hK1XUMgs
GJXd06ogVEUeLQL6JJqti9BV6WDGpaZC7ZumRGNGYvOz0fhB67mHSbzwlvVMs5GimfQuRUJG0iR6
SRNnEs7ZvC4/BShVOdARBEQOyPZ1OHFM/g3Zl1CYeqIP8Hk+7a+Q7N3qyuaCX84sT/Fn/wcyrrA+
oiUbROrHC5ohPqbmfOpCaxZGXPCAGiCXe8+hbDXGQcKLOysFIbs+elBFp3RotNEVxIAgmXPf9Rr0
znt43ijYe2LBl9eZc23oqX2aSZivl8Oz8y7ixk2b3SXcYOYfkzX2Ax0x5N7TmGYS/zphPUYvRKSt
quBUTJV6twtgx7rAffLiyqxPzy0gw/tdPFbQWWNgKV7P+dx0tbkf/wkA/JMDOPTCW5LkovDs7HLk
3PFz9fIobd0ehxon8vxwdNpqFXb4/LSHYBozyK4/4a3b9eIDe1DH4r7OXyMhYav3t4Sreyj8rAS6
GBGHkkdSSXdQpXFncYm49v6GMVfc/BaeSm1vsw34nJztvwxeWY+drwFuBvBzgyLdXccLs+h+46Ib
HfyV+QSd3PLFaXblVQ/1v5fYbIMxqVwUpLHFFmU7ytLNJnUoqpLP72bDFNyra/STsq85AAKmTaNB
vyDnLsh2C9j+xZY3R8zqVH1U99Wxi+PTP4LLLvx0oJPOdANi35cX9vD/2hGmoIo9ZXUAeZbCBEAG
GYALVl6M0VzZGO0+dtz5Mtzjn5Jub4HWrJbMYZa1FfjKwksi3o1WGG7m4+fiQDeOxzV5fzERH+Bw
eXv1w05+wbVO12jt8JSdZIiRklVE1b3kajlKAdwdUg73SL6lhtfnInNXg6hnknc9AI4MQALE3p8i
RPLyCKSRkddHAsfxHYGHxQyxDPE5kiDP5qZkmfO1SBzbz4cZXaT7J8Z2y52Dlo2VnXcq2dW0f6YE
jVI+bGthDMdg9KhCjc1LOhIaWGTNJOFREfCQnE8DcOQirihcQyTKSPCtXskUQpUK5bJ4dwKFFlG1
vnRkXyQjOCx8QHL9D/8D1ZCtuht2bNsxH5W2bEJyshKHQEIihbxFprMEPKqVvE/pki0S7Qn2BPlJ
GF03E+c3OZklN05rlb9cr51SnY40oVhlM7OAxdwysyzSrkkTu2mXfl942ULb+XXS3K8r0lmppW4O
zO3ZkufOCfmWu9z2fU+lyRDNTroyG9ly3AuSGb1rajrYU8FenZH9bbxzem5YaH5JADTjqMIz6hqV
xOZF6+QQNL48BLBSXoxIWW4zyGwYSBAoojFdMhx3+B8U+sHcjHtlL8TA9Z3ZBoyQCv4VNxVwfz5y
DNwAACnw4FP06DeszIwkf4BavdxAAj+sVhulwNc7VmdRCSxpD+jFt0h78XMlHo9cSNCJwifgyuCq
uvU6CVyLMC0uUadekXSzDrNG+Jjm+OVYNpdXAGH5B6/dJo4dzRfyFXw9OmLr4IeVhKjkIWkYB12j
RH67FqlDMc6KrrPxupy+mkjeYYUnTAYuXCSpk8x43gOOkeHcC4LVmCwLz/FCbx7mktLp6wEmnPkb
cRk2KHQZSWM6/HEZQd551rjp5SCZI9Kdwe7P6PMv/0fXMZl4KLM/tve+2dp1EBP0o/z5dDeNs6jC
2DTVwnNIo2OPXpfgb0fu5XqCpoWOF7XOiuZynzYoOsUS1Ldpqj6+aYqyFfLB3D9NRtJVcN8r+ung
61HA19itcu3M0uOSlvFK+GeHc/jjST6RKrDNywxlDKFWeokmkdq5OkALcpWr2jUHGvZXpnnVDTUj
qW5nW3NbD/vKnea5tzkgDtiaIN6VyT59tptI7FNQuW1TbiTWSP/IHVDjYoafljRB6sOvU2/cjtNt
r2soM0g5pZJEmGXuLLo1U4hJQd+irZdHvX28ntqXxpQNPxs6fN/9puizLgqYIDyGNEz6xTUKgLa7
sIFm9HP4CxmcsNI3P54g3fkvyp0t6380xbZ/RcFu9D2QM5U/JHlK5wDrsoVUHqYyX/wvd09FuVVs
Y2+4tCexHJWDnQ0/7ZGK52CohjNnjbg/PRBNwAnbBUhcEf7/UMRNgmF9zNI/37Gq8sk7hOmHC3+X
Fbc9yPjkq4SrLVVh+1dBy2T/xxRjpuFbM2rNBD56LqvN4su/oNa2P84JaMy+VzMpKYzSTTyb/tYt
1X+3B8FHaLwXUVFnSPjgwUmitpylQ/9Ep7saTLFDiC0Z/d6FEhl+bILJno0im6VMxTv0drwX703G
PTKK4qWJm1UzQFta07hpjusV84UKw6Q8ZR228eK9NTSr68y9JjcsIK1nmybDRgjmcmC/8UGCw2fC
z1Yr8IQbCFaCcymiDemZhsxDmYjKMQ7IMQA67DjirCDz4ntVPAV0NABatlZs+Wv+xQTDkpQ7rJik
T02ZTQ5+7VpH0wfdySfjrloGuUglr8CIM5s3StO/v1Kch1vNhqAji30V81VZMn8dsE3LQTck/+5b
frrokgOGmyP8qQ616scirVh5GIy8EK1V/ds3rhhLGqm0QsOWllDmZQQew+oJ0oyy2XpN7fo/mdcb
RKX4eFTTTSjgndThZrEhhMGC/HH0p6Yq2/rQ4kwR/APb4cQ0DvdUyczBqViqQkhmhOL90q14OY8k
2i07KcAgQAxhXjnT4Br9B14RH95J5zk6nsLReiZB+y0VfCn+zaownpuGwSzwrcWN9bsT/+lOe2uu
VIZkjJMNDpvqWUJIWhqh75sGdHBt7ZKzG/knic1SIwFNw2AHjWLLt89vS4qiqFF78Tv1xiJ2o36+
TXlfZSA92iKyOaEqMyzP58pw9pfMM6IJ7pUY3bLaeZd0jnsv6u9PDYIigQldPm7Wd0rk6RYqe5cs
f17jDJS9bHYjkB8J3L9hSpbwiWXA7GZIwIz1W6mfpXfGQODzygFQUAeLLAwbAcfXXVAlSloqTr2D
36SvgWxO+oga372S872nwsIPGSETFV54eI8PVkdh5KNeKtBqrTGWWXbNB5DUiZMYy3Jttr45fHTc
mqqsk6lOV59AATh5RQBQ3mfwyA9POvMDFnLVcP1/Ee6SvHlCSz30drRdWwh9WC5XkEU/DemJyZEv
AkVWRaFN9h5pTNUI0kNW9V5H66MNapAGa41bmgjCg3T6ae8nZFVTEGS/TqjZh3hJBE5H1F+qSBgU
6OY7g4eaP3eAL1FB45N32mmpcVoCBiXYdsFJEr481k/gPZdKh8heLRkmQwpeUBKgRzJzqPmQTA/I
3jZO2pCbZ7hNAKFTmRQq9MuQe+Ec9tuc1gMPqf0JOVSglnc9St4q7RueE8XzYBtzouIANMlGLbM+
KupgjOHsw1O6mPUInqlB1zU38DBBRGGeTliIofbZUQM8KJam8graKJr8vZux+zOODsZi4OzMtUD+
42+cbwbPo+rQ+NlVXSZcAb6rGOB8v8PTo04McxunVqoyWvfIR50W6MjBvlTyTaKpdspHJqQRjYPb
RI3UtuxV/4CRTggapEZ0wywdMH6yL1+QRAI1hjR8nn12nLeVvf5saqhmEy6xt533Ner3LNuO+aoB
FABZpRH974t4w5vvekVD3FVjYD6yzohWpGKivhAeJ0MbMEsqGp/7Pmyzp+kgQG3nOzqjv2km6uNm
PRaCcl6Un4LGbim7Tz/BOYDCdHfFqBig3bNNV6WoRLgTFS4IV5rM9SW0U9s4iZT04+Ug+1+T798K
KM/o6uckzXb2E61C8fuEHuvgwjcesXvjUOR2fZs+faXpD77K4uL4qfUJYWlM5FRFoS6b4RKe4JPg
g0jRROeeG9jswEyDWTztaIpMTsz7bntvkIBeb7JnoLfwIc3YUdISVk88Dfm5fA/bqRW5bz58hN8s
/MWw2epOGuLsxswYNEc/kgS6FPybk4JYVNCfMhKAjluXp6R4m4pmmzC2R1ma05L8yxwpQuqAyk8b
SS08m/dqLbBZWle4s4+btWBUANRZmj/F6zAgu+zbBybciympSeXmdOnQPlWX8TfCBKMr5Ys81pVb
jvLpvEcBAu4xhSS+neHdgRR4PKKAAkzsaiUk22lsR1amx7hfzk64fGBKgXVtFM9ZqZeoei7UI5ma
Ap9thWUIGOPIs5N74XTxIQRKQ6UPr6IYqezhotTPPKhlJ9wGEThmrsHFpTQHMMHLZvflyS3VhXra
RpMZPgceX46QUOeBaD9m6s73P9Rt7kMtHaottRCQwwILTvna+92sNBnItl9grAjhi0lywdex5Bfa
nJHhqkyEfEVCXR2+vCi+8wKllOJ41gvYerFNPiATJ3evtSztPFDJ5ToUotejDJOos4xDF5PJj1sK
aM8BW2lmnl9mM4gW3I9flZ8X4tNjrZBBXuxnA89mEmvMtNV1WPtg1ZejOHz5WxWcSPXZnBTe/bI5
YGN3GA9aJyMuedaCdVmPOBnS2mSWfC/eAuXB9Uh14xGwV2to82DH4ERnvMsWgvt6gnBF5XiW571C
lyilgNaQD67zHbR/dIjxSp/9W34Uqm6eDTrGOcd9SfDmEQOdzhoLCUdBb17PS9gAdfzWoZemvdfM
SqdffTBImZeH1L+95GYVbi0uM6Cv6aqFYpGDmyZD9mVwVB+/PbXkMjMDTdsGc/o0aYS+3uPWD4bp
qaWY6ILDFMxz8J4YBlSicDuNoqtxNX/QeWNnUSWciq9nANWUBnwwPlSe4UJepd+KylavIzyv42hZ
FCcVNKT8sKPyl3LGehSczOj/BAdEYK6iIHAQGUpUoUq4HxgjkSj+o8Wc25x4MEuFFjBFbGW0OBMT
WnEzjZDFOIcAah8libIaycQDzbMwKkFtLhp93L0+iugSp/R5LiMwrqJDNNTnO9yHYyDam10WOdbA
aNHDLLYNvt86N4RJnnclj7uYEajKe6XDxBUFS/6yHC1YfQWJ51LzR9qpAbxIBD2oESlc9Z1CUgy5
aT/mNbKCkdwSBaIiEH4CZjkdAv0ScVrRpvOovOEnoLAYILeMuLjT5NBpAD8RSEeQ+Ytkathvtbxd
Uc7+yPrO7RiYx7OoC0opKfH+fYN8sHVXE16wDR6yny2UmCGtJNH8g1NS80OmB1gW5Yt747xuLI+x
LYYjhk9lxN7D2t+/Lbtn+mWtsg7o9PZUjiupCUVECFqhDgbiB04LaWhKJumJ64grQpG0VOM0Im5J
taMUFTfGP9fd0ycZuj+kNyhOJz4/7iAMI9kniE05F04jb7JWUOPvmEn4MIS9e04RMm6IouP19rJh
hFiQFNyCvYoCYiNfwLKbiheojbeWrhfYSTAzWQ8WmnuXv61E0ZsTApzWLawWkQtetDYXsG6PnNsd
Ox8kIvCL+qU+FjrrOAxsQGwCsxtjgi8x/zkcsPzmf7x+OT0bTTtV3NmNqnGV1EJo1q+qnDPDyYdb
rc9EbQmIQmHEfNU0s1gvo9tovO8o6rcfxs8QP4HoP4obVBSPgBC/FAEbXAn4ZbeZV8kz8ijM4VjQ
oG/f/JGfD3snPsMkbArJoFyTikwX/tt2HNU5PcXRLA3eNoEZEtlMXL9RHsS8EybNDaW9qKzf1Jjf
Ow99zrH96c+NJc1WoeMNbnC0QSM5dUOO7zxDZkg2IMhtKboAJpmnVxAQlJG9XQeaLDF8qmneBK7R
so7lgaA5FFNGlsaMJUxhlxs1aQZ5GPt/IynFYpCu3WzbUv8AcSp+ZnMTOfAe/1ab+GpZ9OVlbEUu
T5Yc+M8ysReiwQhIBZtqqDZgZp+at29dyYuBaCdHnMBaLmacYZrDu9lMOjXQ+tZUjnzqSP0bXlUP
PXPQrSeIL1cIXhuhAe8j2uO4CheVSDvY2jjatOKGFxC/3wLuOEcjjgL0U5NS5nc/XT+2IBvVSSUY
1WmSfjMD4CZG3666rn5mI64PyGmcJ2ef+soWsLvhf9YD5l9FTNFljO1H5q1jPbRlaHUtU9CHvjJF
UZuN8euvmoILDBJOqTYp9VDQEjpa1O+g3CGjdtzWvW19ka0QwJKFBOgctnZx1rRxxuxZL4l18iD5
+uZ4C1LwETZlxyDOQloWGxBvzN18m7CTeIcA5DuSq/Oilg/8u604VJEBurrVqsXMQS6QYLmc7gM6
HgceyrLAo9o40cPfyH4YwJyOeUtMruT81VtP31U/LZmwIC1LqmlkIZuuXQg8HNQDGxb1OJX3A2fJ
0dnY2xm4VxmpET3mF4OMPIIKX5wDVwy+tCqiI0a08FTqHZiYcvFvku4JGIozM/BjYNWaH7I+cpF4
xT4rgrqwL2kCccog2p1QvvqzPzPpYmoEOUWSaumKa0U2x1iI9e2XsWqwDRHvsY1BRlsdckCS10zg
OoxzetSljwoMkbabHFEQUfjFfYI8cKspRu+b5ZvuB3xpqPvrQJJsLSK5cisLW2/xnexIciH0zFtK
FJD9LcHkffTHDl5m+Koh4MRKDqS7RGYxDN7FHuqYcgF6BML+GNV7TDn/kMLbsiLbiNXoeREq7Q+9
pky3zHGNnScz4Zm3VAcNyFA711q1WKRqEqMmPpy9ZjFDbY4HkiDaDwZK8Crlt6sc0RJR9h420vTx
h4BN9oCra/pEV7d0F5eFNHGKReLNlS8bprArUw2lpO2pS/y5OemQY2NmizdDWZnZCEOFo3ZcD4c7
vObtwCKEIqMkLZzwrlQfGlJD5vrArEeL7ZWgAWP69xEfrxeYffiwpH+AV3zBIIm0iPQwDb8GvL4Q
C+zaNq/DNLfp2CXVXUS+VUcgVhVU2NHSP2S1Ci9hsQRr5SyL4fzUhaIYmnG1QMSccpSynNnCFXo1
YZbN6EUkjBlIf21ElfIX92IovtG8E0UpTd8tFDr6CWH/cOpzd9PBTeRtDZq3HU3ylPvRwJeGXwfq
6X5+4wFLXkatm7SzvHTJoNdB8/wZMF7OPeS8+riHVsbz4MlLLCuY6HuCvegL/hECDY6nTfmx0ise
dRDqPjgi5eK2RXuwg89lbvWiIwZrjNK0JXRCCIOQYWZzifagbv4QEPCjWuqPa7SjLFgNfTtw1aDG
hS2777JsNV6LenB8tAAmPkPls+O2xFEq7FErdJ9TZl7VwuqPtcg3GhkuUrz1RjU1pLch9B6MarlJ
oLlwxe3fRIgh8jf8JaRnHAUo8qVzb7vAj1FyfUzPdBKuwHYUUVEAud6a7YotTXHp/rzJLPThDceV
wYhQqYaAofBwADS2guW+G2/VEg80KOS0Sk7+pLaNxSC17jCEyXaxFjZ8yIhjPtvkQD4Jt4HO7/ct
o/46n+sRTCYkGSkrr4fML6lqyqqfUHIi5O7pbxRbrXRRje2nIE6rnxCb3LqsnAGZWGbk5rPjIrg6
z2gHrLTYCl8XtEj6l/St1vIdu5ogvnZdDEHIYVR526/dA2ui7swxTrUOJFDmqOP44g2VHTJ1O+5Q
JqfbwE5Czk/9MZzgi/LDuUmr1ONzPZPl1RX9MZINNDGPXq2DcnID8lxJCQ2BPJkcTidIeBn19CNA
cTfJA5RZALEWKPHiNKF8XkmI1kbUkKm2n7zegJJFxCpJBQ2hEiqv8sYELG01DxCT5J4DidzABNJ3
DWjO/dAUxq7UmNUkQ8jQxjVfVOiilSnet3HU6TkYmDB1R9fXqf7Q7nDKiZ9Zv5b5sz08F6xK0UQ0
CiJNbUgZlmukAdYRMUzcrPY/A7Qi64rdrKHxMcnqW4BXtfbsibmtAwgEZcFYZ7DHwusLKefbXobf
YQoukpWPPCD9+x6aPCsDvntyUJ9rF2jaZxsAo495tWnS7yzjFESRqeiYqpo3OMlvTeM1O4TnmVmp
BTfdk1nH3O2pK83GfrISmEiXBRZ+qMYRHreVOMW6UW1r1hF4vhSd05RuTOklWhN5jGRPymANvgK4
6FNMA1r3me9jm7B6kq0Njqpvdv6ojMjOwGK2orszvPch8f9oU/uGV36skb+x8aU6EdKbgEsAnVKB
iTxpClwmVaGapsDWzTPGn9p3fGLDfT0GIOHQbkIH13M3BqRa5ldBXN2Xoe5gskoaNe7DDauz2jwa
cKrfptwyMLMwrOnxlHT6hdsbsoEGuaN9cC3lSCzKfYlUNP5oXq2+/7oydy562sS2O89dcoqWBfNH
//V+5QsbCaFRgTc5SvDw1kSzfxHkEL6Lew36XNE5NEN4WBMuABcMUeA75ab2gAcrdh/6H97GJwtb
n/Gtcgdh4sMT1OEEWpMaj6T9SCVRJcVkL4Cicn4iqg2WGU/cyTBlgEDlMptMgVO8NPHkC5veAr0h
eMfhuYnNSYSh+/OG3hYtAl7m06auHx9RiM75U9sxDeKrUpex2kvtDkyYmUTDOsCsFDdxI1pFTffh
LKQBF6RrqWKQKuUoUaie+tLhPtHa4NmVHapGlhrYmoQ+uHbz9H17KFKKkeRSUIX6NgAaqlxbnARt
WzNf+oFZQQXcM2/pfeCilHpoNVFg9VewUnCNvZ0lwXmQuecV2M9RxBx99UEV25aBpA15aVKDVDqc
zAHCOp4L/xedGZJP937wRhjX8/tnLU6Okc+MqmjwI5jy2u0XujcwOtpkGT7btnq/uglSDMI4LOXk
oKZoi7uj8vi8VSdXMTKkpKI9ucD5TbHMrxBL3r56DSQKMhn/gnfRHnXqMPg5NsP/UFUTA0FpYcqW
O6QEn498dEnADH2ED9G8fHYbJR4nD3WegrC+6lAeTBwkCj9Sbpw1Y7fmNmQBeDmvLioguFbLXK+p
/Lr/brLAWgQH6Clom9tM/ZBfo2wmtOhNRGXgwbiaRfWUishwDdlhHrNvLHwMm1tw5s14VkYXyCpm
w0VXLfWOw1zFjdDDDQjLtwS13pQA+OvioSxslhKwcRqovX86fSzCNYTcAd3EEUswPv7l7JA6goLU
graaXb7pj5u8jp3njlEFrtWOUE5EDlMWCK12QZnnfp2MwkoCCMv6z3UCId9rMgqf1MDBOm+w2qys
AqBY3lu9+CndbhuxM4ATySjCS7crxprH6B6e9ilnQBr4XCcEf9LKi44LJtYtZSXi39uGNIc0T1Bu
YboZPN2fXpff6GPW7h/GZJA5r5V0mtOxmY2sOgZEaFjWwGQ0A1qIQnKnSaByyETXsSEfh7uozNMl
Jx+IZCTEzS7qJ0Q/8orCXUPEoHTbteEi3L278soyBN/dW2rcnjmasIONezeIPJKJNIWglukroXhF
Q1Ke6lZAgYx8A5iQT5PbyK5E7rrB7y3ltVziPI5Sfzitp/I4sv7Ci7oPjWIOmvSf+l5QNS6AoUvs
acEYtIyZrQCO0z91Z+eHMD1BekpTQRY4O4a8ZE36MbhcT5xmcPFfErIsDcRJlmxw42ZZhksxf+Es
7kJQp/JkrrAdPtje/ZgL6W0fTyiMBBTPXnkQGQxpn0l7xeTr8Y1XgX7VOqVKHSZjFHO/dZTd0pkl
4lqyhgM+DMgtyWp+2xYpLQJGIsV7lkLO2G5EnvFd4RUDoJq40cMxtvROGNfVQhMR5dsEjtsNsqj7
Xh0j1dkU2DSq+ws57aaeZaU1LVOpfQHriccrBZk6+y3FrJ0ZwqdKcF0uo+Mqy7Yqn69bN0TITs82
9XG2MO79b30gydDhMpXpVY40jYV6eOb7rjmBSyw7I8NBGzbnYeqUFRL9Bxby/JWVmOWJ3m59XytH
JUxfI+oTXz9SJ+5PYntpReXlOtFtt50r7IyiGP537QVfTHr/vAiAdHZVA0+tfm+23aXZGl5blOzf
BUeQoEC9WBlHrTu21DltY6aDferE9wLzE6uTCww8Bi3SvY3tQJgocAs+PUJZfMyZrvN5X8JXelWQ
yNZW0N4DGUZ2lAKOLw+XmCLjgXFcYSegA9S+OrUu0wFIHCK0grjoglXx7g7KkfUWbIGPRj52BQiI
cU+XR5LbAZ2Txyf3dt3TlWnj8G2bNZ653GWhRCf+i1UdJxZbsgPOXOgeW04iKBml8aADUmHzBcys
GMJrlhKzGaQQgueUJcaKoLmFuVJQCVSgWKAbgwBjab0xj9FQmpY9inUHwC7wJJSiTWc6c9cJjCVO
tg9ZNQa4klFOc+c+UojQjRZapAidUU/0M0GBgYWALciRitmiIn1XEdiAw2n2kLlamtFJq0y7bY/P
WyMEC+9YyjuTjq2NO5wsxhjVq2tkdUlTAbOoRSw+J5FZYktt6mjw5z9M0Pn0Jqs4x69W8T+CjltN
dHl6N9zGzu99o/pZVCkq7YO7p1UGqIztJSnOhLMKEfM4Z74fCcXq01Y3ymQyjoYDXX9ImZvmsK8P
oklQ83pJIQNA8mTFwBVCtCGUUW5zrIPAuQGGn5hzpAac4rRHFlLocyZXbPx2L+LWEy5OrxJ2n3b0
GcPWc2c5KisYdy25oEYwdC7mVPfoNSsRFGo2XaW4O9AhNCMbDZ6s6reiCLicj8sAAqLsf6RCLcgj
b+LWziDe65GGuwEuHKkI0PiR8gEkhvVYMwQCwTUEMEifUit4Ca8ZOcxW+zCsBSHqkcIzZrFNoFcu
O7nOFCTeQSGGTuK6XPJd9QUf6QI2paukCvoiJIB+3Wawn7zGQKsEY3TAo1v61pbmK5Y51uuec1Sx
mwbCo1M8fRFIwx6y51RrZyMKI8TkzxrOFCwl8xnec+A8ekXJzUGEITJ0YErJFu/P6JZqIybF1PyI
q+Twt9aQDqQTSDv09VMZqonH0RBS5lO+Y3L8qC2cZYPyzq514bDFYTxBXBWMN1tJC+cItQsD9PyK
XSBoSTXBCjIqCSHFYrDXQcTVIVMWcpwT/J+zdM6qx0IYjsIiBLlUcsd7tq49yev/5EuHkad1AraG
+enok6554rV/91pxe89jBd3pDg/YhktJCjL6w8choFND5vC2QNQt88s4LJjKv5jDMC5mRxhkDDu+
d1HE0PU7EPUUr6eG6im+SfYWx8P4FwEbCs1VgV2l4Xfb5SytcWHr4Xeo2qrBtjyGBJJS/guvv5uX
XRGXp8bHGuBx+MeHNZd+zqWDrUMjmYqneryLcrbgfxrQnQbj/eKbwdOsGFwxk1XFiGiRiB8L0lig
2ecL8sBU+LwKiHf3Ba33Y0ncexvUP70KQiPZhqezOctLkZLmS4BnzkyyoqVnHX+bDNoMEWts85Qx
/MkzRtr7Uh1VpHGEpvBWVymHW/DJ/aJP4k3bymeG7ffGkOPvEUqwizIp/8QsIQpWkDTlKzviETtT
s+yV2QRCUhIj7e4d6FFyoKqXIj7FboNAv1c6+FkYovPWCZvoh3ZyleZiPIpL1hdU5Ol70pXVnhUE
s8MNzD2597WS1OGYWSoIgqrfsfKhv5wbPRn3SK1/++ntk7/DdtBtFfmsmFh02R0oDtiHz5DkFNCe
CR+oF27KBM+BSFW3NSRv7G6Zc9VPdgsEcaLPDHVauhVLU8fcJBB83JffH1n5pJ20x7/IR5NMJ2En
zJ7W0N2p9v+1lNepPFCdmHNjz4hdTUmvW4Xb1eoqOjv38G0QUCu18jUOtpdxJ1kbDTe8cIA13i49
spE7W6QoM5xJwcFUdOtbFO4yvitvjeTz6eloLPzvFSuZrMtKHoxjPeKMQoOull9uxZ7Ap1PDpyrK
yNDL4P+yJU+LlMmpDWfElHzj24IwoA0Vvc2FKgNhp3opaCEx4431C+dKZY+cnpq03XBiJO24m8cQ
pWxrT7j8z/mRQTUfUOciaR7uoDCmDp+1qAOmYfSAPzd2+s5KXyzxN5Hnb802RVuDYjb82MmY4QYp
Cw1Jvf3BL72iIovXP0BTTBl8KYC5nGIP+AKKnQnMn9ySwQmUV6DEXrPtJ1gDYECDRdlpIWmAdewr
v5TBPAejzQs4krOaDIKTUwRCMQlqeY76G13G8QmdazJUHfPY6gVCRgBxnJ+u39A7RZ8VEQHL/ReK
5g+Vh5OBPoFYn62FCxuvJ/dsKE/Sc3Nev8nTT2yTNUjt/Bw+qHWvgyDHX0pi4bL4lq1a+yQC6x3b
NG2IznFrx2HGeJjvkrmOLOW2EDq05eG6DNdPwVn99mTqdb3U5NNJ9EImAVNv4qtS/DiRH2Kzjw91
8lmObHhf18XhKKt5DXlNb+8eaEpsktLa1AXtoSbJuB/YcMcAcQ+IYkL0T6S3ZyTxw9kVx3oyOQw8
tYj2GlcVXf9QaxmbjWTok+E3brTCn1d4Y+1uireKZDUdEY+C1HcZZ/NXYbWD6h50Tibd+hz/VoEk
TOFnue9VopWGhCZ5cz4gpMn8WVqXA0pPiOiCQK+8DsPUXHDXOYQry1ndMW0i4iJxPHb6h/73LaQh
8qNWqV36VnB5kGJP6Dy+c+x/G9XPbQfUKaTlxQr2U0Lh4eoPP+FYuRkT4gqr6PIIsWewzrGihc1P
ldI+xMJ87fWfIiX5iDVxK2fyhKpS9vNJUAKHUc2Taql6VTJuuPCjqSe4A2wT3Rjg6VVE+KbDu/FE
CqPkR+UJrRqbJrW28/0DIpcYMvRXsb6nJYhyVMU8HBwqVH8/h8b/Q1cs9ceDSMNg1NGRn3X1ojw5
68I2ke9m9QmAbK8xkQIjJHLAFxyiOUOjtHUnsJ8Jomj/CvS+oTDMvpLvBjHcF1qnO0aHUermjkkQ
ejteAqzR2hU8aAFwyam4i5UPD9JaFQYgfwxvU14uTaF1dZbVKsHiA0t76eLtDSCSX9mXvoxUuDCU
EHJjzacM+kUjvOk1zI1IcMDZnOD6BzjlOCPfZAylVQM+m/e+UqBK89498fgs/dMVcM+m1J/6lev2
i/5aKYpnKOZnq7487qU6G57bB03FySBL2RZ596T6mWz9xx2cAeosR3F5/BnDXxM5EqZPZlno5v6k
ozdIT54tYNsXZB5fa3o8/CDlcfUkbHwj7oOI4pzJtbgXnswowLzQWWbr1jL/kgutv9YcpMGgJjCV
YeetGGxrgYgtDFdK/qKgGF0iAetFPdOQiaWrfL6cHCeX2mfblT8CJuI2wdykBjfcP+re5pxGxVKA
eDO4Zk2vNtsd0kboY0ZembqAM53HIYsXipsr940eb+Y4wQjcaxr16wVqHo4iqcMiWz1j3Pzg+/A0
E2EQ5xHNOjrGH8aqbaps12bNTQPCXxiRX2WmRDfPxyJolxkoRR6R8A3LAH7x4JW4GtD/Uj8wZLqI
uUIXvrIPuRsubED1Vs+hemgkZaQjiUKftxU/tPOC1c3yc46JeBPtFnwvGOItQJKgzNxJGD982SDw
gC1YFN7/dtFSyWH4xjDdjIWlUPE8pWYQ/WhIggu8SrHkk9tMUsZ/wfUUvuch7iAR13uRReD+EyPt
exIReGQBKHXGipCbjOUcoekPvng4sPSLzVvndYk5KYAlkfQRUqNb/GUJZSvMFa2QCQXD9aT+WQ8r
z0oBHYQX14RGVJrgSMUXMqNC2w9rn3BbmvG7Qp1ZAfmmY9oCuTCwJoh5aq+R2dpjo1GuzriNQvrr
eBExe2OAp2LJ2L2gxq9hEthW6K86zZY1Ix/UGDJQTvEUF1T3DDm04KyRwyQG2rF6IDc9Hjx64SkU
C+EvanQxta0z/Gnqv6uOwtJWDXC3OEmDa0ddIQa7QlGLehlYBfIFDcFNHMs5ppcjNRr0p7yJBzW6
+pG29XOfbce1FXvqFEldSR5yfftxCV+i0oyPxWVkUnA61GiOhP1mLvn8niTp9v4Xnyn4ixfDtSQL
nmbxNWUsDEqTCmDOwMr1B76wJ7J1hee+stkEcJqR/7mvMPnrFZzNz1FXjydvgX4tA1v8QchWweOO
4ZDU4v+L37NtVppQuCbkri8UmpunFNZdL/aVsC8xpaZRN9bKS1vmKLU0nvtZQ013zpzaMCCwDhdm
hVoj+IuQSepSR7VTBJAEL5wsNrmb4dHp8QL5TBx9GU/lLYSVojnj78c5/CWmg3jWLo5kpg4t+dB8
FaguasPDonu5Shrcc59q944ENF4OqHLAnsZfzqv3GZkICZPScWDCQ0hEEUBPCYu/eY1UPEhNJdSK
gpGvh3qzTubvKsLQk7cO070ydF8SiulcUGqVwWVb7gneWUrrW2Rf+sfUF8SPLSviSKf1scfpzQBh
iCJlurgzIFJe0XCccukivor521X7ve7D3flFbeM0TKUZ5RcQDEKdCCn160kq2Fl+IDSapM/HrBux
zyqPu2Fnhn0NSYvfLYK3ZAnEMOWcgsJ3hPvFrHXqGFE8M2PWmfHUvjBkBjDWVjbzm6m3X5ZnFUBk
KzFFGaOc7A3L3JWysekMD82oUut7KOoFvTqZRJLVp3QoBaVQ8JyWCt1jb9EoF4gVy9boNrO714sn
Izk2ZDHYI9NbtwHIpT5cdA/k/CNoYCWzDIvt3DAle9z/q80DxUJgW/bUSsCQGx/xYoyGdoUpqpp6
8DT+h/jIo1zbSarGO91BgYD5VhkNMtuMijpNi/qDy8rpWx9JOApCTej7f+QDAkJS0YaxB9uftpSw
66V0N1qS9/FIVsT4lyHKN+VGcYauNIsQk9F2wjLKWYy4rb8PON+9Hxxl/h2uw5ToKWjGJV5tKqaG
z9MVHCe6vEDbGTZ6B5lgWkCRbPojSFaI9qvhbVkCc6QONBEM8wQ+vKAPqKGCVUhtjhBOXXnHePTi
6pYyIpHCeZHupsI9CacExsEvkKPCuNbBzWMKA1ENrB/Qk3pEg2NT3M1PKch1NjKgCxNPeYUJcPGQ
VNZdDF/mwNTXrH2LFxw2MUIkFJKUpMReo3DLaZ1Ayws+yED1U46K8oO92ZiPvjTspE6RwhQph0wb
nI4C8aJfPZTZx0JrmpHldOzzkylxTXloCNDel8YXyGFQBvzh5Y7spH03O+ncfB2qRS1XCNqyqzMA
+Qd5pBUFiNUQJ8tI+sJ9ZBuWp1JV6eOWHOrJZ2jsN02/6k0hiLs1JLF6vc47TDc54jehIXFQaT6V
12p2u/o//tjqqGEWkTzPHTZxMCvDVTF3/G9AqLJR9Mg1wcxz3IlPy0xcSthwKh0qiVhOXU5xpaZn
XYR3zSXzDR3MHfbRH8YLSMUL1k+gc2OUZbaua/+DYxfWiNSRyBCEZ1M0LIb5gNH26y+JnGVN3+C8
dmGXmmoZkosAJpt7q66QvE3t+OEhxDOhtQuT6FVtvEJ9ZAbsu+Povjm5T2o3G76iF5l/7qtGsdCi
kIZTQ+5VpBpB3eBi95j1M1gw/WZ/MpUWJeSK21CV5vrAoFTq3rIRqV5Xeowu1zcjDRBE2BA09scV
oJc9EBHJNS4KlScH13Yz5i0tbJB+4fbxzzfTaCWd0pphCjbFWFoooNiclz7uvuX7XvpROE78mbZ4
P12HsvM+sbrXsnIQU/q6TvKZQdSDQt1SSZORi5eaBAFf0NFrM0lToC3i+P9R07WXuVP517iK70fT
txx3j3XZ/oX+6e8UtX/tb33cB6leB44Ex1l1J4eMTJIlZWFPUVP2oz6lPB87d0OCqqlUU8cKhPK3
fDHTBbdMAn3CiHQS5gcgj3QucqfT7Ha4EwbVtY9f+sPyE856x6+sip8xMkCHor+dDXs/t6PSxdBT
OnqE4AZwSDbXX+d31AHTlc3ZHQo+7iZtCIrmV7DyuB10K20vCYKcKAf0ompv3SVJYHWkPyBqEALb
NYMa3IaIxdZzRpjYJuf5BEV6Ub3b1XxEVDchYyLVrehFW+fSOhAK+s6Eob46VKdSXjw+7oeJAO+s
gV86Cu6LO8KVPWDsOtXZ1AvsKVw1bZj8yzGMw2AY78zSEu0tAB2FeFlZgAgPzEd8hRvB41LuiNDy
bYeTUy2UA9Cqsxf5NV4+VU5jhiJ8sxE6I6WJpVoNEn5KyphUJbsp4NXBoisbQXC+ZO2nNMAUgsLW
t4PE18MeBFxfMgs8+uODNfbLEb1i97pMvunxM1diUA0ZjuBKyI3rQRpRkOsORjALZRiV85Ej7UtM
GBPARgrBt3tFJMdSlOkimz02VYoa+VLvP305G6n14HQAxBMOboYoIW+R4p2Lp8fDe1bT/9nqV6YF
4R1klVhAGCUAYlwR/ytfa9+lSXHnsAIDCLa3cEN4W8Nv5FzE/LNSSNUH5ALhNhGwaKO2uwypGKat
159YpIOPfodPhLuGzZwMFlql3oZU3k63JM6evDvFyy3KCq5yv2zBJzmY1RCJqY8Fup4C7Ak+cLxV
E9toxQWURNkcHZuKFJexYtgc4DDWw8zn3EPvpesfPuEgLJjtQxoJfjdA4GpRw+QC/kvUHHj2QH/6
dkQ8yG7G9EG/j7phky5TM3OE/KDZ8hFXbHc8ZzkNQPR2r4JShFci/uU5ybDuvwXKqmzttvWLoCtH
yx2SXRZmRheWswi1zfA0HbMObdhsh0Nghmxxl2jGvEb53gGl5iebsH+aoBqb/imA/G47iVU+GOgW
VnXJJRs9u1u0azwPgR5CjhDhdQNUcvyrCiys5t8zibxIs472qoxyt3MragkUy9BxNWpuqygEQ0GH
2eEJkzMIsvVLz7gF2kY+Hz6YiKGuo+9zfrGRsITmq0Z8rx65ic2EzLFvCs5/beyRaIgt8xZ/IvII
27X4Vju0DkQMIVY7IqvGQRScaA393ZMsdwNBYkDuLCtwu+7fO+5J0U3EeFgQ2CcWmVLSp8FkAPGt
wJARGFgGkoSri+SsDhEnIezbAkq39uPZbCrJ0UtFb+wDxZOK5Vu7U+AT+owVWdMZslxiMtEb1lkY
APUVqEPMgkq3r0PSZaQX695cQ1qa3ywrxhq5QlzktGYBNZGv6CalkgW9ymUcx4x25+26eV0viPdk
aUlpQuIhba2vaxsJmlOHXoJannMNJlIuw0cfq6rfYaWYt6nm0W7d8Wdy1e93y72v2Oq7fHvq5HVk
znYM1R9w9qYWPA7SYEfs2QTiRjjCbvLeSaWR7p6gHPxWmgCPatfHuKjn0gmeXRBrgxXPqJNUxr2V
KQjJ9N5b7rfA6PtzgbghT8Cx9OVn9FDG4fTb6THNqqG0zAJtItJGl4T8OQoy423eqJQIYBuZEj70
oV579qJSdglj3rzPcHs9XIzsL3GzM+0HEW15RCiwmDHaZTSVJiFxqPeHZ6TIpyPBGtqniWFQYQa1
k19Lb/0iTlT2GE7xWwMaoRMcl+0bMK0SwYnBPLMaqI0QUxCR0nvyZz/a11kejWQ0hGJyuaTPSKVl
7xw6IoX4nXLc9gWH0okJnePCVcgUnb9lKXe2V8+YfzLqvlEcz1ogOrCIWA4JgMMntojhQAd4mnAp
j/dpvnp+SwsERpgl993i9+qO/lw10dBu8x9vdK7ZTbALw6Y9yW/WY4MkISfNFGB11ArOnuanlo4d
ThmPMjLFIOOxuUQFE6E2Ke6vmSIH+ZRHFjyIiwXgBAONd2D7PKHazlXP/Y/aFLcGRNnEh1+ZsDEo
fNr4N786lQEL6Icaa1szifqAw5IVz5daPsMz6wD7TzTWyhbTjaKDjdeK8n8EtXnSt4kCTz7Mh7k3
d9o/14khfcK0ejFxwBXmyteqXsmL3U8woxOqSlKaqTJDvP0DGGvqFUAM8vm2XVlGC8kspDlM44cX
AN6RCmDDk8gr+r5NlMkh0cMYhg3eZONf2AnIKOrwriz1VxyBta6jpQlzS2p0PCqz+V25rcRe8BD0
ONAx8bvSoIwdp542V7JAbvcBCgCkFEEEqxuU1hKYQ+y5vkmdVqqw/ooGXhjd9WJiLFjE09wYKpDr
T9ijLpLB21Bmpu7qK5Gs8yiuMPDzBO0xdik0XyJrY33Ney+Fjp2snly6dseA9nL9hBkMqlqhisjJ
qLed35GALIUc5HNIn9NtoDuxuE5Xi3ZxWv8jBoW/tWRP/uzc/My+u0va6v2kem20yHR5pC3GY+8N
WqLjjwySELKcSFUEPhHeUTUGxDYvsR+mjP3pUzGgRD/Ki34l6WpjXZoPrJJvYnFRs01ChA4aClBo
yIApgdLPCfapMvNv75BzQhQiAOXvztD1w+plmLwA2i2rHDRebuksdw0zZvsEzNsaYCB6Nesi/h2I
Pbu064x+H0uJr+0v9zN4T2mLnHc7Nd07nNHRQEUciAZ7P06pCFm+Lyovmpvi1KAwTpwX0dhg1kZO
4DEpIlqMRM79v88j4BkP1nVugrRakX+xQCYUePGGAovofd4L4FigAIvCS3Xs4aNBF4XG+i1l6K4e
rgniNDqfbIvY1uU0/gOwpCtYxNt/MQftUp5YdiY27yP/2MkdLq0QMTE1EdSxChvf80dcsmKYO2rx
czUIT8dC/0reY70ugj3vX7wZw1tOCAaIrj5E+lJQeuSsBv4rRtOWAoUxQDbRN8lqFMERzfRN1MpW
fF0Q3bK5jDOk4LN0cBLjr2UXYo6ZFM17RVgOteKojU5kj1FJFjBdR5gHj2JUB4+qPTI719rL7nb8
vAS5vmQELLD0zWDTwIXxcewCEt53VilHqvcZ0ClLqJQGkEPMSX9uv9ixnyOWWbpZKMYsF/iTeUI1
MlWxP5RmJxq2C+DIPHvNjicFyyBZRPlAa6QuNyMu1dlKT/FGCbrSF+lLYFO0xee2WtRy7kQpPjGd
I4+VUjy/wtPxSkyjaboMI4syGx9lMZYDohDP8GQNkpGY6dpqXaFzYV2QFfHPsvhkE50vVfc5/AWZ
4UeuupbtCQV/C6p93+CM3hGylzY1FKnZTUxtR1mffVd0XyR8rcZGmBhrbi8OI+qQxfsEZTMVuYvg
HEj5C52Llkv94yYyppByBxnrJQxpAmBMC2UIQJXLzSjDo73/JR4rUNmTJWLa/Nc3aIMjsnb4W4Yq
gkwIHjkRkA8svPa6bzIT2VTkkswQqib0/LHAkRXoFfb7de+jHZODTq3NykFrs3RO/e/b35J8WYEF
VoFtinbMyIdk4atUtCt+HR2v9RCh85wklqW+yXuxyWnRjPK1FJABLz94a+TMHufOc6CJ95GTlvEM
ZZO3ljgfinnns5jYb60tacP3JPLHdGLDOBC0KEb5AjC7aBFF+VCEklgQSvxVyLAqoQb4DtMq5x+w
0xgAJ9daGexSnEPrEVoqMzUz9yr1WOtCfJxiDuJfDSFDhtubgiQJyi4xs9eEeD07anp0UWoq5JiZ
tWjpjsIJK/3SMIf7pYlC97kgE6ssmN93oQeiaCdRaE8YNAwa7xHbDJUiwQ3M8+YZVMw9xdkid8Yx
jJIjlelgoOIbvK4oQytPbxXEWCIHYyDNZ07t5iQxb+nka58L7NNm2oNuWE6R6MqKStjNPjU5sKt6
PADfUcljDYi6w+ZtXDWI/9AvkmcjZfCkFKTsK6TsYmhjjI2XIHWUuOWT6OrX+mRA4IcMyxlTOFiJ
Yt3J12CoC+KdM5qsp/EECA8C556sCKKme6nUdgDDIYMYlEt9/mbdVdCEw46Vcj7o8GOnW8I2Yi/F
k+bccp5hBU3/X6MDLHmMkrb/PwXG2tqmKFpBeiml1y99fZlzhABgF+aYqkECHwiGRbFr29i86spd
JAJ/gdHpngDQ/gz+P8qyNm9WtO1DKAiHXEQHy2Glmof3jxhkRGq0bqEQQ8MS4IxAXVAj7pMzO1wG
WI5Uty3ZEg3nXNfbVPttsi1XDzl6kO8bmnF5x6j6W7VZtVvKJdS5J3fWy9VWAaBnDlyPGYMzxpKX
+hp5W4FFUB17Ppaecm8IVxm8/xqh56GZl0Px5jr8UoXXeiVNzFplNRtP1wEd2SB4ICF5tDxr2BSf
WZjARN1f6l/3OvYzX0lF5DiZx9W2o8CYGvIDShQdhtAd76tT1eEAVXzaR/N9BakgmgVXdmCqIpKp
4NoCmuQBl77AeD6a+DSvy+pen8l9FTzDaBv8HJnZfKYFN5H4m6h1EPL4NMsExcRci8iRD39a2b+F
M3PR0w542/iN0Gwhq16bgN93deHnR5o3yP5XnfqgBDmi7KsZlK8sr8cqtUedHa2Jyq61pZ3Xz2ZZ
lmK+v4vrZevqyBOc7bV0IbiJfNPc4ykmKkD4cOJInSgea/rLyNrpT5iXkGXKDpkVL30lrtmjXDcX
rnDD8a7r5kOzkAyBFugkbGlO/e1IqKyPrb6s3NEfjzQEBKjfN1sMRcnrRQ7Zm0Y+csuqNRfmw51S
F/kwEZHvNmE85epOPZlgB2GWBOf1VlLIKcWSSSc5UQtf/5kkcMEdkCIpNedTavLP0S01XcUw/Dzn
aMq9kPweOeJkh6yWVoQ7jpZKC6VElf2AcmSxpA5cOh17qxOmLWAXAoiDSIVHi5/A7mDk8Ty+MEVD
Cve5C19ZtFhmYhFAbQytbVZ1T/Jv/7ZA4/fQyvS5ij1v1reCmQsz+LLaY9Fh659eKswccUj+xJjA
lgc+61qfmDznuN4MhdjL3VKtNVMeqQpN7W6WXwHR0jQY0gPKadqRBGqw6acos8vXrrq3tmwWQowc
r/uYRyZ//DOmVMK72BNANknudJ1f0vs/wfsHKzoarzCag9j7ke9mIyHT4SryTXTlGVgBqJGmBUR3
fEo9V2W2CxH8LYBwKBGCqXdfj5CLssKSFZpwS/sOFU3B09nX4bbmIbytg6+vv8Gi4v6aI/EjPnB6
2l2bknGnFfDDWsBVH8Fcnn/DvEJqpJzj7WSTObO/igqK7ETkI2tlc8PxPpyJrqf5Vz0VVa5Znhzz
NkfJgM3wwvuaNkYGt+p4jNhVVr/wQlDDBPQfSZ3idfmhP/QfxzLdOn68GPaF+JLeg6Zbt/d/N4Qh
LdL1lyMqKTgfN+PjcC4+nAU6fU4SZ1y/5z+knxXGAWZPJwGGqkEN2Ff6SFoNXleP3tAP5VeY1L9z
NKPTClvYPHz8dRxkIiGRjigzH4Rq5P0+qWEBq8TL2Y6h+V5T3fXgznxGilREL1LayuvbqcA1fO92
ov6LL1kfxkxccCqF9/dIjqA6UugEPCpOHfk2R24nqhJLMkXN7RazaZsezRXvkCBv2zDTnHovMvJs
+HzY6SpgzVWuGG58vMEPqMM8hbX4TlV+Pr/45emsVWKLYCEFCxoG0eBz4A6jjpstj6NSZQh0qsDA
vxzjZSOlR4GDa6Qi1j5pjPFyR549B8ifofm3wx3y/GlygBafd025UVkiNaVkd07EuQ3/z6FmdKtL
BsLcAOm6LZZO3DAuXGFAG8Fv6o84XLBNaWQoKxpKIXxzHjwE4hC6O1KMrUzV4HxLAIwErvHUL33L
6rhXShNwABgND2fw1OFEOcst4CEI8Y2P6vM3dKUjAlaKD7Zet3Kdt1H96wtJzPZ5CacIR4PU5h06
91SbydVnuNtL6tip3O90E2SB4nhu6y4hFM87NXgmDIdIR8nokPTga8lYaEoXRMYPNectV80Ruu1F
twSbOadXX2nbaG4oL9mB4HOg5TiQGStDHhb5o9d+6MwcfCy3GNKWaOyalFh6zcRLN9x3/wyn1mBV
wLlkzIdwAvfoOUdm6/m59cib/l/u2ifi0PkuRUT3ltTzdgVbSzbErVhFNmOKTQnj3n5yrFQvPRqp
WT4ClxtNuRv6jg253iY6EsXHJeJkLimdBRuM9CJkYTxT4w806kSaSbAqJzmM8GPo8vTyDhW3kHs3
lUoPI05ogeP0JOlMLRtNV85SYIbk9tgUwO+1n8S1RNrn1pdvnBbwEBr4zcXkI/oSD18B6vn3SH7c
ljfwAwN0ihDrwMoo/LBqVOnOJYGakDFfPurP7N7W/aPUwgEAUviNhtnQpxRUZojjmM6jZt+8pvBq
5OBxNWVTcU/Jto+U2bZuyoGsH4TJ3eyRMOSm7bkCNadCHFZhMRI96QTCrQCXFdOV4a7OC8SXtHo0
UoonHhuW9YdnknyNgVGYKjh3pLqbNUb6vgypoC+95IGTyscdJwzFL2XKxUZfJaIXEzgKpvoTCYJn
OvNfHUWE9hD0sz/ydcq4OO4kdo0ibMWZLpKiJPQtNf8/mKykJJfHPUp07FHpKAlgbDR3I9SJltFg
ZHL8JKU/3YSCjmnbnjyp+Is7MFWWbXE8k84/uEeX6+h7jIa8TowqrqfJvT7gh3LDgvxDlJrJ1zk0
x6TJ3Ud9XEOdGPTmIaN3BUzAu2xRtQL4UlK+/dilPSIVycnszKyODIL281dMA0v4ovCXJEnj9AP9
6du47KA6GAcTurwnOstIPme7iLlhVMG77eDVKrvMkwzO2dHMgF6xCH2gD/xE5vaEPpAoUSKcAwCj
ddGlZgepF7AyYNFAUeEX0Z0tpJrGesI7dFns40sBDtPZF5X/OtgeEUMgOLi6XAMiKUbAA6cGp2r5
WjMY6Ur1RXX/Oek4KyIxiz4I7UlloDSjls7yF09qkGGsqvx9F63R6TROTt947VkQbT0PTrlf0v6K
6Was2mh5Tj1uGAyyX9pbEoSXznMPLtWgs4X6QD44pyNn6wswsqRKgdbRecVkJFjTFxMkFK5VnIyN
2C7aqid0nMosgdhZlup8U9LJUcdkrsLwlxVH0PbHS84F4COi0ZXGYMSCdVdWV9CfqSXHE6e4ekAv
lrDHKOwe+1zOk2PMljQShKYELxr19pW/2rQnJKF33+wPs9LiNxJ1xRsev4XQ6naolm2wcWc6Uik8
Vc94dxV75ryRtslpp7C7QuhHvtXoGg3HbPK+0W/kl4muByG2t351UHV/Obi3oXK112yJH1d4Kq8a
Tspfy6KqdhqaU5XDfZpT3lBe+kwnFFbZUqlHarnLi3cnHeN34CXJYY6hgkF+kDv1TPGErUZV49s8
fTFxyQtcqhjKt4dmNE0Ut3s1Tsvl/twy3UB+EoFp1keZgXMfmBwgF29uJXqZq2rey0E/d4t1Tarx
iXXd1ERBrYKf7jmPOO/9eoziwGt+3pk8K+jIGZTuq2em77SgGUJRvLVsNEIaGaMWMcjaPA39r2MQ
BI6XltCWovzp2+cPOPyr3Fy0nf6LRoiWKvLAsHij3+kldsaFIYjtSsceYJI9b+UcLwOdqvmcL9qj
gTqDeZ/eNHMg9+M4Qx9SA5MDKTGY1CrXUsxQrcLopFr01UFNnJpVdYH+jv0+TAY07C/9Akol+uUf
IcXpXr2fOPW8A5Fi8WGhT9qW58jNb5WmcnnnDGz8KSUcNyb02q1zFwimSNhGYQFcQwIf2fPqZfkU
H8f6KJOBGpUnRiGMYY6lV1cAIAiA/dXt8m7b8YgXygfFlmm/MWDZ149RvV1RqhATd7bbK/rlfgg/
yG81k/lf+7Z6nHz9bYA5x6S3elUeUlUrv3uTWRXqDfL2rmpM7iIUnvHReFz9oxVvFE8KjRpaKQGO
qEnOrGKLjHsSruQy30KVe2e2xKJRcByLHe6YLgM2KH+9Yctjpj5/NTaFAlikTUdDiI+4q6lnvwQY
exMlIZldoIBx8QuWu6nrxrrq3butilNZPdVbpxM2zHtY3ujSCgw29J5NCKF0wzPSTKD8O/Y19nc4
kLhHPNWNZMRXN2eQq2PIbt5HRMocxmPyh8l5C512aVvV2o43kJWJ8cpJVbwo4JFswuWBkmNuVSFa
cfHE5OzOGhwozvQHZR80XQ7Ygns7k/70FzZTuS5o6prXLso85nLygc4lf33YHyZh3MR7XcNkvdX9
7KpvdZ/71iezqcyLgv258XqPjgPgG+iovXMc1dWFbNSUYk26vXdlEyKWc++ewCYec2yDcbeAhQGr
bGoqHweN8hEzlBTvd2NeosP4GsEnDrsFov0qpieugqfz19WBnyNuaFOBq5LgBt+4BUGTOHh/L0Gn
pCelottAxEoOGJvXrkL/gfG5krEDJL3F0QwoA+T9biLeCCylIOCz+rMSuppr9BWGrUNJV0yUeeVT
Hwof5VLXO02wSTmvcdwmaf9yivtnVmRGMp73Jb2CFCn2kJLDUxWh4DUV0bf/DL0xJmKii/TQHWKD
eJ+b1k+Vt1cHbW+NhMNymwXjmZ1QjhgjCti/FalOOOu3niyEKyvcafY998+tF8zFV8fbQ6/Fgzdg
NP4wjUZdnFNxm0hnjqBs9JJGmVzdLY4j5Qc5N0xuKjbs5xhWsvDBs4OhF/l+oqpwYcnJwSbkgjr0
/odAo5rsIha8izJpTdt72c40/yynEWG1qQS//GdaR2cG306AduD22sVDsCfVnv6aaQOuOjgDWCR6
I7DgPY/au02BsRuOzUkLKH1ahzgPXsnE0EbQPN7Fax7c5VjMp+2ryG+5w4ezziYIsD2gF71KxqN4
rpHgbgpDLFoylo4PJloWmyotSSc2WtMXHKKGj3jRm2v6yg22ppYtqhZUMNH3xjTdtXQLkIzOCrsX
xoUA7G2KtqP0fHBX9Zu/BBeGoJYsrGPURGCO0H72jte4ln7qOZZ5FymwDZDyJEaYX/KqAOujba2A
WGA2as80gdIZUlJBryrvh4OHXqcC1lkjslAevAr/gJ3JBu84IBF3iD29CBhcyh2OCLqFmTKSwK6g
2TeJ5xicZcuSFLOUBO+ty/9CS14eW8l0dWJukmNwkvS1dx1Kb+0VhbJR7FqMMJzgj+9sl0u9m6RD
KTuCOVpT5Ac3RkZiPb8rTYyGddYypHSftiWO4EI/DFAwc1nvBZ4t8h7cKzBI1CGODqNn/oIyAUzS
Uktez7/5q4xHziyVKt0tljjv1Rg3xYSQ6oOvy/lQtZ2jHxZ3tSnsI4WKT9m+EGCGUkV9C6KZ1Wio
+8/dAl2CpQUe5hxLnfGpV+WP6fi45bDgWNz4aHkvLpUWw7m+euy8mjMEpEKZ8TOaOWbA7kH8HjuM
z5jjrpB4ZyuclhCmgug4kgF+cOdneD+K+zjKWshF5S5qf9XriWrlp54U+kLSIksZRvY8lNt+gh2W
G5PIW9k7GK35YrnbvRpCQ3n+z1Rae1f+Y+5EyB++i79vHULtLNXX41DI627dQBJcWnJBubPPbyiT
dAGtu2AHej15MstBzyLiCOA/Nl743vShqYQGJIF7Qse0INVvu/MXOdQkiCc2gngekvrLf4aA49J9
7EuRXzeLLRLXJEoBWNPYp22slnHy/VcTaPRezwJLEABwuEaIscqBPCg8d3X3qRjnu1ol9ZohQ6VX
+fG2KTv5VtdD19XNE/HJxIz2DMc3BgRe7yA2aSwQaaj9K4vZ0MSRGaL5nGX16h/q0LSkqkhsGVip
wLbkYpJfVRb6IyYmh27bmEekLPkZ5jlCWQQcQhG/kE8h3nVYLVpTEP9DcLCHN7mRv79XXKVjclg/
Oy5zFRKClx7CLcKYVy06nEFhbBu4erlhUcpLBek+Fhh4hHLyPkVApw33I2qXvwuMqqD+dRVrdSrn
Xu200i6KJCQetwKBZWySiGoSNkIn3UMW6+Eqs2pisEJP4LeQjtlNzx9Vbqj5E7GU0zW0re2s9kiY
tDQhINxPM6m/47t+f1ECTGOA4dgVZCAbe61PcrhC3WP3cC0e7Lc45Q6AmJxzhzuDqxpmOOVdQrmw
D04WpBGreOLiQ+9k5QbUXSSdd9yz1DP0pWwcoGREaDUePqMFqjuL3lGyEycMYG/LcQ3WUS3xkYx3
2GyyZ0hmDY9tEDMtQx0g2zUFP682a+X/lCAQKWIWMZradvbzF6YZet1o85dy4kk8XV8fNz0vr9qk
LR4TieFz3lVR+q1zb/7QrlGHEUZeZfa2loSXc96YNPU3jRM6154IIN+qbwBkBiAd8DlLV0RfE7Hp
qP+v9ApI+vDrkR0BWewa+KqtKEISY3xlBov0dN9coO4/BOnlOGmx1UV6frshSFTjX/Za6wnVSOWC
fxOHjf3tgFREJmIMw3ZjtLF1BRYGkJxD0+KB+zGWRUI3RG9/hfWbChh4H/6aJOsZ/kmY0eMdjSs+
KUn/WqdVaQp+GF2UhWwbDYmb7jhQfRkTVlIwyKoKkD2UUkP5TfSUgAaj608CXDdgOVvo7Fr5JJUa
Pza0sp5OxFi0jsBhPqNAw8EAU/sEGWr98RLYM3rEcWyuKrpWIMe+s32nlZ5zntyoWGjZz3H1P6b6
0NrrRhqbpuCTwg1ZJiEG0N4YxPU8VtonLsAWzHHICJGK/+m9Svz4Ric08Q1Ggh8oq5W2rEYD2GpG
8apvwED9QkUh6PGLoADRKZ1ULQZz+FeW6S3p12wCoKjm82F/L0XK/BaMyvKlT2OHUbdaZ7g0VKSa
eUkwoYA+7UPcfebEDWHHh03PSpcPUZgvnV1P/UQkKjL91appSrNrNzCPxYyKB2+xhmxHQizCfqAb
0F45PiJThrhttz8evTzh3wKyalM+bFBnLbDtFG+Xd/iGhV5IMMi2+ZRLfqzUPhfaS6tIo9gxfG6l
odGwDTCUE/AyPxLchrjztRNlreFuyIvckqRrcZy0EFXwmgVscerneD3JMPhFCQ9iV4hwb51LTsJU
hYruvWHXNGPZ77rSyjlqSLiHcfAjJI+dY6y3RjlBwaxPLaG6UXFWIbhMNBiWy06srrfoL0OoS8DT
YZihYrb9aRx0Pno7WqUHWHN9J3rRBSS+kj0VKWjB+v5BwehR2kPOZh/xyfEAdCSX+SjtdId4hYcg
aWMpjVqL3Cd7KuRN+wBnVW/9EDjAVSqZy6JG72uXjXljp+ane3pJ/+2TmXMOTaTRAZF67P8bvFti
EdobHk0wi0k9J7EaLVhrVxxnt+kyLbkjc5pJ4rhYZPEHIZt2YSV6SL6BdiRI8s3pQsOnlWfHJ/Gq
Nym6LBPXg3FlaUg+YEQi8bRUO6gLA9Yjm1C+ZtOuZrK09h1v1ruSeueSWgleWuiDVt+uGgK9/jhO
AnX+j/Pa+2IqC4wrNSMuv8GO78SPG5YIL+7Tjn63G0M+6nxNS5Te1HG93atbQKXs4Tr3xfUP5Rhm
R09/2aDjXf4OIydlGxL0HP3z/W6Wjge/3J12/j2rPe894WIzOytaRHe4X4T/sTxrTZwzJGebrquC
3oBoEn0aM8L9gU2YyQvgK6lMwlu8YSg18QcXkg7OAe0kIbZXImDSaF0GSvQs47uCtbYji8v+gCtK
4y1NYp25tLmUmgUW20CGORZqAn3j/vUF66g/JY995Byk8HrTrVm2QnvrUchgfQmv60oraNbup/A9
CSL832a4gr06GjBzO92jLbRbs/u/W8uwK8b5uJm9dovhxiBUCalWem10j/SLABlG2czRSX2Gw7Bm
6vYHGPeDqLQY4d4pH6RZw6UwVPJUphwwYIpxroOFEV/3QrURM0vG1BXTyu7iT10pUTgQpOLNK90t
woqkyhUYuJ51iXSuPPnDSm2ckRiS8CeWTOmtPY/9LRdKa2MU8kC4D78yCeP+Jv3XpEMe9sL1lksa
+pFgXuCFvurmfPvfDZNyFVWmNIT/Q4zq8lXPpTu0lJHAnu9n4kMOPnCAUxHt+uhew6jsZc1XyviS
eN+U/szunDYhtnXStA9tvs0UywOc8aTeypPlv/oqDccq6XWu+EpkzZtzrdNK2ZxmWWbMTQOw+Tkl
eDaryW3oOXsH0UM2GDRM7Ia8WAGYmqmX4LMUhLMMoEi+22uEPqfmQkZIOvu8Hntj+Dw9zN/rbCsJ
yMiMX7DHEiaI4giX5uDIE0d05tSJOzl0qmowR5LguIDwl0/gVjqj1Yb9GshbpLUt9JLy3mdTE4O8
CHD83lQVt9l6yyIw8vVSy9fbg38o6KO3k3jhbhhf0pZMKdm4jL28Z2sqJZAfAq7bH4vZXiuYBcHx
6xVI86kGAUoQvoQJ+ZIVnac8ohzGuC3/D7XREVSifgdGMHx8xBQeSIOn40Ca5jAshCmVugOhNoQY
EkOWBptW3uyOmqcLkXEcZD+9EFCEIGxCnWWixbp9aIU7+Z6EAakXnVOEPsgqdIKLLB5VPra6F7sH
awwgYnm2vTMiwP2R+y08Qz9slsV7CGy279RqfbkQ5fxfaNQ3nT+KYWWMoTHf9jf69Pe1N5wjlCsQ
yRPOMWFk8RQcaZSnaSUq37dhWh3QUNqDYXzDcGMYFEtoZHMwa8LDgguTXXaOtZ79izHtgctoNM1e
kopjCjV8RcAcEJhfq5GAuw79qTFGvviPXXKjuMONrGzS+irwUwfgwHAIUUCFJqptjyWD5iqmdiHx
yGt8n0QOd5zW/gUs11zSdj0lWf9mZdb3KnuAbXBVVDIYKzLyOtVRuCKyDvixcKui5gxQShtMEmaY
sPM2bV+Uk2oPNJnSQvJ6mUV0Ol71qZVWg+dfP7c/V3YJjtnHQlEeuVltN73XRGq/Vu5Dls9DMvaz
YSFWyIaTHAZp3TazHzF9yjgGmu5NWJMvG7VaewU22HtkFY/oFWs4Swsefe5L4G9BPOGmqan3zoGK
lqbf6D9e5EzAqVJKnikFqmiQ6r+IjIjWfOVDwu3YPxahQfG2nRJTcFsSSVMK/B8W/Ugo+odpi6Fq
HuDccL5tgToTHPxlW9KwJ+eyuJep95doJl41m+PNAdErsE7aQXlmsvytAxbBOSHl2FRyFvOChaag
LI3/CT75LkrMEtKNdB9zr5zfDnTKScV+1Wj3ZzUdtUg+RYeMCVbFuCsej6G66nP+sjT9Xb7nJylw
ED9XctYJCh65SrWG6vc+F1KYI6aPlaE1zNjVsqghGdVyahX3F5Q817JTT7I255E0xRlWrJx/F8eD
wsuPfIgicBFoBGXnd5azKj/pOnu8vRGlcKpj5ANwOEyEvd6686oQCGgK9MSct3eRDBo8IdAn6ZZv
f4Dgcq9ERgdLtuPryaA9Rb1NOL6Gp8AwaPrRjr+9OnaD+Hj1xgn3yeeaqmzAr9RD0bQ5MvjBPo8J
rtvl7mqBMZMArzAE76XBJpeQrZ5dQFTN3pMtYd4Ymti0atJ6Cp0RaCj2W8rhI4yerQVkPOJqbbIe
wwflL41/6LfbQkyGYHUluj4aDAaRDof9z84zyOQfZ7WBxu0GgKDfipGHWHHp/MRG9tPCvC+e7rin
ulCbKFtZMfymiT6bMNPGuxZsLMKvh77g6ss6uijgUiTr4LB7KmNZ67M4TBqe4rpOy5D02bob8tBk
BULRK+ARWF/+LWX5XaL7m3gTylYMIGvgkb2fqr8g9m/lhMm0oqSwW7MbJtjP6GesCIvYiUkb/N3W
Rs6Lp27kOnfHRcgcpZKPMJCaKXl0QfQn1n66IlTmiuw5pXLQ/7OoBoT3i1xEUo717PInD265ZNQ6
x2Bi4xGhttnkl3m3h0UI+vOwmZNOOPnHfuG091zXrtvG4b0lQQxBhcP8S0QqXH+9/wo6Db4KAmid
BY8EYPukpU7DbLCLNfkqbcK9KWzVkwTo1L4i7BfiQg20MzfGsGSB8VdNeW6mVItDWj5XQ9akMRxv
CR8EJ+Jp18epSHCPxfwtfa4i5pEYU/sUcrslC4kD+K8aK3gJQ3cM3MdsM4rREzbU0jz/KimCLRel
kGMsPMFw5V20cSUXeonizKZRIZ1mDmD9sZ6sLo/BpQulTFo7RkTVPDMlbTmbZfk1pNatbDI7E1fw
rDbMIasGFoYdQD7hpYOWwRJOjzDl2pNUiS2gfYYyGPB8QN8KEEJ6jSu4bwMzfn5pdUCpXMizT8X/
NZQF49qJuoqZudtFuY/hdPiLPKBvUFJ4fdWy2zYHsr+1L194ZIicWk0XYkDSrEwK+JnTOJSo2CEX
JcGEiLU1jvI0B5aWhMHanI99yhGygaOHcPPhlr86eX4UUztVNYIPN88ZnqSdfxGM4gMwU49Wndud
GJSJczBsCJ5ZI2HFop0KrOniHK3KduAI3YaW8M7zqT6O6Pj5SPpHpPhR/aC2r+zQQjxbKOnSDEow
HNAma1k6fejbScKjcV3G7O0jlKsSx9Vdmf9Fp/KgbB6yz2Afk2ZTv+nxKdkT9UsqOVkGIAXUeRzQ
3cxx/fpPy8OkRCRavzLeVzeGwue0BV+jnOJltXKJcH3FwaO9AESYbIgTwgNwXj/UrYVlWuJHcVXp
8qv0CNsU/ZMDWLExDo0qSJ5MXps9OI/iNiVy0xBGnvPMUCBUHXph1Wl9Ol9UzBXa/90NKC+o6pNP
HaAUT54p0sk/75rZgr094XGxjs3IsQyi9tLUwl59n3y5VHjxudkyhpDfZLSP6q3a6JbgXVOE3oFn
zsuKNBVUODzpA+RnsthAb5RSqRU5mJMfNFinADrG9Ijc+M7xHb/CpPg0mrrMaqsNqwoKZldyOqbt
v0M6UKYVmiIy+Z5qIDIwy6MnC1ypmTF7YCYL1wVNvkR/9bzJkv0TmBV7mhVsWff5imlFWNBUKGXh
INqQiE09BmymI6NYQn/uJ6FMxIj0PiVDh+MOGNE5ReggwDdlKDoyOKRbBYuyjA5xclCPbwZnAB0l
01RwfSQfAoXHEudZ6Vq0veox4WQ2GMUbher+5VqE2ZPVhx51IHsRpDhkB2XUu80qYabz4fjW8uQs
37XliK0oXWR4Vai0pi+2NoZqaourCH7xzkNbeUtM6VLNWPOVKn6vqB/KldePfJAHQEuSd9Koh/L2
M3U6KJbXro4+QimcGtxG66dc4NfqZ7iud8OKIHPIVN3wirYjZt+NZL5Kqrk9NTfJ+Ok+zLFWR9oO
bV5e6dYK4ixpqqGis14kfySuEqntsj/5ePtQXz2OgD/+NGBlY8JO4SPsPlQyVN2XCqiPoipXL5hB
ln5NbFyXq1Jpr/2OFsXlPXg+cD232lzDzbiEWCKWxzJQLNr92QWl5cg5Flc1xIrotRp/RU/PEuce
Lhoh5H1lnYtp+4MLWVu8MFW51g9sbjVYNimC7riEnMpw6kIImn4TLstFRbp+Y6gu+dhbSrtFFZn9
AlzHIqFjcJI7oiNBX0s7hyEm8+Dd13oSjUDFPx8vzRJLhvfmrOZwU99jc2RmflZgw6+H/TigMFns
I57CxIXS8avjkJBMjcoEgfn2GTEFXSvVAOTgD9hGrk9uL188KoHYCizBKFMQkJR9gO4uGtlMbI9x
7T3lVHKN7vcZnNiJavAO21oBcuhY+AWNrOjofA6SPkWh8q3y/ql1DXjPhmyjzYjtF+jBc6kxrlKX
wEKzBZCB4dUKOl41kQvtNzJFYj22SsqW7aEpJ+xNYJyM8mUMemy4nHWE3RCBHYxYnXnORmQwkILy
s8wTkepxj8BGyiTzY2piRZKN0c0iNz87DYuTpsbQ/tdkJj3z9fbBZo/QzZwiNNIiBy/Zi/m2d6n0
xbdUzAa5oI840XnSecuUueCOzTnCsNzr+E0b6JbF1f1zTZBQHnr10ZxfbXEfHICaQqmYKonQww/W
Cw9jnZwCJTjK5GmlmhNNdtYE2FdFhZv+0KW5Wo5K7BHIM7azIeWBL/Inbi5KxxQWxO8I3Fq8KDSX
o6aCiEIxL45AqlCcW3QbKuoOpjZFfO4ehsFNhDouNvZaVyIRydxYOp8bBou0JDuo+dTR9uc5dJMp
SQ7ZXY7F+U0x/dVBuGYzTLB8M6k0LJCt3psk69K5IdO9PYpMwI3KzZvCRUZRpsifnMuwLt47//r+
2vypVqAGrXKvgkLe0NSJYTGG/IZD5EiHH1wgFnNhi8N/CynljMwdKbD4D9jOLAnerVaKrFuMTPaa
lOzI9VYIo/t+ZKIGBgntgmvyjv1xWJibddDOeNWqFQHSJXuGN0RYF8VomO1NRXHwbtzAXMk7Ny5W
H7mmH+Ful0KiPg81oyinATtS2uyTGosLnzNESZ8zT78M02VCzaMiztSHm/F5NYO5H25Pw2D6oRJ1
gSAGmclMl73fMMddjcsPQOusvEvNztjRSXKR7YDiu+LyOLHJedcPgeed7xWebXAfpD66s4icYVPm
gmEm0UEpn9qVY2Eo11sWbWCSHhjNiSoZ78y7EEeSU3e+BIcyZtHpQhKT20yCrO9fybNMU+J7GKzz
VMCKbNczdFMubkHN8GjK3dj893VrgO8SRcPkKe9D5ADyGQB9ldZeoojA/0I9Xipd7Rj3TXw0luMJ
vGwd1jN72cmvJSobvV+erv+0xvkrTHMWDT5NG+D2NBKuJNbTDaTLfVEtqtrEbOvj8df4qFE2wAf/
wGB5cXVCMdJkSQ4GT24D1S1p1CNFWV0EuE/+XD2FQ4sWkt6y3caR+OPQzLPcEBLiPRtyawpPPKcJ
0yFhHWXGavxKywqQNp8pcOgnQK0+WH6bwCuBgrijlYbhvNUutstKHl7wbx5QqzNXfWOrfFMo5ey+
AoABDRBBBiKKQTNU3+JjCK8PeJ3MUi6lBjoGSn8YDye7EpNUnABwPdPBTZWl5+GWKyQ/nrMDyVMD
8hzLzkUhR5rcAgBrOYMJuQJw9CfN+4EvcS92QObez8Wt0UNq9g90Hd8FCpcZ0WKynWm4MKsjyxlm
m1oXuSadDaOvROurQAPHaKq52bVCnBNpiPKx5U25T1amqM3xxPtoD2yrf7apA42BB+oho/b0yQz6
MKxqJMeer5Udbfyn1mBpzRCOvh30uLzhax9tp6IRN3UcnmVPsBpRjZ7rf8WxaOY5fvGmK6SfdTmO
dxY7A6axyn8LMD3fpfDSKMuECDTkbfz8L3w5sQ/sW/7SYAJ2S4zaXJbQyxsTdh5i35NtsoWT+Jpr
xB4iSdz7kmeWsjGEXcaK7Ikyb+AbO5iuJBBB4fUaMe19I+++i9/8+UC5fcutEpr1vG1KpizCx0PX
FJ/8tCcddusBi1A9KzzZsZyqum7wLYZnsb/D7ZkMmVSKW6r35ws2QdHyfNmRpHy0Bv0+D5yFeoYI
2YwhpnzgShj+GUUkSFyVbXXHjgetEUA6yeiaQcRBHDtIoNRVqTe69bQyuLzD2U8yIA7wbVds1PQy
IbOwtSBDxhwixVvK8LkzuQOw3zb9JhRAu4SjJbLgcNqRZG4SX2BOw76FG0QAKZ1PSL9H2R7QLGog
V84XUaTDOtHf2Bkn1McOYxooHFFtcOgxbYFWSmLxTGXq5MYjVOpVoa8ef/Z5XDaTkajARJPpLZDV
1PN/MBu+AxR08prexX2QGezGF+Zw5cckB+u5YBxFJtbpxV5FvMxeIPKsPb/g0mChfNPMHeAR0ZqG
2F2boCs/YGpazvJq1ObUpauVc2uBcvqPoWaZIpiIdbudNxLrtKBLnmtPMFCiiwiz6yMIbljsJ+cd
fYJi+cgMvDlBZxjgZnPGbTMp4oWy4KXWkAAXYJFOSD/Wp6W1W9H7cGTnv+cuiTPDGhWlMP9Hjgbw
AAZ1EY4MGRGsuTd9z6e6mtGPRk/3PIIQKEb85z03WrIFATKpNzybtjQV1zLxn1PeKiMSVAjRh/Ig
AB2IKYWtg1E+94cCmCt8qhpLvBxdUgV/YRsb6mIRPw0kAZWJppBadA11r667GylE7AgX53rqNyHS
BM0qRNAUnTr11oe6wuD4jgX3MewpDtUQ0Eg1vHhL9s7UBA5FKIR9peD9e+WGSY7TA+wMtSucLFga
fevPXXB+5Hq+ey1P3zlaji1IqLBIrbpqcXrAZFPP4Z9nGWztf3CKeE0DGwTHy1C3iYFfT4ya+7B6
Qrv4Dxt3DfxQ4EtNcMxpXFOmZ/OzwYH3mod9mF35qSpR4NBNBftqe43PNPk9Bg0BiHNLSivMISdW
YanELT27DFFezE9UTxqj0u9KoWJGZIIK+gev9qYfeRezBwBT/rovIY8utt3+ObiK3ubt338e0Ck3
+vq0eu+PV5aZbLGRf6yWpdwTlMrJkBLMWhpfAn+AKyjDfkYLIJpaI6kiYG/nmM0um4vuCpDgnnsK
URukLfTflCtyWgIJ2fAkmYFjQ0Xg79ScUF3ttQENoC3Qqm5DQRG0LHhB10FQXGEBXv2Hdp/5lJts
NMrTCsyJumO2UW7VTbOt41HGgfPowxNmH/acf9UGn2A3KD5bRbXLKAu6wLZ3R8PLmUCkzeDBMfTC
6vJtPPiEB5Rt3UyVAGSfTahSvBCVgQKCVi3vkmxjWEYdUgvLNMa1ZhH/y746SC2MC8cyfjPMw4vd
HyEal4NMxoJ3wtiB+qLPKOTVR5GI0aIYN3TDkvF2mJn+gmYpedYELGke5xbJms9quvlgoeKhuQZ2
LXzRYOg1jvy13yizUpOsit/Bg1HYN2R1Wo+diHXiCo5FxmxBiednLW5f8pqWQHb3r/bwMNMjCj46
zgV6cb3Z+VznilYxsSBA56QnC8JFOogK0s6SGbksBYLNOKLnDnwgc/fbe3h5KJhpOOaD5Vw9LjFU
KIzj7FsRdtD98kxm/aS9LXuZCR0rYut7inQdXDuNbDQPBWM9Ij84WhXuyFQ+FBZ7EDvZFNLjkzzF
u7lDJzun9UWyOZZsfmLK3P3lay0w2jZEAcpWWSpfFe4rJ1o5XLOUyKEAeL8uIO+/5rHrG2wRGaRK
Mwga/O1Zl+qDikRBmgq1wuUeedbOO8sokzPqumxNATZ1oE7CNqyRfONY0+1ZrhRMPjktsIy1biPj
mh5yQPyXXyiH1RoUetsjocPgPyVdHsFdeO+M7GpE6fsPxD6uu5qN+NrgTmwe6MMMU81uss8sE13E
NAUk8p/PqjXXSvvhjBB5UZXqr+Tu091ljWneCDfB415BIUNbhugD7QwesWR6h7onzJfoy+LarUkR
lGYXSsw1eESWty+iKyMRCjDP/KTLMQn9FN75xJy273cqlbJeYt/Z11uNaVcjOV+SMNwhhcJKROc+
jZ5bGMztp9bVnR8CEvcvh6GVhB72ua6g60PnWDsNeWi1JTLyQ8vm1OwFZKNGMt9gmQj5Otnk2SAo
enn19jeeIJVZ1/v0kiLCIkYE83wwRoVKzi7RksMed6PkvFnM6SRfFM+4KqUzEowKOufEcA4KK5wj
HyyNDAdqX7mHTVRhFMzB0pn7VP6hyVyXCPgcU5yCSHWad53FrNXD2AAoWEG8IYLqxqg/Vjj8py5q
s2KnAmxUEA97C5rWKE2CNgv30CnZDgSrLtjLLN1GASr2clmSnlIedbypXjlBtEr55EEIt09GQV40
YLYQdxu5zv0jjxitZ8Xlhn8ngvKHgtXZsWufOIHb6yYCBvP4GlqEthXgV1lNTfNhd37Qq/2eISX5
urZ8xwl4usbP6dwTz9ofLdpNLNqp4RWVVec89WcsE3fWumgDmQiXQtKu183wKt59eNz1d+hkZQpp
kwuzUjr1sNiZ2YS5/AQrpaYxpGpl+WlpqKr7nnl/A9eInKcS7/C1uz53Jn/5IxL3uHJ+OnBNIB3T
NQTLPCMVd+mpFCG6/9N6FRQx8esedIXzWS7kFJBKRfqjdrunAk+kD5f28+ytnl+w+zy2R25HR/lK
0k3DSF3G1iWsVtIWBYRjwU2ck29vgro5Bou9GmgIzLDKlpKbIR0s/EzwYYOQV9uL0OcUaJwzJ0VJ
1L80qH8IqClmM7lpKmMu1sONKbnyxDwFsWhz398KV5gHt5cwLfuFpOEKtS+cyggsdfO6SrKc8lF+
NyFRfiooOH1sSLe7217TeXNEyNPmNjDC62tnLr+6tsNDsc3KVG2Pzvz1Tz52MHIIxnlBcCy4VdME
hNW92JJ0924NIbjVf0vseaKm8srcre3zLeRXCKukUKSqG5oFdpS5J9gZcki43XtJFOAdQrWf7KO7
VYFRPBILNj0dARb7angwHbUPU0SeL7pEe5Ii1/tNvNmF0i29ceoh2cQaDYOrppjaAsIUInDgWTE5
tN6ZtjLkCnWNx89AXpO7Bl+rc3GBC6HMRwCfxTtcjbT8Vfh1p3aWgNIvgr659xhdTbQC7MDGHoOQ
ChcP5Q0lhQLgNXQ9n9V02SXeasv0o8SlvdvsZfUbnH0ZJ8TuffQkmtd6TJut5Lf6uDJB/+/6p9rt
eLsqLmY7KVxJRuXU6Hvfe+JO5AJTtSCBLqaM43jZuiN70Szzk95tNRZK0D59wzpJ4lDJaf71U/q4
4j8kII2VzvPIdh4ZLL5IqOsgHpjp9FyL7ywaUEVqgyFp16XvSvziVB7j2BOdiKwl1MtHupLkSrDa
g+DEUGJWaf/qLCjOtbGZQXtfJypwnhMjIges1RgtFsh76AIumLr+8qGDizSGLW5jAj9tIvaeTzKf
jpKUTf7CM6VORvDPncCsAEPNYPS8qtl3XXa43PrOYnYIJ6xw38DHUfYkrcfU3lMNKT9eEhILoTa4
V5QWq6h59bEgAsqT0NGxlyECiRypXBV9E2UIWk//iw/UrGwUjCiF4BXJ3V2MDXTyl6cF2zNrsj+y
IW8+NJAUirzlSUlx/R/akFzK21GTu9b5AOUPm6n31b3mgSlaI5BTTHT+E7xYEUcOUFj8jwwroOb7
8fqIXcstLdyax1oO6o6wy9LP/6n672cfQvd4Uph7zM5KozI3iFZqcd9xefDFS3jFF3qQ5PirP0T2
TxKGCQsB4puI6WQvbve6mtrOU8Wu8sSnDOTJ2mfesTAzucCjhGr8ceFTdcGy9bdT64fTuKiuKhI7
UqXOCk4QtU34EBKeBwpsCaPENmWbpyL9ulRjo1uIg7LY0+JaZzPUxnb4ig9Sh2EZZRNFLk1pZDpU
z6dX31B3VgfPsJrCOMzWevXo+rxLeR5jDCcI5fqiRuBztMea1czGKfnYk25Di82y454CUra0Prhy
qJC7TEkp1Ozg0nuygI5mIw4+YZoFS1pIxq6TBfmJ2FTjpmi1CAu/EruzJOL7VyUch2e3Kvu7RXoF
6UnnDiz89TjGddbXn+/X1aYt7HsL7+180sI6Aq9mbP6lV3tCBwis+42ObHtkFf5MMIH4g+2Koi0w
tOO9blt060kgUJNCaP5Ne3w+3GVt2cGvygOH1/nrgszmBE150TiC+W9YtG/tOcILWWCLp/JTlYr2
0MH42At2fjyE4bv6zu06J9FLWq9WcpLSUEUxMjuKaDmAqQJx7/+pyiz1MWTbxnuwQm5IIzu9mvyu
FmdTqB6iNSY7D427+CCXhw1Hfk+YH37loPu6HBXngSqeXHiUO+hHvHdNpaykSzO+m0RENij1MhMe
0KNjqgpg2c3n5d2xyIfJiUsA88JfT3RmcSkCSrKJhQRbwFHROMm/BlcqB5+LC8k1CPOm3r/uQB7K
Pi9YmAGmJGX0B0Rlq83jW2SE8wt93Liwb2Byj1U5u2M+FtRxu7XmVbEXFZGdjRwjR9U4sWW8GU26
w7EoEut4JkdUMjLNlHEXU0KSdd88nz6aQFkahQSPm3BO1dL/nVGhb+ZvSgf1ZM77JdfDLMC6cP2i
DWQoClT5JAJNgj0PMhD5EzTdWQ494H9JvIz+JtO6W4Beht3373ndFBnHGBKAkRbWnouBzpTPPeuJ
XpWiwCz68OehBaqofcfrbWBW4TUEPTenu+kl2S4Sgks6DGVlPY5QvFuUapX5uy8RRuMAptIlReCt
0nfa9ZCstDZeEmAiumulJ1v5yo5jIkpL8UWlkAncu5Oe7sQMvsAZR0nnQ4MrZS7vHW3qaGPVXpoK
bhEn7eCxNO0UIb4v6V7cPJtCZIYQVtzr7QgiMSd+phP2Xj2m8SMM6zw1KBTNKQ7PxbMsYbhAAMoc
O6Y1cG/Ou35F8YvV11b/IXel4wfr8ef5CB0cGz5xXId0lKmG4y/vdwxd/pu88IOg07dg+E2OJzcD
v7eE8xPks8ajOIiKZRLxIvFNm8HWQLUuWPqNjg2oUqx8jczMqKXIO3kjeHhKtLuXABr8L9gpgnpr
334nFM3tspdugVq5O8miaOWulgnD8b/qqIJVnqyZOrILFFylrYiyKtwEXfsLnfsvKFDKs6D5tRj9
m/I7RNdJNKriz6RvaRuh9cqICkxXi6FllGXB9mrf1SxJiwg9izqdz6MPQmakNol14ncpHKl0+qSw
1eMNgkrMQIDZ5fue/jRS+iDJfae1tTDKeeAQlus/b4R3UNseNVLH3J3LgR/no3PSt7niuElCzrWz
lLZjW7kjSxMRKWr4H/mITRYqRO8YjiQXTMcXn2kerfmY8p6zysf98Os/pbUXKqk36fNgZjm+MSJa
XL7PdnoepjIyw8Hgx5k0awn1fLxZrKJTo3slYa9l085ZC4doiH5ktwgDSYygEILtthoJ+2m8M0Zi
vOAiYmMOhSCcon0+Ql434PHMbCEy5jV4hOARHjEaAdL0siIDRID77iulIJVc1RASLcmjTTSijjrF
uy+hmkGJoiNvQAhKUapsJ5rFB/y74oNAvWFE4c4kT0Bs+Cl/6wcCmRPcqWjhrmhyYpcEr6fg03d+
7pBkQEi0qQn/nwY810jRrOrLZX6Dl7DLDcbwH9QrMYkcIhwtO+IN2R2F0DByQu1fkOxg5wM7Nto+
bCRaf5kHian7DTeDlXb+CPR9Y9Y/c7ZoZeQsAxqBg13xWNU1F6BjFABABwSUwyIs5M4Xlr8M3Yk+
kRDd71g2JJHQcscIG8sFJhCdwBhU5Mr+JvFJ3iEdV8i4LQiaSdLkXFMnas+HU1EHhkpMVejo9Rzb
H0H5lUlLHXuV67QNKNEGHPfAiYmi4gKZmN6tHe8dFD6rn0Rp2K8MII1V/k/M9GnsnGr1S4hBq9Ky
HomoR9b8nZn/FwmM+M+WPXigsopIf9P88ngzRizsXXve90rH6WUJxF6m4xusOcp79R6+sXwOeWMb
LS9Rw0O9VT1rci/sC3/q74X3xb+00wk8bM3DUH18+Yu4rFG8qK9ULV2bu8pqiLzXh9bYveSmAQig
K1WGTWdxLSDb9M1ttytHRwmF3U+84aVVJ3ELuxcFmgP0gbk4bCnJx6AU7UbZRrSVxlyZxrODkdZC
vw48V7QWA0I2Cg+IevqbCo2E2P1SKyKxZUUA7cQYcW10dggTkZSKDICgsDzQ7wRGWieQFjxPWhEK
hvYwL93b/g3BbFIXPNs9BuIOy93O+OhD7ul21woaSiFxmbp0jnh/g/7zoK6x5vWfNL1h/OYghi3j
gvUd8+KfwyJ8S419Vis2TRMHK6GDqg/60+K68UJwQz6jz4AjeWXEsZv629YyoSvJE4y/b0fg8O2V
gJzcq3K/y0RsKKVH59r1cK5XmnRfdLbfIKe9byK/vwq1L0cXtnBwK5RHpf3HTzvUvmq4tbwOI68Z
gHkkZ76WV1kj++YpNs3SeYpuhmMCgFkuBXx/KIUPOLQrIyDkHDwFL0KL2Jo+t+DFjSZfuOHtTewh
QEc7HB5jkZFGkV3GvplnnaFGzMwMm7nmLerwrKWthTFgayXlWKcvLmLp7aETZpLXzr8JO1Xf8OPC
o2FZMSBB13p7JLHymno0nRH3y6fSD+7sYsNyfTiDydMkTND0Ti1JjpJYIJdYr9Ny8E7Bn9+Ap3te
BBqxPkRtCzMXP7tdoEmwbDX0SxwWMBHZOvLdS5PQcKxHEilVp2OxBH9d8XVxLwg6pPdqpjzoqBjx
cHcH6cuuC85Z0kG4QW/mOeXyJyOeoG4ae7zyfXBhTIL3KLbNEbn/2alVvJvetNCCKzLzpi2+1jap
se8m9pVwL7r98lm0/Sbh7zp4VEq3EZchFT2G54uW29OJFwSuf0he+sroVcDGqkFg5tEOiYZgfnh5
luR8uqOgUb6C395fUK4GgPBYW1g+Jd6NHJLytxrCU4yFTX+BDwT2Gr/KX0KVeFFv3MvG/sVfkWsc
BA9kpToOoF4p2DnMm8WRXrhOFL7eCPGjllZkamkYCTm4v3zk47TpdZk2Et2tqc2slgER1FzAtxeU
1TV7M8uF/tD9N9GZJIQsHF7asXM02lTFfuOVucCB/F4TIZlnziaBhfR/NiJtDXXOz3EeL9Qe88G7
TZE9zFiyALh8cuos00XJ2nm/6ZUdTkRr2Qpm2CZ0j/VUKND2mRq/AJMKzSwAVbxzpmoHLp19SaE2
UB3B0oPA8Ks8PYu0FGYKPjvQxccn7FIqSUXF1G/ep7+2DWbbPI9X1CC0bMW8bAwujx1MB/3qvapT
vX5NlG1lJ6cESrv1xGNtA4b/4Oafn9gTkzVn9WC5gaU1noOD/PfM1loWuxzOyW5HJxSVF6mBRQgV
0mfcanS6mhDVlNIge2iFgF7f+ApYDrTmJehf4XPoolxzxq7PTxiXrbvb/R5Sfu8K4bl2o5zBSgmR
6GOJ35P7ESzmUi5m9btoUHTi+aw3R3xcyP2Oa2SZygRA5DNdiD91uaT/qXn33kpQUe76JyVghMck
3RVVTk/HaF9ojqnHnuRYNCi8L05iaj1CQND07Kb+1tmhLYuRL2LFajZpFrlZbvcd7cx+R4yOZPFV
NTOMGOElc5LklESjHn77BlvoEun8MWkY5N+YDINHyElfAECDfHIbi2eI+usJhx2ZjnDg7I135LDB
Gqxs26s6pADL40NSN+0gluW26UIYEhf1Wjrq1SsPJP++HJLiB3ny6SXwjfeghK1dWIY314VeLLiI
bEyDBFqd2QN55oF5DU/m1imfwCiHYoTumI5AptgXJm6E5rKewkjo8kVc7OsT00CouHRtkSs2rWJA
kJUdA8YeVUguaIkPjThHzyOK4WkUqj3lIrZsFxst9NXFYrbDhhgrM+lVjbsaSaXn1LGfbpuJ8+ps
NeGcx8G4A+q+5c/7f5/DBoUROXbQGYtJflKhSDdtsGv4fc+9Wy0PW8qMUp6IxpY1Zse4viP/htoj
GLWrkg1lsSu3dlnpd6LLtg2XDk5zPOF+4o+01ByuV2FDKc39uKcSqMVnI8I2z00N5lQiobUmoiA+
3omd8XcHVgVv91AgYbMLx1eSaRfrHbkgGTfs6I+gWLSIxQUxN1TTD9s2xltvLOZKf7FG6bB3bBSE
tdCGD4mH4aCDmS/Fmt4+O7XnyZtiZz1ylz7LYCDQdGmXBnG2jT12X3FlarfIAamPpGjebNTCernh
ybfeCQ8R7qobsjIO2LcyMHiCxbNePeA1C0wA7gasxEm6lCyrrjAYgJKzMoaRfHJqJBnBGUuKYdZo
QpRsXABFHDgARzXOk2AHhfbArZbmNRg1JEfOo6ihW6+kEtJiYqQ3gnxeBdRAx6icxSokhkwVN6cO
JN5zQB/QXdx+qmaO0Y6qthuCK7VBytxTdn4G8AQiOlAaIdo1uTA9uvs+8k5I4+cljlzx71KmsBd5
co+m+vAc7Ksjrbb2XUulKhMPfCkdqcaUlJDBLo5LW+VppzIxvFzPXJrmidpzKaFCpcQ4VDjvKMv5
HlamiXT00yHjRc57E7dAzCc+GUGPdDVqkgxBb32fCH4mdedWTRCrfQJKzuablVW7pn2N2h3cO1VB
HfoDZkRgpbp6dj0btSjgJ0LCxbMCWyHEbi6lmZt27w952f3nzu599vv9YxMDti2tpw+JxfBSx0Nu
xtwfFInBt7baNOzX6bsuILoMUxzMCNHPFxZBobaoERBFMTekTbIciwEK8iqs5SYtP9PuD20u+/1A
Pc0rf7L8HCekWZ/riZJ6kmEZ6iWZ5oc1hKgRqIlIfUtw7HvM01qubHxRWGMUIrUomRhgXMfyDWNF
+e7ePk22IsDfwe61faqAJRdI1fhQ4ep/nB4FGbZbVGHilZzmzAZc03EWe4/Tx0FlQf4sy5dgaSSA
H2uL+rPwffISpvxcMhOTNGJSWMBNyTOx7WAGs4DtKpfcf1H1MdEbcpBF8ZxYp1ch+WHrMYSU4F4+
opI0iBpqhmccQzGuZlWC6Vm1cM6TT+IzYHMZD80cFMzrFensUxMUe7RsMgneWROucJBplpoS0Cmb
NKU/jvPlFdu670dZAjWDy/B8ezYT/FnIYrev4UHMhvubGaIUYSQJrVXUfr1tZdRa/kKvGDb/TnVW
rLOCeNJaDUaNrpsOoaCT4BluPEjTSUBx5WhPnBL35bMD7Rr21uFoA0b1KAKsQMy5YI1dkH2zhYnw
j7sofRbjtWJEy4wmFVbxgmxYCc/oZLulyMHrtq41130CkoQJTI5yXER1W9nxSkqwXRwQKHyXp7FI
uZKUGD2WQWZnT4U3WYkFvanOohjSYQTD1QoJnJI9QEKnVqTl0ru1P7P6ydv7URd/oAnH7kYgXP+o
WfCUEfPCsYCHE+npXKePN77dp2iBcAY2vIW2yur4LnuQmt82LsFX7CSfXYLyQ+ZzGIYU6dMf0Ac9
Q2rzv22hUwyTLg8HLB9HIJl3ECOBq4O2GfZck+6QfJAW0yLbWy0K2hxwStPf3Wa07tErFbs3Nqfj
3Akw69AZSR5RCPqD0UvaWnG0SdjH4W8O8Zgn5MJLCkhV1s6CwMLTmNckv6VbgmMKYRAdbcaBw0mu
ezTiXfqkxIv3Z40jXdwWn1yiJA4jMcNspYeWG5geiL8razMZ+MwURJUsnY9Kt3VONR/LGaJvxIIh
65d5vKAXHpI+VnfNHbMXauloKm/X0h83MIUL14meaS0xacNDNDb2n6XeB5BC/IeeZp3qMu+gONNa
x/2vHZLOUZvxn1FnWYNUbyynSy69RW1NrneHQFsxJ/BE0QKLygnJggXy4iVo9SIJVg2hMekHFlY+
+c+woNzQGKkYLwqlokHosYxNgRsX8qhAT9vVz9273O7vHWLOTQDqekS7eqLPFrw3AQdMQ8gOacER
ST+wtOEDrZxDFb4FBLv5406r97vCW5/KcEdNRm5FL0u3kZJJmd8S8G2mWAyEFXEeR8Ud/N9wUCEX
h8mr6gQ0EKDaU2EdOaY7soRmv1NFHhWdfCVvl2nVXNrTypW90JRbFMmW6LomH/mXSk8gXU/0rrTc
JLwkeBH88s0hIpbrkIyo7d+wd8jaAe75MIZlIyJWwN4yiFNfH8WZdEcJmfsr/Op4e5UOBu+f4Zum
rXeyvGGRaZ3UrwvUwqv4a6+aR7Xn6uaTKINqUnMIzasMwMWXWwmmMuFts1eYQpkphcq9xb5deW8Z
Ay5xcf41XLQAno0I0Tihnp7zLVKxNTBc2H43YWBdQSZgQqwsTgmg+f2pMyn9ja90ofd7qjzSvRbt
XaDgyI8UcUYo1sgRZu7FhSlwY8ZQgY7eHuzMhqYL4m2UHpQ4w6cX5q+LFPeQyZwPKufXfefmJQz3
yQr7Y9f7D0TtILty4maFE8nhEpTvVAsdId4be7vbJSy2hHKvMROnGaxzaa/hr/StVhmemua4DpTQ
8qcj2ctxE53xKEvcY9eAVW0skVP3ZcNKSrrlSaAF/B+3/ehEaXAyViZ2XMoSR+DwzcuOEYqDrAuo
AvUn+BFecO7yZkHFDpYswDdLm+4OlOHVaWpwbUt3qMd37C7hmr4RYUT/Yo9i1AqiUcZR6oVfsKgT
PdOKQj2C0HHRlq7rfO1Ot2KoThoTk9oxFcYU/+HEL94ORJX8IoK/W3ptnq1f3q6gW015os3eQ7t4
nmHL6crhe1GBDA7c7uhUoy9xxKY0wDs/e1J98MX5R+pk/m+z+djOX1WXTZTfClJfbHzF0nyvlP63
Wr2wsyn2snMijhfkCdeAprv+2nbIXu5xG48sns/YHuAN1Fh0bDqAF8Wdc3rbYLVHVn/9P6oKAkbS
0g6RlyYLZamtlD8avxtKBohOzc6FhT7QxCxr3/E292q6xUsN1E2QWK4CHN0R9XHRvVfmMzY6M1Eu
1WP4WNNPb5Pk9m4blPEOXp4mcSPpgVc96tLBRiWUvra9bvMB78viH9BjMAkgkXYT2/zV8pXcYTMa
uXb0QuZ/YEu6X6VMHdJYQnJ1Rg6kvaJauD8Ls+KYaS29WLvT3oNJwLT88KAOEK3FjbOMpDstJPje
v5LaGY21awFlxnECtE+MbiUqbh+3dzI4FQQtnPLa4X54B1uO1Kn1/vZzXQ0Pa+FnXifism7gBa0x
SWGdFizELppsfcaVPwpIP8WcRN7YJVq784Hwfua5fwkJF4L15O0uecgtsZnLxEuxw8+iwutcU3z4
BsSQP/Zb46nTev6kCDf91Pu60AGRz9qyV80gy4EzAM0t26DYeBOyfY+rlOLNY/jI+N573fXIUWJr
9eSmvcYyhhiqH5nBB1oysU9nTfS6SBlfAZR8GjUXvOI9ZbUbAlhChRAhdjtBJR7ARrtjsKGBc2b5
g1gYYUOcpo1Z00vz4FJKk/XfZfzTydpLzNIAVkKBW1dzKIHeJ0YivulqIblZfXHAuyCw+imABgj2
Z/aP1UM3aBsNax49b3CzgTxsO32XA8Uo1yUuGGEjEL9smSKqMhjTUE2ySh7KU4qLTGg+wKj4ipGJ
lO382ds76sKgv0sV/9tzGj7+p70+TL3quQiQK67+FRhE7wgCkzrDp8fWRW+MNBuFW/0164KRhi/p
hk/wRsNP+qwmH/DzzUf+UCyOlL5TbjS+YIkzw+TNKElwiV/zL59MhV4LBDuWl7wz2KmVTFv/v/1B
GNvuGIQTlIHN8cmAL5AVxcoLIGugkw288Ib1mBP/SrzLU36oX3qJPIpMYO/OkPbmjw+Cft/pI0l7
2fnbxNDvu9GvJBejQlErJ3LEQOt7NVMFsRAhOaQiJ8ayyNhKFqTdhijCq8eSXdviKRkXUJgdZXXz
OdfDL5YrAaGrtmRy6Dk13KRu4bbGMKwnIiDSSVl1OARQ0VgZmmOHGdP3IMdwjqXr3prYGIuC5UUr
8Jq/FahOfxjnQsQHZzJ0fkWvPv18g3gIkcQuK0Ap4Q6b9B3QXr7wXR1obYiH7YN+phDdVDk6fLvc
tyNzSN93y0K/eJ9bHZxd12O/fEKE+WZCg/nG/DsN7b+tfUUhku4ck2b9mfQ0cbcQgPqlnPFAEOBI
bPUGvVZbi2hIpNxbIZZ811tElUPNDWNaS1xoDPBTfuzdNm8P7yg5X1GDKwq7+Eh1SBR18iK7B57z
QJBnprAvjw69TDfRxt/DE5/fh/i1w3VForql2u5z7Ws9sHq1aY0wMf1lk4VGQOjKA8KGIkT9CPtT
MyEHbBIO8DcC9/jApBGIwWZsWI6i12Vq+p6tYqblveC4zL7IqcLBGGblFmNX5d2mHiJJANpQLTOA
hyOYLE1N03ChRuBjcXR2Vkkr/NEG86qCVY35U/TtS/efPB6gX6aMzaES5JLJ9aUJp5o+naIhQ0ka
g5KCgHYUzyAURwWLRg3LPqpf5p8M+TFsUt3dBA/tvgFcjhJiEahyHgeGwAwqCadYYpi+h95KMekO
+jc6aUDWTfsj4/ByUx5ica9lSZKPMy/hxTaXDzcXrFjHQTPZygKT+dwI8cw4cgc1eAWVVp8mduU/
oux2n641eSMQUWMWPOZPLU0w/MW7Fq8pIJ5Q0uXrHiaPGHEmQCWLc4JnfP3sPhPFEJc72Ad4lAB1
MoSHbXVhd0lPmjseuMitp5TgGfgQlvNp5vED5tGGEeIj7E0a0gyzbEQBnZuQLxdy5VtwwiGsCOrc
QQc8XTWdRsHIUW1oYsMakhwbIHs9Ghm8XJJ6NwTw2T7gWpiydFb3DKp2QpgD8Ek/u4KkS0Qee9Nl
XYmEngtraoApVMMAvZLquEJOy4D+V1tMloF1Na3/cygy/Qjr9t3Ank5aQZPaHPTgQBu00NWeW1hx
IUAM7clwSJi1Owsrg+MyDaPxlrf5ExmCGjmT5XU1LzlcR2+Y4p7pOgqqg7NMIg6zv5gvJkrb3alv
9Dy7MKdca4nDwi2cLBMZ5z908N5wOmieFHfvkeDGOnDaYPQUtXAbgvDvMIk52mBj4+X6pqqAel8K
6ogBvBCjMm38Is9ikd0lWAR4xV2mQbHHrVVV6rf2kG0LZ+yZ6DjP5LOXCvEq7fh18bsanrGE4VTc
ZF8rYr4tnDFvRT26hjaotCkqDGGZxoH5sAnh7Dz02S8HhYcnobEP7gh0ULLhQL1vWaT94EJgWCxa
1dSuB+1hvBts2RojVQhGYRE7SPPJZpjbKQea68Pxa6e5nxtCRInQGtrUAeNyBwm3l62IJ9R6SRid
mT+Skp5ZM36N0uscCnnZNjh8S0LUgTPqvfC83wZelaE2Za0sHSpmVmBAOOStUOOxXmzRv7AZBv0s
/veqDkkuzLtz073PHnGTjOfQQiD0V4Cl75K2VW2k2zx7wWgcW78+WaMyKFAPbE5/Jor6DrSR3hi2
hj87j/KhaBBTSAxEVgRClQlMF8/6Vwfu9Px4QovoUCHXutiRaP2QUfl4XYHbWw54AyMSBzpYsg7B
XtyNSHlEc76iw+kNrQuoOpYsb0UxPGS9P6FRk1gtlvl0k9OPyvmTbKV64ROlrG3kG4NFeT5kbFTG
78Zfoe4l0sTWOweAxVaxNSpAsn8K3GU5rT9J8Ly8msXw5RamgGMvZ69qfeNvxSfZ+7SSsrLc5/o7
iYWeuLP8AjYITUMj3+qZnq9xevMe9PY/19ooLtPCDVNgjODRMxucjwOCELgIKPaRZXpOG5ND/rGx
5t3aE8iesQsTR4RlmJPpsPaGFvrV+OXnkQSymSgmDLXCHqnXJcW3ZKHx28ZQJRGhEVynC248BTT2
uI/WpiIA3O6jrxE773ofg/esYo4XjgX9OcNN8bf7rZ3hzXMfKOOshTBcgs9GlLyl85sT03B9wY9x
t4nNErVmX/J00rveM4Cd46q12SVdbXYN+q2XpJ14IIVfP1UnjKA9rpQR30xfOsS7wlIaGxaMV5aB
t+Dy5vDHnCIzWzDgXP7qSc4h9i3Sb03NwXMCWAqs8hy/zUYzX2XaB7ncchvMlqNB4lQyGJaUciA2
9PvGwa12jKGF+Gi+c46ImnjZAtgxZMYtEzWYYNWYh03nwuD2IxgB67j7ljIbOqMVGPypJPxEnWHH
nkFs5vTA4wdHtCJYpL8bU/D81toHITfGuWIBdNJOnh0ePP7DL5PPmk5mJ2abosoZUkyiB+1Elmt2
iG8Hfw+NP2THobZo3L9ZJnERgv5LOGmEHjoHZcV/URmNGHt+A/72mJ3r2q1F5dbdU1sqrH6ydWrK
xFZoKgHGH+JYgHOuGz83PgOcGKWxfRaJMNagbkCflq6KRMlHIibfxEtr3xtEfuQAqf71wSzuYqKy
9VFS20oDN1UncH+dF9XBukedezop9Pr54E7kuIzMOd5n4jyajCNDZ8uUT6Mz9QJeFpnD0t9e2/VH
ftQ8JPtaIEQDFWAXFGYO39fH+uV1VHbIyMXVxQhzzJVh33dBQ7bIL90maVCwjc7BCzKQtgdmOlAP
MtZdt8Mj8gPMu9HYmZYIavhhm6jERrzWt/koUW8YtaJ99KRDmQmEnm/++0y4y3mzVNeonB5F/XCA
mEPWeSAX/JHMRAn4LKX1GZmTDu97nG/59uHXXPm0YmZso8fHaPy33Qs8eIxApawVf8oSTXZlk/uZ
c8LlH2HUWBaXv0igzEDcleaJm/udTPMBOmH+qtbRPDmdrPRsO9lW7WTOKZM1ISCwJegthtt06nf+
zEl0QGnKsl8EvwWIskh2qDvPfmAipfKFajA5YzgD+cQ8njqEML9pKQOfPtrw5rt0tpXQkn9muBCR
50ZiKS1mnq90cWrjSmPoKFaay1BRHADvWffl77gJAfSNN2Az/zSnoTeI1KOkphrTv6z82d1io+pR
qJ5cM+nfM6HIOwoF/K32qP3GeLF+mZ19sbDACMjtyy2d1UE89r+fB/9UlGEXafdhGv/mExxbv3OH
SAROcLsQY9wAZRFnERf0uC3vAbqg/H4/uhS0M/TlCM3rcKDTW0jS8BJWC9RVD7JEvDLq+W9mopGj
DIfWCcqKwMYCQatRmZfgjSdC0T8S796AntCLxifStwjOH+STNKJIWY7kjfrOXAErCTylNOG2K14g
M6VAe2W9OibknmwxZDjgWmbh2B8xEtE32ZNgrNm7ttdEwjirfiGemagpmoS4psk7Lg5IUdTA7S/1
6KWGv7FucRPZn+w117opLrt6CSNtemcflihhs9EUAouT6BdZS75s093VZIlRDdL0kSzYqrLAGQdP
c5UXfBpsJyynQew7T2QdQt4XYtsFvQ2ukM8thbs2O2vLmkpN0W4j3XT35F3XKtcnZ1bM09WRhODM
TBUKtUvw5wY1Y+0tkH2DClZ1g0MLZSUoxm4M9+L4opUY24oebGC+MOGBaZx/RFDAVkv09sEKuVUA
W00WugUAsR/X+MB5O3GvDbn6Lxv8nBj4baf4ID2w/eRITutXn7D0limErxNO84ti39Y0veQv3stU
YrYbTmclouo3f64pwuwNREpAAC2HmyH1tuIuJtJe/aRQX3/Ri+VdAmdn9Ap8cpzNfEoXMDFjv6Hf
/Wnez9cHUnK2UQkvopwHPG+vRJ6mc8Ivl2exhfrwXsvIHF8Crpt6PuKGvbPHHx3zM8onTXkYp9t0
vflmUDChce9ZzKWtnbyMCEcAG7MbQN0tIfjCJhp/zbJAgUnLBUlub9HbwWMbHxqRja4WytKAlYAj
cPDRJucNMd0WjvnRGrGuQw+tJF0Z+T5oHxX64JxAirLdHzMa4yZIJUPjJIAEefFKdvxoqf+EyPf8
01057iO/5E521C2tyFF54OYr5UL0suKT8DAGm55i7PsCveEOxkoSlb6VtgNktR3lha8BJdJGi24t
Gq95aZnlf8CXRiBT8cX7SRUuSCgJ6lf6j1zvwCgYWKxC11DxjY6MDSLvCDf2zC3+mpzIrgZ6wOyn
yzGy1aOeKLWshuFK8jIuNYxDJiMxiOpSYkmliB4hb95+nWX0OCViFSOiro0Zh3FVhjQbhjvoOfyU
BUwQQQvA8kGFgdcv/ajwSEOcI23ZVBSVLQGxfkdAqWbntef4RYZS0/CdJdf06nkUEWxD0pnvzrKP
t41qHEV7TjPU/klB+TaEof4sjqezUdwV1NNpBxYjCKoJ8PUXsJthWmZ1ddS6yJuK00WbkJoVvBIv
pU34vlgE7xnCSpg66xOlJxCePjlzSjdUY9EZuIAqVWmna2aZaMbWK3kCQ0m7cslSVQuSNEwjEDBj
PhsiS1TtvqZavQGeyPnXbYtQ3Z0mYcNy6ILI00vpSD1i1mM7hrPqEqpjJG/sS6kgLXUKobCKFE2i
MXnXimJX5JM6vNl37PDTxcAkJcyS4jLTGB/upSS4W6Tt+7VWsbU4nX1TJLFX4S/bVsOujP+FmkL2
f6G+WuiZO+5XaapKEW1G6xu1qX4Cwk5blVH12wKBTShzIW63QwRYTKeF3jL0eFZiulYGqK8xS70+
tLcPvyTDokI1uszgUB1SSoV5hkLdr8MiTSNBbGwtG0HYS/wrgvny/ikLjBRbsZ4EQ0sBN2YHSPCI
hNpVE5sMl3JCA0Pui29CbyoRLmGF05UZwirD7qr98oJUenH7iSmtAb6AYVhk0xnt/hBc1VSrPCv/
Xa/lUnfWQXEjP5H/rZBdrHTIcCcDn9erTTc+LQkbZHVUKZ6P2Cx7DcWvZn9d+eYufwP1TFCO5dCF
lbXbphzymW3iGwWR2HizvT3fGrJUF6I2yEb08By5f5+bmYrr6yFknbsDxGBSTAKcTpux+ZdtXW5R
uBRC0I2iy21rcz7ZOs83MUQXCapUdEwax4xCllPofBAhv6wykkrftLztC5y6lNrG7l8fDvxEXstA
H1Bv7uLRcYty2FP1TjruyVclYSxkyt5fOd8l6+c4KLuwpQ9frTo6oPTaDn55xiWiJxQq1n+BAk4f
A9k3s0pW1NhUq+TTD1OoziBu6MxheqqVirUDCwRoGAc2Mee+TVocOqQMwxOCRCNfjR7hBHXJYCSg
rTq6Df4Dmktx9AZHYiR2GxCpdbAIZTK74z0hLr13KuGp2admrJhvSaIQ+0sa5orzhw58QE+lVG3W
5asExxPp25rOb6bNLFOf4cORtgQsCul642iDFI5FDdXUTMjYgxz0P5+v6AfTq5W5L0uYiVUd0Fho
5ENF/QIpn6X5xes4OtjrD/xvlfC1372KGLdBFzY975A/gqPEXc94B4Kf5UWZzjHl4SuxxVCpPpy9
SY4Koar3YdWqfiEfTkGG8SPXS0hBwh35VeZdmSlbGqguaxvB5fTIB+w168RYPbLz7djc93D0Ezik
Pi6YvPQCeU6ki8bv1XgguVGdoXYPyEwXuyVFJ9MCOGAly2UVUdSKdr0dLRWmXjjc6asRKIIZfGwH
911MN1dNH0NgKPKWpZBQ8fG5UZ+TKMWOZYc1zmX1tcF6TcllfSJqt9PcF470Mu9UEX04CBSPTb8L
VbrnLB8Ek6x9sMfyAlzNaFEZQzvhG/ncpO+pPk+nx/xfSxZkej/qrpxMLHZ0AOAefsqgBZ6yuVGu
Srdff7Y6MS7nS43LJPCm44DvEXZAgbnPWrISQAHVoMjtxcQ6i0DtOD6DKqecDOYfHNxRXvIYNQad
jwVYeEgBcuQxjGtKvEkPbDaMUrnBnYtZ0AipcI6jXCvoV9/MwinQdpjzGumAMQZ3veKpm/CekISs
0ReTxjDdLQ4W2pR8qgqza2Th6C4V2uVByA818dCnhBhfQDUFvtlI3wObNAOteNOyMdvKZffAbaX8
gcLk/E0eavVuPG3GkViJH6UdJgGHZXP5eBiK2avi2cj22BCGZY9Fem9ac6r0cQj54jtOsoForQTN
1egIDcoAFCJYShuxpvJnwjz5tZy7gKRycKRCzCgksiNY0qPOslL9cq5f7yxtZ7mh3YLtv8hfblcc
KzzLD9v64UJyXjLL1zZWr9wPfd86s4MAuC5ToUgh2VLVgrvoArwJkwsBgepQqrL9ty6RhLzh3hWy
wftam+SpAGJ1jw6TaXsbNSE5hH60ITASf6yUR9qTPtCEu4RESPmM9gfq8mh5tOH+9YuaAI5IeUUj
0Y1liCJDGW4BtWg7rMMQBFk/WeoGakJc6+k4tEm1FWm90l/+JWtveNI/Blp4HyXRDvNORPPL0zo1
LwmZb/vuVN8oC5FChXasZ2bF8JabjIZouEs8bcrB4sR3ny2vPO/Pbqh8jUYDjaWV1BQLVlkmd8y/
+kXsGkbINkeCztE/4dsyay4S6KtqSdSlxge++kyxNrRXcfV1wwNe9cIyAleSvEcuZiXppbeSaCB1
ZNOx9qHjrYM25+nlRAHp+yybiVMOqyes3aJ4yz3YYHhkM15vC5qzZ0Nhm6NBa7UteohZT+Gp8/gY
TPuuHy2JNR0bIzcmYG47+SuI34hOK2MDCKtgx4QVUxvHTdGjbbK8r05iIm3XpRn7s55zSPBvsUNY
llsKkPYypha7r7n8A2+BApgtkr7nm7RZd3UcrFTyZ1lVWFmATK1RRiafianClRYpguwL3fsivo5C
p4QYWd9jmpD7gu3Tz73ybUbkT08EtUT/0Hjb/TyRQNne6ISm3mALeh3LcQVJBB/nNv/xddaEE99E
rh3+QPTAsvDZr/C1lHmA08s13r4V0Xs4VY92snzRvk2GJlIJppxdalKFmsFyqPjeRz5bA2GKEqFq
Fs7HFqJ1dyOAySxXNfFUiYKYe0xsi4nMB3aUzi71rIuPyx7g7O4x6Dp49lFS5C+2YQGBEQsdivyg
gsurytaikU0Xwgjy0/E4xjZmWDh1+MxZPeZB7j+ZOKFFTVjAn+udqWb+ZKRd28ExehOGUJMg/OQ7
oNcGW22X5Hjez7eoYtz9KkN03u46j35Ts5Vh8kHzhmajV6HMsWkjlzo7io+omIKeXcggF3PTMGk/
LcYsQoFMXg7huGBsM4Tb07X3uU6E7QimYOdh6yDK/fjiw/+ZiKYyKgxgaY8d5R2+eK5/kmnuIeZa
cskMvyxmeKOiIzu1+0xNz4DJKDKzMYx38nAHLoG7Fkv7J5hP91ZXQRUR5qoOHKoKZH6NnICe/jDp
xCXMJqEDyGmZ8JBcRUvuty62+QbLUJESKnVF/H9jixiwPX1X7q15gwt1PINkDu2o7a2jkqWDrMTj
avjief1AEeSpsZVYDLK4wBvasXlHoOiFQ4MCVJtPMZyTetYGu/YxaqOzqhofgQloLFHbTysHJBTc
i63+fewZ6yBcSfMaO8PKWAZe6JfeznW0os03HIIxtq+YKFkpU5/rOPP9foc32WbVmwzZmgbahNje
nG+KZvduuX2mzsiBGIt+gFn/qS+vjZ3Pl+l/B3GXe6Tly/MxR/dNL13Co0KfMlVXiGp79SKJarhx
/bL2z4t/0fEYQKmbcE2UKylLWhqenA/MxQNRpW4ZA+kXQ2BErwzLbV8fGnN3xQlQSyQQ1OotS03h
0PRVMZpiT4PRCAFnVwTQpJc6nyL4r7VW/5vIxk5Dc7ASWpyA2yFahAsDFYYiggFcOpeU1RA5wuop
ms79fMjPUf0JUnEb8OgYjlud/6XDE9K6PGFSGLnJiKA7/Uf1cPC2VJB1I493vjNe2O1IfKJMyCA9
nuLrpXPhAETJUBDnMGkMgAE92q+L26742T/yT5O2gsS/uU3ZgvZmCFpWS9/xHjfhfYMG8Lbnf0qm
3p2QB0shncdjHeQ/AI1Wt0bB3SyljGkgloSTvcTjZdq18nxYu+v6wkrdykYR8xbA7XW1fCH0VFM/
0grvCnFNPKwC6Ha97HWZYJ8tWDnlyoW22bdyFEwnrsKnaTvAU67NIU+CMQkK66+/QjzlnuMrV5UB
+2ogQG+zGtviSAVVMRdA0iKK7W5CFoZkZZ5oW/lYsGEBHMkp3r9XOx7V/JclCrKH6cOGvQZX98C1
t+XM5S8STF5Uu9DtjHi/MutwZMiFSITw+LklR4aNtf7CQeSkByy4Li2Ai9qXeDTHAznuDV1bRH4k
b753zsmmIZE3PyPvYtTv21eep+gkeE7aGMY655174hwJSGGMXAMHl7REIKKb9F9/FMqqhZRh9nqU
s8anl45+HZ/lX3fWrQn+tYeHSlixVD51hKUS9UCrp/+TfULi2dtD0Dsf0YeKNpGVN4z5YhN/KZjR
CBxV2Vg290gKAdhxaYhu+nQ9/Jo7Ryq18vtdhdZ9jF3B/8YSg3WXJK5TeDTIbNte0vPoDsRPHptP
6RsqT956Sp1ByuQWY7a2m2buhXuKUZz0tXuBPXbeF2Hin3E4KQXdf9XKMDlJKQ3AEoHw4ag8hC5x
jfCRQa8Nhh3xJci/+xOVEexuL+O4RzDImAWaWfv/mOfbJURAdEk7GyYiM414HMAq/hOn/LwyS/Ev
S/2sDW9QzMQPO8ID3KqGXs34wa8a6ynjPr7GG2DUXjNSJCamd29qhxou5TYICgqabs/0MJ4d3x0v
dfR4OAIg4RCX/F68jaskzqFpy/0qtDGDSAnv3mOEiAu7MNY00kJRvmkyumi4snT+W9u0DJBG3z1E
5G/fhNPqpPzHDLkwvOZ4t/ATmyODHQ/+PSFpoyQf0IA54dKZrc2DUjGtCWqxRAgYg/4AP85kWDbP
591SxjrgdAhXyUHFltpCOq4bPQ6xkmSTYGqEVVECSL6adSGY7Zl3PjqEs+PIhQKRULV2AU11RSUL
JKOua6QLYlAWTyFKTAdq6JLp5vCAYU/7k4gNYgbpj8zHdT0Jp+GR8fSoJP8ImRE6zVKAOIRjG6UG
7FuT8AwtSZMPrTPLctQqh3gyrITyV7gQm/8UwuJQ6PQ//FP2Swf2hZy9xaibYSjcT1dbHtrbl108
pLJ6QHZWGMKxzzmi+5kKYG975vf7wIVMm1aCTcLyOZhwlYR7f45pnfDKR7wafAoL3kKvTQKZMzOM
d8IIAP27apAvXN+rXhvy/G9eHCS6UT37Xz1Q+QQbzUbbUnj1EZ1yil+Jvc78d3RSxICeF5VCQtbk
5ZXL3qbN1ZGLNEvQchhHTiEnYZV9tQDJE/i3T0f4cTVwVxE3QQuWdU8AjQ016ybd1/HwLqpuD5XC
v/i3gKqZZ/w1rUONZwxS22bvFct71P+D16RsgvbA01E9CXyUqk2ki2UKU9zZ8alR6Bl0KGU3Zono
OoVlay41FasjurRgGvzgJHlmaBemNf/8CQcrl3HtGci6QZVBFOLgMpmGuCzRx+miC2tmcvJRgeej
VZqj3VhDsqsGXyNk1NIBhDi2PIlE+iAuKS8eTIdembIVPuBVKS0C3pUpPPHtYzmylVI+X5QbAUoa
m8FqP40zEnHgKf2Au6Rxs2LzvNoszWn6oAfKZVJ0H9yR/0UXONUNpaXBYYoh3IzwGhDAuCwDbLWa
71AjOdVAY2wuH2Jsyv29WpeWFA0xQkp8r1VcqvHKpbUWwMVwYmPJPXsBF7oFDcpMbKVPcfVoqGBs
9bNwvLFl0jPoQqilOB+iCD6+wZheVFmvw/V/9edoq9/BhdqSnW3EDitbQVT5JWECpof5Fy7KuN+L
IIVjYhVbAil7Nlmaf8HJtg7pu1XvnTyh49ZZMfet4q+VJyNVRCOQ02VK2BjlXqk9qrmJaDNTMmFV
yew1Ody1UwWqzpy0yVVG0E13UeNlP+/z1BRCuYkHAIOtDP5OI0B7wipNqErmZYvScNyddpyrU0UH
fB+As23Sp4JEFTCkqga3VYaOMIW6MlO40llAhbnHJgBtHdFvA6o0k5a+4e8covUqiPTdrk/Mzf8s
NCbcqZ9oVTstyp//9Ag9Z6qsQ/mFEQ4hH1CQ9xOybj72fH6tYP+ddpruN9p9UeWMRHW/JW9iPdEf
IEfC/AWXGvxzDezjJdwMJf48s4KDVJRGclMOGkJXcttobP3ZtObcge9tb4N0AEi93W85wWD2tNxf
GLRD1JzIMdg6hcQqvuwDchs6fJFfrN4kP4jPQMLeyTy+ZDGZ/UvRESHiAn9VT87r9yMemmMxW47m
Ck6bjOtxHIiKGkkr5LFT0/k1j6CzTURyeBsOMfNviQ12OUWqQpbqSytmG0OkbN9d6PRK8kM1D4oI
L5A830vL2NrXAEAAD9LmAo9IfoHlrMHStcSKJCIrqR5ep+jNwpHRyVtu/G4Y5zll6tOTWMsxaTx9
ufDntDhTjLykPkODO3gigcnmh39Q/qB99KIYdTsXvolHoTVGP3ujkH6+Tsefer0mvXWnMauqiNj9
RoTg/Va9QkJniVKJEJBuJYL1XSJQvq9r7ZS7ip2KOgXwLpydWEc3ukQPS5tE7Doc5cdNNLgY8EdY
8Pra6/MigQaGBsQbhPDd5KnuPLZEpNYhMGHz5FzmK8CeawYXoJOMfs0QleyXEQ1NkDpYAHrXb5jU
THH981c8hbHRoglNN0DDhQ7SqnwzxcYRhfaXHSsKqHSGqcJ096jXatU+7JBp62M2KeyUxv549LNv
CCMN4pN8O4fJikvW9+me6bgjLZlLSuMyjLyO7aF4+X1SLIfFkfBeQG4v3VaqNl4C0x4EhPUP3CIS
YxSsVb3sspr4p6zGvlItwZqM65g6Y5TGkxcp/furkklkgD340Yb3aRbMy0n5BDq3YIq2pMX8hmqG
/9tDLJbnFHsyeEJ09RahExTnUtUUb6CCiy/91PJkH53aqzwgaW22OCxJZf8hYgaKlJoau73uShJh
2vyKzhJORuE2mQkkDEM1LtEJjDbyTlrrcNTZ3zlOuMcgya2r5yJENOYVveeJtulF2tYUFT4Q3rcC
Lubug2padqlAB+Hnvx9qqa21BzUEpM6qIuTM1re+91IltUddoqRvzLvF63xRmeh7iUxWzEnwn7ws
CjZ4dYf1/klZ4i2iJpDe2V9ZIvUpudUTf7J/isJe1UZ8LX45gHxZzQF2jHngyHRcJuNzlWxhS9wR
zJ+on9J0nvyp0TxBYzyzwNBT9IHW1doohU5hT2GNaR6dk6mKdlFurmHBGJ2G9E9pJZzCEjsLTu0v
zB+DePdekcYvZ8sIDwqlDulF1W3W78YkYm6sUo8fD06PVOkDUWlLFWyXMa7pXjSroNsLaQjf3urm
/sxy1YVOII1QM3t2JzoHSafgbAsJ8KWdtvryJuRh+8EWqFLD/w8Je1DFtePCpgvZ/kFGt6mXsf0w
s8MsCfUXP/tdWeBsocrOImWKM3UZsnVQzSdovS6LRlIJ53/OpZNP008h6MX9m1kA+q1ZgiSr0Dq9
wN5ZslH70GJ7xMsCGkZ/dPop6YnxTZJIf4s85qFG7meo23BVO15LNSC/1T6r+loh9kCS7U7Kij3g
qSHHnLG4KFcEuEfDCLpjDOeX/zuKAFVTwW15nNmu3kugdpnod6hBOQfXjqTRR3SshfgBy2dmWuTf
I3JBwhHKg2s5iOFDp3YDOUz5aqDcGiefxNP7z+oMDJtnT1+mKQtdOjAyJBui5VVWeWdnU1KdTNOp
LpPGyJaNMw+wWN/f7Jfc/xHPi7QWDihQ00JtsQBTEYbB2oHLKH8oiX/y5FtMGnnwp2Xaf0pLJgNo
MNE/DgEDLwJ6m2bnViria8Fa3PtD8LCxA0ci0yENkQUUyyjaEBsvw3/s6OjapDmg26i8iCbSsxx7
x32bEr1z0hcg1bGlJZuztWH1pYFD2jUM8Z9WwB4Q4PCaZQyjuBmV7lgifWAjvBejg1t5XIGfo0zA
kBgl22ARnUp650s31KlRAqowN6tEel3hu9DLYeU5AwLSBok2sZ8CppctbuLING1xu9THT+6rwA3/
vHGafVjK3zxb2yM+2fg56217Trzdl7xpCbbfcWhUwfJjTiGfsMgL6KcKju9fyX/AAMS2GC20WB8i
WG+mk4JgmIbaKpbxH0hC1M64AjxuzK601f2vX2O8H0aCY6rasa+zP3EDWmb3XA/7cPsfJFHHQ2eF
GAcz9BbmoKdH7jjyiXswsh2g7MFGRfXi69+1EqFOZ6gKDgK2Vs6XiKBYDcwL8IlKXe3rVktvGjDe
wluGX5ffzNvs2Nl7Axfef2W3fH48/JDiRak34WTAJEjO/6kKCnFRgyE6HZ380AF4MhQOx4k7LQy0
p5zAZh3NwBvUltdxjLe1Mcy5k4cJcYYS78pEkwUZuZ3cg52xsimeIJjSEpzagL6nKCOL4VrfngK4
tTEyV1IN0tbsoTlgVJEYHej0uSu8ghZvQ8weUzVSqMjpvSL0uBy0/cue8ZzWgwo9nu6nKvl+hnl8
689b8SLBIsp8CMFv05qWwGKH5WZF+pskHlK+FhgYsb80cLagAuGZtkBn3kksD/EtPj5+TkDRImB8
uVQhFi0UG9pt6pcSTMs/fOzSK1taSB/0hYZM+9MzbLXV0EgWCRAQXYoslMfVaDZ5q4z0yt2LoGbF
7p5Uj68l2szOjfacP9bI/q9nZHqJq9C6UF/Qb8tyUiYhgWcox4K5DULwi/lxPikfBCRVUfqknHji
qowdUk1f73JgslVga+npH0IF4TujERoKP7xAxggnYYDIUu55hz+DnXiH95e4HmUezNZ81JeNBaA3
3ErUUgd2CJF73mkr89VcP+0D19qGUSH3CkCkPuS14NyFXeau+WAq2joeixyj0hUTO1nrIH+yQP90
Znc5qA5GcC2NfR2sYZfUTWyE/tUhCnvUD0CJJ/0lFBkJ8BDPozntTA2YXLz01RXql7uSaSQUVXaD
YjJ6AN2ep7YkK92+gajnC21/eior8zLcmFkjqUOiLK2+gi+LP8Uf6mAHMmu0y6kJrvhNGMtqTkMq
BFCW3P+xAturaQ3GBA5Kd4IB4Y2RXIjFOt6jhTYqvEblzodbSL4TTxq/czXHbACXRF4ZgHj7QGa0
8Vr0BtmdEOjp+kFp4fw+v6X6h9TGFGSXptkgadWSsPg8AhzATTWh9yPfkrfxRqZSNj+QgqVBZpkR
B93sMcUoX1MfGoaXsXKvdBE83iwJThrzTlChF7AwsZ2kSzW3Xyt/5QugmuApKKb9jh/Utv67Oc0R
fs9Ui3pZqV4ZHanKTJQUuZopkbEK4rn5EnEA6RjKKUWjeVYDc9pGV+m2boFX3NAYU29PNQwIk3p3
ZcWzVu6u/ELdGBIwhMZW3G6vo/By2hYlvAUOZu/0i/mIVNl4ik953XT2ovpiySx1efOczbSjuq8w
iqPEgK4Ec7QsGeUswUSaNRE7n6RiEjaxBRtsguYB4dt3nlF1+e9YCWAE3hKwoSEnwwXb9pXXTBsv
uFcKqydWRqEpxNb6GZ2IrWqRPN0glNfe3XS4GnIVX6zyFyV/JoQC204Ghoi9LC/beRsgWyAToKdx
tMe5GFRVq/SLliMulyZHwBFFP2M3ONqBfttlTd3X61HW0jftRef3tcNjNDbQ7P2/ipc640U/1NFi
POApN8oWux6XIS3ukRhmJE1dOgJpadr1G5Bv0Cg9M1hu7LrMLKchxk8M9AEYuPBGrlTNHG6Pbj3N
i9QURUIjllg6zT3wyG9bFwuVqg6Cag0+mzgRxjtq5TYhLI986gRJv/LMsoTQmj36otDOWwFZTi74
ONI3r+Kl4w0nPmoF0H26VFJCCD59U5dmCx5kLSXEkBFKggqnphHzHUU3h5o9/qTd2Z3byfQ/sxVU
TvRGNlHTI53RSy7aP5hDMQJoZTZxXjpZDfIo0CqwyeOLRtH1nMLt+wZJPawkztvnFSp/dUIh/nKp
/xAvHagv/9DVnIoHDe77zE45R5hcl+PbNuulvMjo2WrkuzsmIK1wEiCPKDA9/JPM+OGQxpmUUxoN
+xehkmyoEB6eA2Yr8Uq7UxsiNUkysMjtE7kpxDKqBTmHLqdWI7KW/Of65NMPDWamim2ihtRCana/
I8oryBYjQB0cvk84eetEWs9loBYvhOoioob54FFRXmstFD12kQUysnf3Dh6I8k0dsHaFi9kvl4XQ
imPVbiVUPpEUBt1GyBawI0doYEkkw4oIKkY7qpd+IvzI+egJr0Wk8iTSZ26dXV3TC+ZRxJ3wNAk0
cGjO0Upe7+GvI0v/nhbBZr81f8JD5eJNWew5RLGETQlVj5pUiJI3BhRXMcjMvrf8smp210k1iLRW
qqGUqrr+UrKL7gndi7tUqnMvmBkimtKKVX3zhalcAusgDRLnkx/Gkpb/iMdrxOm3L8YprIRAVA90
ifi20aAXucnvf5J1bQHQdBFIkziUt0/JKtWAicUt78xsgjTksFgtCZ/f/oQHoZ8mZAb0BacjiXIj
oEWKXNTsxb7ukTBCs60w2ispXcYNWx34ycVQWKdqpqzoP7IqNLdMTPwGxul4oQgm50rmm7AT/j3J
JpMvEQbIWbfAX0b1GBJeV1JblQiJ1cbsuVDwrBMJNkNLhGyeo/BStGZSWGm2aUEslll+oj/6ht/t
xaqgd5LCLcac4r99lGGBiGLw1B5co1cZpKYjj+BmAQIFR4d6Ri5x3XYnxaxpTAcv5qY8pnC5+/dm
QOMFEN4vM7NIbrwoFDLNUoqq2SEw842ABSXYfJ7bHEJFt0eHv1WgAKIwRIh+WnIYrqf+yzelZjyk
FM9dLYt559hWtVebIzg6MVV110EAVfLvT+rmVsahjC7QnNYGrPto6hgpy/a5laNqX3zjbtjUT/qb
D4s8hHnYnbJyur4NHAOwA/9uW12/8FONCeej7is57L8h/xB55KzW8CqJ03cOJVBIdXO7qf6xEIVT
hzGjqMBkF8hoYLlyaIi1LIJldEBJ8a44VEUFivdTWjPQjwllNNkUNxA5QXmQRyhg0apnPJskXpoO
rig1EYEcPRT9posN5Zwq1YrRYZKbx/Gx2VdhCOxYr/5GsfxG31qRcRW78duhy1y2G1LLKQeSoSrj
fm8RkADI0W1A1fYqJNXCa8CeMwgAT2lI/iLgs+DjC1Hv1v9swNu6mBwPk1HWYEzecZjdvK60u+Qu
lW8evgfaADbM/GyA0w15KOhdIR4bXr2f0gPl0KzNUjSpJkOmDbsGlN3OgZHQCVhevkV3zQkUp+K2
hHnNmcs1712cklWAWE9WhAls4VUPLxdyida80aVRFikg4CwozWWPkDQ/S1yfVMZjJGeS7H/h0aBd
I0Zplr6GIwjpIWQWZOqDJmEViev+OZTwcC9oM+1VD1Z+nrRrf6+ITpBu2nwjfims4GSne6V/n5dB
fUy4q51j8lQ4SabD8GvP2meBoFR23+n7g8S3EKtlRdnFcv0SO3zBkQGYyetPqCOHlkim1BTXw1pB
5L3tgq0gCvSiTQ90ljboIZu/U9+PSr9rVk+UFYyQ1Zgp+ywZ4kmXU3jTIH5rJHzrHlSpjYU9WOZU
nZrXuUlQyUNtK3c+1N4abEW/K7yn20AwkgO1JiqYnh95SX0GmSXcpVEpoGb4FjNLDFvZi7IqwrOJ
YUGYNZOAz0UTNYSXFfpF0HjLutUqoIT/sisT8MNrwDFGikRv3iTgcLcp1opqhaeLMKKCX8+wUl2q
XTMmAQE4iTvsXRUqiJ2Emq+P9bOOOuXZ4NAuyGnU+ceiStAr3Q9G9HdbPx33ZgdXoqkwn52NZfjt
Jey2DLuacNHDz6sgQNkbd1Jvo3XkkRoK5gEyUN4VDcKu9kCX8J/xkw98N/6iSXufP3Bkil+tDtDG
BXhpVC4pKTHTRxLqDVx3xy08L4/kmaZ3slYa8mAzbwGLiEWh9Kcu9FYV/MCa4dIW65eUJqHsQS8/
TIRCR99yUtkBiGZfn2T3/S3KJ6F79iHDOLqv19bJmHgZ8VL0w9LrgfZrpROAY+eZiFkh0OF+2SQs
VLQQoZ9vuUnzvtmx5buMsk8POHkrb7bJ/yZDeim2OGZsAY6ynZ1X41NrTpHe7d/0t46/3WmuWsON
C/PEPLtajmUQ+rIExwnFOOb2ZJFqoeA8yMbma/edp4IWln2Bvtgr7D1nhG52IP8okVt0K7vl+IQ1
5CzW7PKK9nRygkOsNgaqEpeVG/TVBPGiDK/hFy9q/gIeNqse0WmP2cgn3t6sgB4myAyKcbwez8ey
5vLuObNVI3ioDsEf0F8+Z/DIFvy64EmN8Ba56y4IeK748USCf4elrmJdMHoTpSjHIo74/9eqoJTu
/SElVI3SAcZEX3XAN4phnB9h5De53ThMM3AYOGGOlIS9pVdQ35tB+EeTEy+oeUE0SEBLhzKBFTQl
0vSSsmNazjvn/U8W5lLq2uxf3+s840ngkEEHmiiVyZh/4Nl+y3xNvR89OipjpdeP6VM06WBMIMNA
tY9zLuuwU85AphJZW+6Eq2Btd2fWUvBtU6it6ax2d3yPhm9hRMmaYe0ZbXMQ4ZgVdeeVXg6a9SrA
o8tF/B0xMPfVFHs6YhSqU8rLaAqsKncMnw9YaW6XcUkLgGtSwtD8ysozkCRdMZ80F3A6r16va0WH
POT0R/mWfZYhaQ63jmdjWvuDSXn///V3jcYUOQLFj6Qpa2pipsqXLK9upAKs1IYaGfB9ieSq6vxj
2zqQO3XsAALSFVRpoigHvx6HwLD9RhNBvLX0vaYN1asbf200Mtue3JYlUa3epDofh8eb29fxbofM
ezt96uBBVvNuIvY2/t1f77MbS0Q1v976/DibBcuJCYkicKPAtXSClr5db6MP9qHG5EgC4RDPWjJ/
s9WB1+49sLb1fLtpWEiYiNQ1pjzSYCh16WvjiCO6s0nCGd55Kb6Sp3kAD6j16QJkZbtv9Z7v5f04
z7J4qJisdDtntXQJbYmo5iGXTSN0U6wcs2y8cw0an24vhhku+4gwO+InNExp39bJrn6/jykMV40s
yySNPA97ZBlJ2IHOwT37CJRS/lSZf5YkTbKBnKhAwToMXi0ggfkHb55XSt6XhIFV3CtZR1XUW3gh
uhab6EKD1x+67IjGKhaijfiv987O7EZzjm9/ieZijVtK9kWtbTs2Fgi9pUkz7pxd1jC/lDslnS/h
tE06VC5ccfgqo8S6U8hHjIjQ1unbzaFdSsVBhi7FDRYR9r/Af3bps/s9wOX7sTyGWrT8slPj3DMC
ycEuRYCpdC/Kef4WMwEm+dKXK/3F6L+O21MS0pXAue2DLo/pSsIDURJ+EhG04VFmIn3BBHqLDox3
t/9scmvjEqQtAKzsmCPPofzZ2rwl2DYRp5cfoerTJx3XMvVS8ze/PIpSX4rxhVFe3fhvz6xjxaE5
yigWCsINW+hLIqI/Axzak4cvHwDdHW2N1deR3OlBBPO8vN7PFZ10ha3/E58tBBWYgiO5YaO/b5zE
5T5Th8IZlRJDk8H4syeKQwWl9iGbt50G8sDYZXW6BkaTkHFox8MrtpzvapAZfDuZgazyhz8ydqDq
/1hRN5SEowEfS7QCqc/mvu+Gismh3KP2k8GB38TutpTmRZ2eoP6dL4cf2V/hY67YxxlYDqS6crRE
Z3On9fJNqshOQhAyHahItqIsE6LyxIbYbZVCtn1IxEdRUdsA2PlKm1TNQOgOAlOzn0FLT2ySldD5
9zA7aU3svXWgrAKWAPtBPMiQqKQbSa2rzxVn5ZgYY2ywxeuaPzQkjmMsRck2FQDkurJSl7an6sGp
DmqDDZBmlldj+RPUVIfHoh+HT2oxIE8XFeAGnyY0/CXiuIpMbuuMqNSpZsSrBQDuMnrw9aJyQgEm
UTJCdyWTO31HRLqMmQ1WO1hRwiN6HcjZaFjwrhc21vYCcRtH4zsYMgFNKCHd4qdfJDxLdryJEwsv
7kNGhAUhZfwupHOEvOAJ/KjZWy5+uWj82FqnmLuTzVa3Tcm3EVV0cksQ+ZjM2WSV0oWzKM/4/DPD
ccZMicLALvCboPLDu58hFpQRuPINsIoYepQMM8PjkuZ9oixuZUSEto2Jv/LHKUakDQJJ/3Y5n8Tc
xtStXTnLoOCq6mE/Flg4BIjG571eq5vg7SwpBYPWMA2l7bNxBdYIp7QqqxEjGdlgmX8ri092Osn1
dXVHSD7X85Qov7DJMxxcJr+XylUvwDxFy5diM1TmB/P68KukBUDnU+RyLTiHY8CtRkKPVGy9U74o
oGERkOvQ2Yaycp9f7bLpzqapImx2ejB6s0CrzeV+1rgppVmwbFl0u2hOnG5aReCd4qXyLEoxgFrc
wjDbEs18rEa3Ko5t4EXbP7gkz5kaz5evAvUnsllMF/ONOP/jncOWWciCK8keKZhtSambA99FJd6Z
p0x78qJ/749v73+7dlTksVZVwz2cIlZObYRKLhGm/jwbLVtJhNI02QyjbZ1Ht1lkuzkrg7vSP9Zr
tKbqzSeO0E7m0AQx/PUvCbjTa0YFBRes6YBjWa5o+LXgtIMzrcKy748MzNqiFQTIt31zzhYnksm4
wGkX9Q0O0SxDfvfNzM1sTlOn2ee4UiRgNhdcDqCa8nMrI+Bo71Ak1Y9Lx+gPpVTOjKeOd3i3pPGJ
8IQ9RORLASgmULRI5Ijj9VB1xhaTfEch2nzyNS6LsSSIIm8s0pmnsNgq3z2ICBf5gtPTc4mlNQzi
dAAtNxrjV9st+swftDlSXuaj2taD6EpH4Qa1Xi/6Xz1F2+3nMLQQPcPjByH/9sOSLGKd3kYAWkFQ
sQrYgNhFEtEhXqCl2FkGmhbtneqPflKDZgCOs3IK3AjR/qi775n8d4VNnzy4lpDDruIpNzIsviwX
TgRvbTmGYwgaWj4ik0aBsQJs9gbGKt33Le2evFxhkMKaJB4M2ICL5ePMYgq0WBPZsHbgOi1TI8h7
DioMWKAqdMV1psZrNzDWUV6dJQr8848TLUSHt+fPeegZiRPedlpcCpwiBfK18YnewyK/QRias13K
rbwRU50RHOEBLg5oGSZiW6e7/s0233bpzDXu84m9wW6NQ93SN/t9xzhF6rtU6KujzNgUpx5DGAFF
1ede//o9m34uokngjJDebSIPDYpBUQYZwfBvNuseMRPOjMRusJf5Rl5GefiuklxrL/DHBVpERbhc
Sgs4uJ5O3fsFf4qJLsL6Z/tcYGYPLayKwxJJJGb8k5z4VZYx9Bed8I3W6MnphKUSyVdY7ib+2g8p
lVaQyIJeI1Q7Dc4+J5vuY/XQCqsMLZmmy/oBJN2boYv46Ps9U/BUqcS1jMGd19Q75Rw2S/YyR6d/
wURagfTSuma9xL0wWHRpo92gn1uBUiMx4fb/qXu5/5Pfu4v64sEskc3VagcRMBmTPxyTnr3FWjP8
EKQws7sTs7jZh8pJG9ZHuUGpYrBtf35t/vovI4aNpwCHX3yawoAoSf3sHWMaVcoOnixR3LzPpO4a
5HA4zGKr3KfyS0ar2EPA0TrljRb/6xNZ0YdVyBwcfK0vH+BwyX2Lqf5+Olx3epNlI71Y99ObwXtB
n9Vd/mV0KiFxSBE/fVtrqwDzV989ZljK9SqfvkTkgn5/3560RNNvsnp7snuDOctZRu9dZdTWjhQ5
ScL6G0z1T7f92glWj0QNAGYZ9voj9fXpUfrTXrLQwRX3SQFhuC6LsAWf5Rc6Wk1PtGQKTfkPIOf8
rqFls9gN6FQc4/d3hInncqERJ6oOb8q7sKPh9PhUPt6dZWpVaejcZ0y6DpnA/hp7rFa4qgXuxAYa
DqfGHZgezAHalHwpK3ZuuTeZp3UQVM3P/QxbLfwbQzZ6gcOs1BanYs8OlSLdQ50jZj++3L0LmY5/
HnG+cututSDA32Vu2r2dc5TnX9FsGcsJCY9gVEy8sYUvC7GCn3qi2qUY6D8yhJvxzh1g65WAwdCw
NY46AzuKZBdYMVKUdPhwPQFrQL/6pdb+DMRZzfM0V8A0MZ8DGEUrsQeI38X0ZW2sVM1Z7biNVm51
Pjnyl84rWiwFYWjkFMacRTRhf3MDUBaCQC8rQAASpMtUrCEUnHebx0mTZj/64U0YCA26C3/EoytE
Eb1w/cERZ2YTM+U+KbLUEGF82B1MDzs9tUWLAtmBj/BtXEU38Ml1WqHzE0vy9lh0JuLsT4MpjSYb
to77FXa7wPgkAeq/QnYHChaPpV/p9FxAEUTgSWPw3neQEquBSVUjLkZNTIZTsEPjNiOYjk/X2xw6
3m3L03Nxy2Pg7+MKcc4p74xCf/EnyayI0dHtOZudagfVHTs99Key5JLZkZ4PLHeNz+7HfPhitheZ
v+/9ls1nZ17GfSCdHntyzgd4H/Qk4SU/A2Ph8T2VlHXhmLnZPOgxv+ycF/cl+hfm/G/5DuZUuAqv
BSME9B0sVvaTUFiGEM3m47gSyOXbIWrO9PcWDmLii45QuQlKyFJdm7QHMvsxiB3xOvU+Y2m1Oly0
qD3OFeT5ZVwxBp+vCrw6hxBOQXyxwTxOgv1AGi1btopfnMvbCcBz1iQhrgnq1tAztJMfTdZ+JtBV
CcvC+IrBHYtPis+tGyQaaioT8ViQ/CDn8MAEPZ0qPysCEroASYbdq7o5RLf/AMPdVEbmw4bFT8jQ
8jKHsLx3VWbqRwDK2NPw+jl61j3QCqlSuxkq74UvmIq4UiNcpgIT3c2OKB7mYYd00W0FwFq/D4pM
DSjP8czuJmaiCHUSji7x1nAOkgsUAVkvp6Qei6E+LNJ2JpPCnqJSGHhb/FA/Yi2TSVUFWpfxywtE
LGbArGbh0ZEBej8Rwv+2vs+WoC/wmIf7l6GNMHUXM4tPiOlMCrBdjAdMiUBViTDhrjXJurtsV6pv
yNmQww1Ti9+sV61MFXJufhEwM0k7FiymOOfUZhVtsXYkAPP4kMuY1kvXWGBIEXDo/U9NP6K4ACC9
9yzyea0vbBtMSGZu9MAU7pMP39jv33WgsfTYfsGAgZyiXXyDfnvCPtqRl+zPRpybRxQmPHn6cHOf
x2XGNNVGVXuwaRDEqy53jaeVK0Lltbpu9gQw0TNZHGJDpALT7Ix759ZMK86vTmXoWKQi0vZ1fM9+
SmEKYr0/daWgXnx60etTNm5eZPojydhNYCVNbgvlD3qQsr0qmDyEOCKShXnW6v5v5Op0UQWypc9T
jUBrXTLfOyDbs3GOS9sPALM6yTlGI9YK8x0IQt24uegVZ6RFjGeqiwu+4ys91FztSYq7/6WD0Uv5
EQIxsuhKiW9TdAX4a5gHBV7gyVenQn0g91Lf9Tj7g86FTID+qmWqOLp9xGP2D0hfUnop1R8efAx+
MwGB1sfKrDd0j8PCHzHcmloM7qTl8ZRRWpwhnskzXDq+jCGFQKiOefQa9/3t2AgEiCSTtSijmDeL
U66cSkrms7ZQtlKCiJVu2j0cwKZ4FwSXm5/O/6XwCUenKly2kKta6r8OaK8LEcB/3k4UTCy39HBR
ogpSLouMrLQLzYsbCUpzW2Lq2vwcQBabqMrvi+7npekT4BIt0B4RIUjdl6K0oh7xnDB417eHf2hm
rR0wu4358ASd315RugHPN5DA0dAcKIhBi1fqqSdMHFrlrVQZWw4NyMuRAf98vGSYCZRbk4lA4tXI
ovhJAX9ZWc1ta1Xrf5lwGszpTV8MC8LfVV5as6m+ZTFyl63MmQE8eIwu2ZrN3scEXhJtgE7E5YP3
exSOEpA+EKqRsrQaEiP2spvZ68EKe7CyzGrjm6DDZ0iPHiQU/3xRonH41PWJBi0K0DQ9xDDVnxED
kSGW04vdS7qi/04AHFw3GnBQBznGYGM2xp3RP7wXp8Z2bnLf14JsJSXL7ODRyMlZjjuKIIn+4JdF
ICkQZ1JGqoXx3LpKOYlTCSsdeHD/3va/ox3iejfZ4kz8j9244YOxK2rmjQe7Uaa4zQiBIfO4OHJ7
EGve+BBoJvRYZ2u1oJU1YT9VPVycUTaakVxqkCe78rsO0jCBemgH9ZOpzB0Yda8RqkwmRUFT1r92
RBURJBGV34rhVHGjBg95uvtjE1kJf3o4Rv1MdPUVmifZXhRmd7gijzCMer+Z9qKsaD0TKNI14buL
WR8fNoM0G6a1YCenoUZG99lCpaTyrSsEpvVfaQqT3cHzie7ROMJgHq34ZkYhXNF2U9Il2spj7mCu
2BaBk/HfvYWT5t534Vh3PgAfwbWsPK5rtFoYjT5TEDJ5zLyXOW+UGYFfcvw51Swz9Siz/aQW3V/k
yBytOO0Ci4CZZ8DHttOZuHrCxPFBS6G3hqtDirtb5jBrP2j/TQhdJjAHxoBVNzHt0aiu7/VNvkhD
NXtHjUS9K26s84kzt2W2J4MjqAz5o/p1BY1xNdLFKyQXHe1lkdIvVmy3miZiHiJljzmfuUHYi+ae
BAWSzp6ZbGJvw5l2wRNBALu7dlq3O155afn5sRS56uUCD1A0Kc//Y7m21qZBH5cAydH+lMo//w5x
6JptrRduzD2vFVn69vef3ldoDj3lEMXrSEW3mJK13CGbK64ryuppfbxKOacTHgfb5Zo6oaJBmXta
mbWA+w5XBMipj5IbmWutR6+0TitfJYr+kO/vxauIzbfPbtKhWPjG9vISlUsDbkJAGtpqxf9Cpkjs
hfWkqohhRwuIBokhl2dYDUR1ya4iEzAxSjXGdMQIhm/5gDmuvnLdYa6zcLFn1D9mdzrZw9BSPOJ7
imy66h272Q1m3L0QMVhgApDGLFKi7LdWsjfBhBe5T53mBfa4FDulSesmjFMwHDdFFUsK6eYrLoAc
1VlcxPerHechf+1v+O2t7aEJb9IqTSjPm0dSivVUEBn0oD5qEEQlqiCPCjN0A9AGpZo2U++9Ajra
yyT1N9DR1N9fwB330JedDgRZ3i4KZnnadHzlCMKjNb4ze8ox+6nRcjgJnSYLulYBG7g++XojwbR7
VayNAUpxIIJZudA8BL31e3sr2oqMHdEKCHSGAWc7bXOvuu3E3AW7S2KJfLuDdlHCeugR6pOiajFH
5lwQDCLJ5naO4wv+xe1G8YipC7ivPEVzKF2GHRQ1aXlri+nex/hJ3O8Fv7ik46AZtYkgxHJ7PsPy
0/FS4l/Nzx7SDzurj4s+Da9UNXo4N4MiUHMrTq0EiTWiY2WetplhsT8dRBNRuw4vZ5gFTeZkbE12
0T25dhb1xt7hVZtsIc5Pcjyg0gXZ6Io4CGfOaJtIus9H2Gd+MlHb+ecKii2HehB5DbCnym5z8frm
T3oBjGeWM5gXBKkSviBh8FHk1pqQJo6zhMDhO67UMLxz5Toh/fwdpGaNDNfFYOwvJgIuRj/DmIGc
ceib5hkwzbX9tkC0nB9FQVfPKoxG4s6P28JLfCnP+bdfGpuKxiILYUU1v7pcbGHhg81opFdNk0g9
rgTnuJXYulRorJ7x6OTGo5MZIfpYBWzePkfM+fwP4Kae0nMBx2T0Q3nAHivBx/74cEYTi64WvfZF
gopHwgIMlFo0/8kSewHyWn3Y3Xp0Zhuwr56kkEZW0VwSte7IHk8CqqAjxg1KJcR6Mj2YWRiJ2Gus
8ZyvlkjBNFga/SSbYoS10UeavTHi5hPl7spV9EAeWFZG+wjsbcnsqh4KSsg4qc6t0CQ8pi6q9WsB
W+/Q+vTuc9hpS7cZGoT9jGaEikJE8udcR4wjUs8klbdpHoNmpibhPvdzIN4mGzeNYAJSDzMAWCB9
wIvynW6hQkiRuOeIjqUvRhvpl/HS1l6TxdplOEDsFirOA3VRzfTAOd5XJdHhxKBT7IjumQCNcf/U
KYiHgth+nZjZbLXql6DkoPFaPbH2qD7Y8d3T3VoiV48fEqCSb5K2tM4vgS6SVdx5WtA28sSUU+LE
EEwP2u155XlCqVLhtcWvwwRIlxSn5xSpdabOXSW+abhKk+wHm+ZYt/3u0/0ts44sh3gK1hqN/NmK
jwNq4rrEOAcvYGsFK+AwxIk4z9qVdqXhxf6aB1eDNwETnU7zSqzvNe6VEOFq7JIqKbm9T6F9t/3U
a5QfKkz/CYCLpqRZ60ibVjZB/wwlzEC/6kjhLluuTCdboML8Qv+s6AaUBZpUgp3c6sBNt7/ZfQg0
izBRX0VX7jg47tLI6R7ATNafXr6Kg9K1Row1oxukJglbKBPXQWHehWQMiACj2JSTzcwaUwlQE9yL
CxjUQMvokoZMcJgoGnZgpmPKdLM86ltRZ2r8N+zXd8yZfxN4OL4RL7CbvYptpGE6GpGqzq4dyVa3
ia+noUPMXHv/YaGI/TbcVW1gWQgLIu03KYBcWbHuYDbkold1DS4nu1wRaqShbkOjRt/rFjQrjl+I
8RL0q6dq57RO+Vgv5iZIn/5ac1WxwAspupcnYbGMljR7fNVsWS5IKQUF+fd07fnTGQ4y0TEztWvk
V/qfTTjrl3gcX/XMcUdZXkKpnMNbnOaKZc0tIxWpvkdjotZTC/A0ksOVmR+IVsHCZSf74IxVPEZl
kJwin2UugvuyayaJ25r8rvF8TQEbwgc6FkUF9j36wYR5hZui4yL2eghxBC1tyuRKIkRYOmLzDwv0
FUFoZLvsA+JQTWaX42BDgvJJv7EX2/wQ4Lta4bZoDqm1aB2NeCfaD4lcuTDG9EdMMhR6jIwA4xRb
/aZO7666S3SKL95OyFFJs9ZVxl8OPEIYc59B1Dumu3eWHo19qk3l5Pk6xvB4HwJODhjjRUCRNp4l
S7qt6lZfTiyiw/LRfVQyNcfxhM96yU38yhBReCCyUeOENKCb+V21EJ0hJntSGDMLYHfHdMKNcMZT
yAvKDXEaQxYEabSbKegd5CHwNZCB7aOqrEus9e1pnX88fqKf8nGQJuVoxCytO2/ubmSSFYrGJJtl
qOpYo+vDVXweN2vIeOZdZsM8JFSMUkoOodHAh/7dsek8b02i6uoYSBhA0ZsoiBqpqpjjUosyfSjw
hvqXJ/35IJwkQCeKLEoRv73kNlTsz72+izBFFT9fyXD8ZQ4SwvxylNqjF3QiGcTE6fKrHnz1eF2P
76RRjjw1K1tA/3j4oIaVPMhXeMQmJLpQf6uKWnRArhz3xWLFynEF0zu0+LF0/5dCNdv9msKxuAB7
1mMk298D39hgBipMiEM54+j28q8uVsy7iCciSi4ko8IIBVBmJpQ4yRmA17tjAeNS5TnwdH/P64G5
QWWJU7mEq0C6MPWwU3fW5EYn6dhQQA6y8VOwsAEDJCSeuJZaHzlgEqsuegIHfyiiB+Rive4bn58v
HLhlscA/pFAmk/p5YdBXwdoeM/c1ipY6sGjzWq5aeCrbYrYXo94AI7Z4GPwgKKc1fS9+C3Jas7LF
6AzcqXhxk1KVsj7deYXX56Ikzs+4pDEfL/AOdBPoomohI1bOb4unT689fk+z2fVrMGI94TKU/4Yt
DrYOjMxWuhEhAvwWFwcBabJFWr8/rUdBJzKHHoLZenKBUpNvrSgKOZ7xkcfxqIeEAcYDP/aibIri
vxgiN1495UPWVT+ya9M3SXCSPFmKLBVa4PgwQiUghUUwJBy5sON5trjuICX7VF5GCpGjQAwF2W+f
zkQcFx4SMsFzd9LUplnUbLrztsa8Ys64YC7p882aXfUtZ8PsGfSyMtyEgUiJeG3tLRoV1WtXS0T5
8HkkW8iHD1c0hccmxxB4Hh/vRTWb0NFnJGbQNEsmx7TNMa4OBWSnZJe5bBBSbgAGC4fcqQU5fmdc
3xwgtuFI3q+BlfCzbHVGrgHErLJIFBPbis8qb0bjoRNgynWR7TqrwmIGkHpdp4CMWo7AlSbwwwSq
B4wgWHpXQJ2oP6H007mbr026ozDfSXNtwa1Wjzbm94l6Pg9AZaUgqXS+O6BDbNgWO/Y9Q22OVK4V
Z/sEgIoNnjiJmBl87LkFrach0KaUFPezkS9EN+EwSQKXBrZUEHZJs/VOkeInSL8Owl9csMHGcnn1
5dBEY38YbJaGBP3RXTbrju0uslTyCcbtxO8kX+5ULLXxoTTIknaXeEKXqpp2G33igePJwJox3l1b
YF0CApzfoNGUrWM2RzRHuqW+howOBAVYKQXWWnZONYRDDzYeqgm93kVHYWdVOYe0KvH65hbdAn8r
65mr+BG2dL/e77xUf8LdykzEoaEOX4WI57XTrzgfcC4WYCFrUtw9+Jqos9XUyL6QHuXM5jErUfpd
eO9A9TK2dGFACQ6vPBfprY/B7ucwOZVd7Fthf7VwEKVS0vELnwpaJq8J1b3rk2/wgz/8Ev52cyxy
Otcy7Svg8be9hdgbJIorrV3PMX881tOvDT5Hu02hFAht7oqbcSdnS5NKjYCbLcmHeJOlx4160qrc
331qwUqwnK+1S9Ri9BSTzCPGMbtYx5dLKsHuThyioy/C3H9map6E1ERmr7Msz0uEAXuX9/8bQy+5
5IFNF5bv+7XFzh8fAe1djMiDjtSWeFE/khPoenEySe6mfdg0Rm3vKnu64yn/CnHkl/RafMGik1GQ
gnG0ehPocwtn2IMpwXLhvMghEYYcNKH5VQz29zF/hCh3D6stFye0zoS1aO8SCP4FGPfhx+69+EGb
vrJqKZ2hQcImeJEU34kYQc1cn24OHRObNVEdIQftNsjesEBtdZNxBCVwLbOhY2FWDjj/Y/hZRD90
PoXKGN2Nnfl3di7y57bEbtvb9I3KLGRSYZkPLcoaCxFPBUiqhVPZb+ZBgVoJRzPIjHIbU69NuImO
1rrS0S4rLDPhlixz+l0eokoQrUPXos4UHcfO29m6x9MZcEgB+dBpkCOezh0whUUTsfrGk1wqupdu
tsZdJdgD7gQ4GpXPUpUNlREISvKu7nkrw9kZVDKc6eCrmeCDD6nzQdhzgmjvF3AmM9BrnhL68gdm
IfoiTUZCrMt1HyadJv7qmJJ/Ij9+piLkcUk80ZpXaMakck/4XnaWwXtRQdHPLKf4sv2QbRoYx7RY
6Gy536JF2NZpFc3jRy1eu34nJIzD7FaWfco4M6OZC1XsyDr4m9/pmu9vOjFS7FXHILDza4itmoQE
TV24t6C6H+fawVvgxGbFaqZRhHGJ0yadv01C1FFgzh4Pd6er1ZWsr7sdw/+oLLM1Sq1TVywd+Jb9
tpbLSCIWWnBWOtIHG4WUqKA78Up0nEKiwAp6tq4X/mJbFaBR6hxGABKXkQ1C2+OTm+hBASMlmIMO
EVyCdoEHISasQ/1/kUvcY6GwFOVMY2Affe6EOmi0QczVc+E/nlxnOM0uXChFQMl+H0ZIc/xIiD9V
xfHV37BmDgk+tL2Pan4xLjzR6I0psc3CCSvMkeCEnbn8WyU8hWBaeOuCWdYIKiY6pVvf+qLVAPBt
W9XW5BkpFIrLCHgE09BnAUI2QOXAEiNS1P5BHKbSAVvcR+I1r0S2idUT0CiRbMM7hqjFiiQm1GLN
Iknlby2t2s347uuFLxLj3rombFAOXpBAvUp1aw/bTDlpdLnf4EPbTKBjoo7qObgXtELAllQDs0lU
4DhUkVk69azzlZkbFaDMISRzneFScJXq/j40TwdcAmxeXUyfGpjgqACPX1CU+GF1seiVhFKno0+c
5izESCpIuOcAOJfo3iS7npzsgT/mcCdQr2wnjI7RsrgXeK70ukSU0n+0kLWWzAAVaCX7PFLSdknX
DnsaWQKNAsxjDOtlFCwmimeeAGeikAEMzM5lDsyopmmAyDhuPKBrHzDmlXe7PWMqumSUJ4EljaHt
0q+WSrSmVZBl3japslvY37XNVidipZ/DJ+a2IQl0AS9fCfqycwPjJAH0pviHm2JoujUHIldoEXLy
8BVensr0PEAYOerJIAalJASr8allenvPpf65PEsGkDbqCcyAlm+VTokDBvP7t+VgUPp8IjyjlaeZ
1CbW/rzaxgQuct7pxstl7BXs85gGc9ZwuB1Mbe2qbxZMqwE/U+2YzYi+fex2oqlYER758KPNCY93
dCAbY4p0FAZS6kfSkbNK39RnjIdxbkg9N1z3f9n0bEQqwCOn1cRAFA8sRccY+9CJznjryPqYiH4O
GXV2NtjtNp1ZUxMXvp8+BS3dNxuU5XyqB1n4hh63So1YRbvFfGL2YHFFPbh2vCdkTtfH2B9j+dCP
RcxLlPgRRYOnFG7WGHMH3Cj+C5AQrtdBpD4rNajYAcTnhSRn427Ynl6pjbRm+gxxdhssc/S482FM
JdSVvn6E8UBt4vIesgFH3gvjtD4rz/dWRFC9dPyyPKwbxptnMADNlBTJOG919o34JgyX1OtT35bx
GH3VIOA2Eo3PvknEDeN+dg5UJ3eYDEj8G3dnDusPhSITxaaLT5vZDka/fRp4ns3j/hidBUyr0jzv
aJDYvAZba0M6gJaV61xy3Hb+lEwcZP0dQmbpZ7CpEz/nCptHf+w8PYyzbG2NHn7F8B2GaGNfB0BI
jlL/ewMK4kFgvvrpe+KAkxlRQGqL6o6gSYOjU4lGbBS/NVjMX4d2wxkj7o2ZE64VQGaU2MpEVTsD
QcED4qqKCR7p80b4aMwubGGhgbvCl9y4byRR+F55I9Xj4bfo+RBbH+I/eZJiVhz6WusKQT0y5Dsf
v6M+tRWJcvFWnV2oylyFMAeMomcJQEtjDVs6nFLed0lOkVb3IIUddrpvf68cjf+CINt1btgZmAzV
9nlI/nHLfqKK/R6Y457e6yCs/3fI0PHC8auEe0sO0J+TPVdCBGWbDpEMRgm3jrZBrs/7Gq/JXEcu
yf0/bnPPmCE1iVZMfRpcuP26HzkZiEvfnPgYr8ZJQgv3NYFr31UbhETszpocwfxtcKHG6z0J4JAu
Xq2sOisnYi13eK0hBjmFLNsd3vZYzKYznykFpli5H0Htm4t0XaWnAJiOI3Bu5XelW5rn6jqYqDhC
MkshwX/sHy3pQGYdtDJzHmus/Q7d8yjAHrPq6oUQqsbE3BVwmkM1eQEZuT+sNJjfJyUDvfpKEBA4
ya9lyYXZHvGUtpB0AL4ASDPlHlpX9iSrJ4il+xz79HNlEVNxp20PzLKxWk9H2njvvEJYPukLjk1u
Aw/Ats37em+pMOGK23yNm2OUToz49z6bBfgMOtn6uXZpMWU5RBpomjfU4d1OnMkYDyU1mHVvrZ2a
YuZ8GmvEjz8ebLQIP1dechiiJH7LmbIN0U9JSlyG26CD41PDr8Sci4QMcnuZ0E11oxUhjb6T4wCI
OYUojBjLfs5nDeNVyxczEsA+vBPanzby1BoqMvOfcQUNyB3cUewv3fz5gx1Oj0mihJup72NfPUHF
eJuv52/HIVKASdKf3tH5gW8um2fuDslRZYVdJFfg9Y44ox/wglrNkSCFBY3A0g55mP83yqY7v6UY
1pqzIBRHwI0Ng7vXamCUjgpPIhx/ngkc7HMHyMGBTmkfRAYOif47n8I+GS1eOG6oygnfY+bccZYV
3FCG0j6fWjLpHJjy0pnO29s8R7UkAUtncXS7uu2PqjS5/jTRITY7ev4ANBmX9Xz22MtruYl7MU44
NDzRZo5nD4V3hYfj1jC8TPRr8h5ZVDIwM8sDUJ1FDWz1Vk+vybjFjFTGWeZ6uQTrisqLsh5izytq
F31gH6wIeimB9OgyhJHOWG1Yz4rPEBAEuN1CYKWup9QHHjrJ14aWLaAqKzTnSJzMW/6Q3hfvqv0/
GCZ9qsdZBtHQj83jgIX4pXfM6kK9VMiz7aZwbM+b51p7iKC0DCcuSodYxPhA9uRQ5tWt31nPJ2Vd
bVF7Y46VKd/14DwazghBxJoLeS9tnmK2oVn63Wa14PtHmDk04pdK8fPYIZzWyyr+iF8fvVnzhJwC
bj26pEj1s5bfhlFSbfb7F/j+RkHbk7clglBbaVQ6f/sR64Km++w4k/2cyyR+tvWe933JE1Ln1kY7
uOvjNnYXVNKV9jknwlB4kMTTJ3ZEw3EKLNbfOjHnjLxmFWpq7FW5MdAi5Be6ZNjpIo50iKkXkyy4
OIjlPfCOL07e/BUE+AU0DdaQ9vS/0X2JHqcw0ienvlz7UwsyeCSB+ILcI2A0hsES00YY3a3T08ud
oeobbGObOAZZq6ycGpDKEEWgFzdhHyf6mBtOxX9maSn9Npex3yjIdveZTcEZiAFwk2mq2r6L0FKq
qr2VgZdGGAM47CygrpL7KXdx09YPwtIMQOtuaxhqUYsKLRcHtT2RJ6JPGnbFDW/GpVpnZT+CMTQA
AJ1Fo/wbZCJ1uJ7KocayngS35B/4I4ydusECWbShslVrocO9iIHQ/JjQevu0x30Q+10GZWIfoRJJ
f0W5eiEvhdUB4Cki//PsfYWQsc7CKXqxfmhUQDKBsAq1godIUI+9OnMkeK6vnr1AoMsrM1hAtcCw
ik8hhiaxzKgU4TezTFV1IxQzCTKrce51lmYS9sChsx7A+HMzoFrK7YTBY8ZFbqLt4T470tZtVXVR
BUYGtNNK1vWKmtpodPb9FQQiZfYnveoODXdJqmghl8m9GQioKkMKOg7plSs6E7m/TEyCdGFmJgze
H+7cXQI7q2LMHtlny2eu/bJTn1M1pkxX21OIx66O5azXPRRkE6NTaABwxkBxTIkxdbdcnR2oqEqF
oiGkUJlO5dkq6jewALDZV+NQVkBdFrUQw6xBoFjY6BLhi/YZRVEGNlSrqZWjD0NNuzAIPZ3LcKpM
zi3g8ahS+6ulWmxKFsQVTWZuCqKrIxM+C3VWEKriVfUhSPJT0/GbWnKQOV16XS2r5TBEcfjVJuGY
EHiIRRKtBVbQwCekf8rvMPBl9unY+5OYd6iV/UmTdovn6MCB0bHGxw+fZzczQIegRMSJi2iORFIO
C+VM9OwAfvaFXIsB8neSywUvLAHS9Z3JraqPIwdVxOT7tQLpSI9vfDAYVq5y2Bbi20bXrPC8rnqt
lTXy303MT7s44H404tZgnYycNtzdrVogrmXqnJ0BBfWbj+CNTHvfd//SAcCIUaxfDjI1mv5xqRR0
WQBJIbVHQxpLINVXQDYNbFnK1yLxIQ7q8yWsQ5USmuWJPJY3pierYxtAfJFzQpyhutbmM4OMJEf4
vkARrf9cN/eFu6j9Y+4m0AM1XIu65OVwplJ0fqUGW+qKXcgISEs8MNzZviRV/z8n9+jLmbf1RAvK
VRLbrAiLlsZo8Od14Uu3SLVZeniLjHbYBV/kshh0Knn9YHgvIugJob4tVY8FcfGlLknqPQlThdGp
gZg08oMK0UOXxWHs2xqVFgp7H58nPvFRyYoMsqFvksOlex6Wgfnl2XpTFudmXRX7qyLwHJo0kMP3
4Aw1/IwoO25TgIZC/VDm3vzUAwFXj4lbYblJWsvBy2OnxujR44N269s0ABx43SsF/YVbkkXs0UBa
VB8+Nw9RqpoejSPE8QWMTW+cs8m08weX1x+LazATBmnpn9qyoWdX+hVlz+vyMd1BGS7yreywta+Y
aUxri20dfnklugLKe+csNnXVLqqQEoGSiNALanIPvlhRSnE3w3g4bvDNVG/VXS+avW2P5w9alJw/
1Ts88bkGAbCsX3gu5l4qNBou1MUuXRu12LvZY/22lKx9JZN76eYAcACKT7bNvfLe1qy6c1KAy3Np
1QIAaCJv30OL8borCMFricqsQcSBCdPiTF7JAzYT65kuHMhZip1Sa8YlDWvF51Cd/nTqCbuGSvyC
r5vUXoeWT38rKUHPTsFSgFBUcIp/udwzebVjPSCDb2z6r3YRe58kblQkL1lYdu7Tn1QLlClOshPX
hb6pX9fAz18bqeJpnRTU3LH+ORBZbBzCr7z0SHxmUX5Iix9+ZAITTk4XysAFM9wQ6fPTocRNVEDI
a7mUzDTfLUhLAUFP61cZxgUr5zendVHX+42za65u4mHJn5MYF1cM206y+hBj4UBgt+/VEH4xQjvj
CI8NGGU4hYfA7bVbJkA6YlTjPKUP2SG5UUo2Es6pK369ITl8HfCe0hXLeI96haLpDY6YJZwzzQ+C
9fAEIiKABKRAj6+dgVio6XOKcn9EWIkiIB1nwiNeZoi7zFHm6Yo1U1L97iCwAA/2fUK9k+J4imIq
41Fllhmqh8MTxVLTm/pHX2HQwPE7ECJzs15jVbQD6qFt76Uhvt+skGdzwA05XZXFNHNtWq8ZRKoK
x4kz1400QRWjsyQ8qsozALznWJyJMyV2r61DyepWZ904HAbXS31CVUX4F8Ti6ixOlQfejTKrAGxK
wbcnf75LLrCSi8gXlW20/xcjD377ro7V4Wzdu5RridneY6qryh904RV3ualp5x4HoDt98BqhTObe
28ki4vIz+//+Jj8NWVP+mJTDnN59ZBlbgnJsU0mOLbzQfNIUk4ACkEoRl40jlgMhYG0YkCG8Xpe+
wDtkJHZj+lrYcw54odEFt3B2Fn0X6J2zpcSd72rkfUnAutxT5ibGfVgXUgwQS4DQDyM4GYJjCAEM
QTn+yEg8/52I0Q9fPbWjMIFd9L8VFX1X2FtVK2kriE48wX0KjeVniywRphSRNZWjpTx5U6HvgGMT
wfHzHGK31ekieEWx/K5IPTL9dmKUhUQGBQfjAuFbddISXiytZgvbkcUaUBPZu+L4LPIy9Py9vXop
nEFI+chUy8U6jut4D9jfbYypEj5ZWo72RrSSDfGhdCBOwRfap1SjyZwn8tsKQzUxqBEeAXyZGPkm
jtQrNLXhYKB3QBtqgP3i6QGg0U3APR9CT9OHXgDs049DTIzEUPOdZoe+BCpzeCg4yLrjfvtts5as
23L7ChZcw0xy95vcTv+ie/uzFN2OaxumohRcF1wltqwM9MlyJFROYj1kEsrUn9ZxJPPha65Us11o
yiHcgSX8syTLXYpGuq2/ZGh4NR8ZiWeK48JCjbL/x7BhMr2HqBM45RTmROpJ09Q0YxqcBLYdcu3l
eGsZFO5HOL66DCWdDjWTKDiaIum2qsIvKc9/+KPDpT3r7Pah5xgjRMC4QCgpxodm6bewQoQ6gTyt
kl3t8Rm03viKWBfPxYGbvsl0CEGZ9egD1W3lrmFyVIehdoXoN8IQegnVygE3qG8yQP9QWtXIsapp
oapW1TZqrfyK/W7ipcovQ36TQGjrzLOmWrNk9uJDMK0jZ1RYb6YCO1ZC0MpxYCG7lfPIY3ua4yOZ
2PZsYELkGh2Xl4WLT6PBanQ2cL85nMig3OayyR/opM3DYYvBIJ+HGoGzlldE/mTyAb56N0N08m1v
toNDpZl8Cl8z2EsEjADn8z4jy1xdV/GJLumWW6cvhCYVj7OIRNyjne/D7KacrKElMJwqF6vDEqSr
3IbsutX5siaYPEWfvxiZS5uA3E1k/HGaAsaXovuleC24iCwl3Ldr4oyeGqDeGhRD18EIgSMzeNdg
4JIobesYaBo8bueuImAqti/++5GKBNQiIgXaXs/7nrKpjlEi+hYUDPrWdbvmxGCPmInSpqbhshVt
6A14s4T1zmC+4azZag9G9KYzFkDgEAs2ohJZE03NhR0Y6jbLXLaZZb0pqgw+pspb1CSGrI/Szlad
TPOI7847f6fbtvNxFCz8ec7b3/0zOW3b4U5Yxo35AS99JWcn52g0i5sk3Q5TCIR6goMbXhsy+ztu
2En4SFHfUEtuh9WDWhlAtbyU9O+abwfUvykiOtfLok9z5X8ceHg6UnEELMRQmK9oOIffz0dgUKFE
nRPxtnEMOQ2M53Bp16ANUzfA21V9A1yqf3hb0oVpbTuKRKrcRBNPBP7L6T30ubyJ7myNkgU5m7Q5
ioW/xTJF1wEPqqy4/fe8aXNcyVaHaAAMK3zPGWwluOm+t6AvtAI7a9H01+KtwlmQtZXOjwT63u0q
KrcTnh+NFi5x4naBTiEBegplxwMuxtbTIFxBIqXQkbjcHOWVnAb44R6pC6NU2RQIEO/UBYufNblb
1yc9wYuzDzez5PtU2x1VLX4PJTsAFtNIuxraJawXrZhqjFeAmtPO2oiS5euHVbJcNEG1l7ElUWIF
v1tdx3BHV/lHGfS5imhk1kmTwLCspsDX1cL7x0z8KM5lzpi51c9YLTaq3KTWZIVj3sTqJW8GAqq1
wQcdJnbYwkgPtx4C4S09itISNpmZp5EfKPgsFeyzwOCiNQXy8uYKJ24qY3pZyM7mXKwl8m1ppxBW
ZEH2RVeDosnIsBBegUbDX8/8amycByn95rFTJHR1+4A44y/B0ilJfIIMEHIxfHpVHnuaPNlGLLWM
KCWatES6gTRvoxujXb+RojMhtvVf5yaGoVqx03ygpc5mJoN3ObTaLmCQgva9fiRv9jEYVc6vizgO
fcMBzACYLg1opMzuM0/K4vWjWVFYPnO7lU9bff3O8oJcnGmLxocm54KAv4k4xgigFdLZhlLQ+mFl
uVLV0+P3EYS/Ov2kgwtO0tn8AT3i0yat7rikeDEgwHBoEzFfDDWWsNPtz6bgmVtg11iyEWt61i4w
3t6WIGcFb13YH5SBf7y5oXH1xXbBSFCFNbWalxqQnIoV702uH1sMXrnoRmZ7ID3lZtl9jv4cFzQ7
ToQnWsuidaalBAtjkttWKjEsoT6nLLRwgr6VYZeMbrOLc2+NugdrcUbFZaFNW5q4izh4BhaNcncw
uER+U3cirqVPypnreTno2b2QL1dCG1g6K2qlqo8msRYjL4c30kZ4hsah7gHZIOSG88I5t122EnxN
z1qlc9Vgxig8yHiBQzHxsHu7kPMSbXEFxi9tKWk58LKka9t5VeeinzMC8LBHiNJEG+T4zrHeCxdc
KVdNF9hpfJ0WO3uFJNsf8l1AXvkJORUCjcYL5Vi2NFeIaSvRj729RguXzu7WA2gb1JS2nn34T/1K
Ltb9qfcLbvY86X1EI7l7CpvPQepJqbkDxq3WaSwWdm+N7KdLJwYTohNXSaxULshsRAv8kdMQYHL8
MYHZGXLBUiBCZfW3Jgzm12j2rVhnsP0X4/zMdLvdeEuEpsClXOxrly0CKf1lTauXWFbaLXd4HzdP
/ZHdWZ6y0U8WX9intuUw0YDEigOj63AjIEVVIEI/DOLKCBSJV2sxk78gMszDEWDHkUdm6XSWJJ07
mDZwVT51/fzS/xzmo4bRZB0KTQvHAaD2xleko4Yw6FUHc6KoIeuuwVp2w2/lFEXrEzh2qOL3vs7X
lnFD3ictFfoEoUiT3aYxbp7/1r6TGRcYSipFlkGEcz3IIal624coXycy2gOLccMP4tnkMUg9iIyZ
BaycTMxncgtmAUcxBbZTYZHIPNH6oVTeL40Y46U4c+IMKzqc3v9R+cYRaUExqDmAzxXgKu9yHJ3l
ZHomMGJdGZQUBGf5KXc+qJvn/OGIo/c3FdGZ9Fxab15G0Hsi3P45nsTM01U60Ydbs2zUWewI4fwB
GFUkJjlQw7TTlryUOD9triJxNsgx5KUhYotWZw6gNAyQr6bN36eFuiGexiIv9Yfmc8Q/bxg4k70/
q/5Ks4Qki7iSFb9188l2Qp0IJ4JukfNclQyQMyIwn7LW/89z1FzpfRLa6/3+3xPRmZfDnnYRF2Ta
/iyZPYW9yi5wtnfl+mDtcFdZ60sC0L4SjhsKM8Mgmqmz7h5WvQ7FR3FrKL5GP1FO313LxD7FhjHV
ua1mQKfxZM8PZZ1jX8TJlY+O6941/N66xeH/9j+0qMmGTwaZ1ITh5YJODktOyZdAXdp3qJF4le64
YZB2Xs3GqIsyP90kPh7W8HL/qVjnKzNAT6xLLOgO4b9Twgq77B/XrTGmuxrXMJw1D9Yj3oiHf7wl
6OMtM+Yxzt1H9+ZH/X77gnD7C6A8IJl9eP+EQND3gx4jgaFgPbj3Tob3TubXLrbsZdaE9RH8oFIk
yF82F5NEDjO1/+xePDQokDc8qf6k4a5Mt5vLeeWj/6AoWHxfyB/tfIQvxxX6cBKe9RBK48gN8A0Y
zg72mGnAn18ro79GY7dAh4BZ6JCY1vMHW5qOZmx9ldVPIovdIlXjU4hgY+yjdow7sF1rcLzni/v8
wnYqUBB4cfEslh8xTYnjXelcXC1vKYsZQZFzse8FlGDZk3ioV9I1zzTNBGaDNRK7bleRuQLU3EuC
InnFTOBR7ynHeXmqkRarfCCMWCgGrmROlv5drioA/uylOf3XtLHwIcJUg6+4B9PsRoMPmaqvd6QK
AvSWwB7fyOkBPSXWEWY4Hs1Y6Px0bPddWbWsFgzBOn/ewB8KocC2WXG26DcsgoSL0ZfkHWJhejX+
WObNTnUNnQN7MEdcHpT3mOCW7DIhTRj9NsRkSG87VcxdKszwgotIgbUCAHFrbDRxhJWSduo++Rrf
/s/ogdnAqJSlxyOP+mvx8viDdvfN6gQMbMisblG8bT4e26yiUqNVqnDJ6z4r9DsAaJ/YrPg+mxrQ
HgkEr9Krc1LUEMFH1A7umbcOOADiSXmXTenHdE5NrxciPxNpl4XNUVi/U3lnlzxA9z7EoLdyX2t2
4zsntwxQ2m3cny1fEflleHsUu+KavwhjlgsFA4VHBUHJqGtpvSggGev6Ln5r5AOWcCh99zYqB2O2
wh/n/S91WGVbLvmEpXGo9ypL4pB/VUx9tTofib+NaabVyGHu2iebY1FOAPd8vQhz4X4JgmtRG1Ey
2u4lGQU9jkmexQlVUgmHCbgfcZ73KuMMHPJWg/lhST6RQNP6+Trq4FkTlKNJgju5SbWH0WiBjb2v
HWFPuIyfTDLiKP3Ttpf9xTpWoqMax0/+7/7LewpjiyjLiK2AJcvlcp7XMe3amaWY5SysdJw5Jg0y
x9IsqbOctrnx8tDaRXftVDB12yWdvTf9xVerqA8/IMEwC+C0TIURlNNaBmCNm0WYiOBPwrLH41EN
i0LnB0anuZinP3UYyYAoZPa2jPzOtqW+k/sZrWH8OxoE/WbVkCfafNLLLNkI/sjQhOcvEpr7yY6I
3Nj7PxihiJz6a0XlMOFih05ZKay09+b4Hddh4UJICXJfZP61HX3ogFFGQZDpcHISQlJP+T4fxo7Q
K4Bz/hQw5oF8kr9m1RzVlxONGK/jFIQhNXHybsFNgkoTMkbU0xs5D3Kih+8ut4Nj5Is7B4NaOzs8
BrqOOWg5htkBvj7dX9HdRLY4x8a3WDEPF4YBAxjHR1IAPOFKO2f3XfN8R8UQEaAmfNQHIpxZ9S2q
p6vj/cd43nDvUwh7/Gf6UaDpvSvX+JxAOhFoFUsFgLUnt9LIE7aowVEdRYD1Cgi7oFk53VxuxBGQ
y/ljLfw8bFWk3gqwkDkmDwsWQepNIa1IMHIA3t9OQplrFMYlYz75mudYqYI47w7wDNiHGHD0kXCm
Ynrp/JvG3FxsIihIBwTxKEbWgH88Cj0bbwHuPDEmFF8BPhuzluRBlCow4DdxZ/clEhohnAhysWBd
ELTgjq+P0ohyzn2yDleMVBC6nVVEEZIvJbj40frmZ0L2VIPnAHKPTVg8JR0lbyfnUVbBCmINdssA
+P6nsUh3DUA5bb6U4j9DDhZiYJzjLZOeung0vCLDDjSLW4jJqvq3rmkrdMU++PQz49CvF7vb0cic
DMY8RFq2ilWi78MiwEzmeuCMFu0hu1gNqngCTtyUygzGcVAnpHu3vjXiRWeRG+PmTqOfiSeixcR9
cBy8uVC1QkcZix7uZi5izBm0YSEZiDe2Gu7B3lquoLDfy8R5xAjNX1uAT3b4xEKEewD8DWoroOMd
Ay8Omw1+MSiU9frwoTO0sV4UC6sXH3uWQpROI4WS0C+DKmX8/DoDL27tkqEpD/VJ7EqpZ0S5iVFd
XBLYEAfnFZp9hW0YrMAdkzlu79RLzSyFO+eVlHshJ2IhEYw927kxd9jAvZoVSpwInbc1qTqtSr1/
PM8QsTmleQVocwHElPWZSD+x9fiWTUj9ikJurQoYmgdu82OrBiknCFWgiIHuF/kFnModfRxjyfWZ
7+1YVP0s43H2WCwnf5G14GVFJVzcFbL+QJBUTxtYb/8z1zfNXsZR1V4iVtwEY4Dz348MEJTIZTbT
HFeuAiTXC0ajA69I5fOQ4iZoLw+3VxOLIQM9/IHhFfJa07VS/iIuadq237z+hfO14N8ePTjfNi8E
ciLJxAlMHfi1ieEWpDmS5u/XwUzJA87w5/ffMYu4ewzbasmPVX7HuH9M/APE9gMxjPnnXn3fm3Tr
putVN/w3PJmsCzT61uWgePW2B3xA/HgXE4EUcBGOGsgJI9fU/RdYfujFKKPrX1uI1p3s3sO/jagb
Uzw+nCMy0Mo9I9/VI7pke0UxIXthxy1fX+2vm7iNW0rozehsm7XuMeplVd+11O6d8GMt9Ev0tWNl
NqNIOGuR+JgL0BxWlE7f6QY6yZoRrZ436tYYlJ0LBcZpJy3SfRvUo9k6QqJtnvvCjeargYFOnZ8T
VUcNyie1LenS1PFib6q151FvX6g782werBgCL355PJuog5tfB8ZLF22c1gOGML/+zpPF++EtFNoz
jxcImSrifQq03onCFNSPlAhG1KABG9vKN3Lh+7U/1K18RZmSbAlPgkgy0UIgCJ5bAaitdV6vu4Bg
Kk5hDV1pKN1C1fIHH+jv7UUT7ykluFB6ln/Gx4SompO2HRtxwE4014X7h/VWvfVglBH1sistIy90
xg3b6zcWUDhH0uXKHB0dR28+HhtqAq+00Wt3W2xnBNROTF0bU2M7cAcAaDSxDp6KL8fNqjEeM+hZ
ZcGM0pN3IKu6RUri6A0oyeUw+2JWZ3JCE5XqGGofpv2JS5MpUpTLhx9d5gfXl1nF6DACtQ0OlxfK
chnByWp1GMUxCE4qdbzgCm4+BUAGE4pt8aKpyINnOTEdqJ2b1GNl0AENz/6t/msd/IkzuwqaeIvp
t6GNez2k3CowNg06E0tDh/PlE+ih1BYNcVtVRvJGaiQszk+9fO4GKuxSX4yzdkTIzZXBUMRIzNah
Ux48pKk4VFzw8c/Q1h+e98TAgczL205VnPow6ZduhE4Nk+xfvjg4DrnRJH73RIdTGE4CL1EsW8X9
POVPeZqkCKCluMzTEYZPk9uECtU1crQN4XVKRB/GapyWtki5+i3/KwWk6fsR0vcGJciT54BPtuO2
qgNAQL9c7e6Qpf3qCPRfzppIYYek560836drjhXWI9VrM95FUrFKioto5sTfKns3PsgO1TZ1Fgx6
p/dfZYRPhGRcAm1NLg6l5Qjg9Koe1CB3VUpbfSNL5ysCo0JLPueLfw/tGzVXw6n8eog7sT+IKoJF
fWN0+0lF2FQrLtryp9JalWGMhKwgEKvcm6USnaKA+BozTNhIR+vCrWYmGq57m1ht/oeltH5qtJ8o
VoUD5KUJ9gev4UrVYzw1BZaWSfrGCwF6K/i3cS1kjczqt96Qcn5ekKY0qkmt/6Z5q+Who+uOd+RI
G3ktaTK8K1SRfOIn9OUYS0U8cLjDgBS2Nc+cEaU8wGMGVOmo8Kd2houS2t8B068laGSLPc7U60MZ
3ecJTwTrQqTXQdCDAEV2imaXnQHS4pLqhajLQZxJCtZXlT8QLFuJZiOKc3efTLg1rlI6U+kOnji9
l4YvOGXyhJjX3NX/YDxzzuf0xxHZ/r/qpr7IHLYhp7F5Xsbk3W/7opfcq9hTNAD0I+Xn1j8Yz407
eHR/yxS6+ztd5AwXQG1sP6geYrYJQtpspz4nqbcMme1aitZfemFcbMsEUyEprR8mn+QWbcvkZPor
XUlTwAW0GkvwyCKY5Br26jbyLOYs2CYqgqzMYH1rA4yHsQv1qvxpOxYhBPntgjlh3a3pU/sr4RRF
qMIzs7w1bz8bwQWJNCAxYGlsJ/t2f+ayK+iyDSJARjxao2lxy5CTEO38SpVdfGSZa5ECnO5MZ+yZ
85+dlwyUfvBjJqSmwqGbl1RZR6xBod3sC8Xaj25uWcPKgzJF5j7rUHIsKJfLJRofgk27cYlQ1OLg
0g4OXmEBJWsanL6O1kgY2Maoc6bu0NdQzz6VUMZwtoCEf51gClX72I6J0l7A5RZ6njdle/O/v2v+
IEwXakKvWpCf2jqPEh4kUGHPig2C4Emp0sijDqaATXOI5oodzz0iGg297fMzcPP6rp+2L02A/QSG
1PMLYaYSg+z0c87E6sFEGyTM+rbeexndKARt0ZB8aixpcYgGd+jOLUpFe96ryCsXjUvZe4G8Ni30
3zViu4WXtJgLLhqeSLuQQhrunLNFsf5nl+Cy5CS/oGFiP0pe6DFrFmEp+nzsfV0LY76aV5L1WnsJ
OcUGG5B2rFuOAmb3smLsKk/7z7o2xL6rHHJ/KFlxS1mPTBzn1yjHm/HXYr9D1VwaAtSwDfPKqM1Q
+Gl4d/4yFfUbqxDribNcbpM7rQfSUxG0zidnw/G1ygBcmgdZHNhjpWoPwh2f6/k9yTgVdxAR+7Iy
3TX1v4op9QaLRokYRG99vWiQCkrOCIziKJeKFH0XdZuHr666Zt/OVDhxhrB5bBbilMkEIY2MDJo6
H/Y3/tNSaod3URF2UgfI2RLjD6qHK9NTligVoXBAvimCtqps9IfRY27euKIrrQQDLVOoLDx082pi
fFNKtmp8Qn6rshWqS7itLZWh4X0u8fuLT67s0yBXAhVmVarVQ9gFgvSvN3FJT33vm8ElATbru3VT
82gB1ZqJVgmhgNrayvCaWfB8zYFew0ta+1Pp3dd7D9NXQSUeGr6o/gdRkGb7oCyIJ97/jyYTGAzf
qS1CC/xIkd7xrMw+onw1wBEYcm0ORqe3mFV9EKAYtGRJ1R3GTlLS8OYrveWI2D/yYI59aurRPJdA
6nF5clNcNPUocjJqfb/ceXZvqFtWd+ra4mXpB4w01uDYKI2Jz28p7FQ7FbSswIVGF01iiF/wu0Nb
tpn0MS5TVM+RQTB+Qv2aDdJuEZS3amcaA8pWsbhLjn0mFvGz2kthFrSeg6I/CSRoiWkqzdN/xvnC
VX4minDJrydn/mfJA1+nuP8RsKHZo1ZLF8UalrQvwjFl834vqumaFFeJRrCFvRVAeEwAR6gi9ZFP
sRYadCbaKpNDtS5ivqQ250fjxGrdB0Znsor1xF3yiTTaWfnIo6jzwiq/gFXmZ5/FxDORlR6O9pMF
+ggTfuRiV86jh+5B874s5cIIAWcjgZrmMtz5mex82LkLZ3oyTtQqLENTTwaxL3W7OOp52LHh/MZV
dUP9hWnnsw5cWp+hH4yTfXOkjwv7n8fapxOqyxarxgrrFtIDfAwaJv662zFrsQAE7uU+sEn74zy3
ZsgOKG51L0whQIn1dGoGIe/FNgYYApHQEIFQCsWJ0YCLhPD/x8L+Ymrv+JkN52nagkrD4FUClwN3
N9gVxoxBs8x12JNssFtIVjh9Kq6HmPeLIKdiYxWUuPlPu22P04GyQBnK0aaktGR7cXGjgru8I6HE
IRdJ1CQQFvrHcclWVHDU7uDzaaFyWiozYcHN1zEWzlkF//MMQ3kVtlogp9PSJ7P7CB8d6xI0rjmL
TZtjTfW4Fp/BSsEr1QnmX2dsubRpaCB38OFr8k0QkMz3tImEM21TYstmtbG7cd7veDRH69jny5ra
+h6JqAMlZAZT0jEQCj+pkrHMvIlO3jBmQDPKo6iXmTNrP8NuwJ+Q6DkRSJzngoVHBxmwQtYTEY2u
w9eRfnweh53g4mv2tFKZD67Ax35hGDnvKo8vvDY4df/Cue1QWYomK1SPQAgTk+TzoULwolNeCmom
Hw+hvuHqHz/39opSA2yVCSgkZAw6Ll6GfrNDSujA9cLL58L0TNE6UEhKtvu7uzVbHLeOfRzK0bov
wxkDa5+UU4tOowJfnIeFlkWLiivvTD6ORMrgu1MDsJbMztEYBAmqX644f3p4S8pqSi5QpUpwbVHu
235rSo1cMlgTJ4WY89bFaGL5R2hOvLUlfZ4PoDpO9W45JWy88q5k54mMnpA5kGxWHVEd1LMgvU1i
u6pxJhgzS6zeFLIzbVlGI+OQbLBGwutNOW0dvbJW7lYXxUusb3dHj1LAtlYbmhJTNT44YBw1ltBy
irzm8imquTnpy2OEjyL8Ta7kmmO1rob/fyys2yF8gCgGNsssaO+QanVEu+6JqaXswjpciV/+fUNS
c6TMbLxX2p0tHKadnwdtcfMfF0ypaOrckdwy6AjCl0HA1WVSIQAn8IQQtOB2dx6Zp4aR45nrqYXa
yX1LmUxL3wIQMtvo1FoCkI1GOP9MdJV8ZhzxwZ1V7FS3DWB4Kasg8fP1Xib/u55dMvkuwE6Bd0fo
lXLtpc6ngB4yo1pRCGGlyqxoAJoX3SdBbSbqNE6FEFiD28CYecop+zkbTrdZfroiZuUUdaOyJgIJ
0zJzvXJ8X0lBY9C3AP/8hTFO0BBhHVoZKCFqNGrJZ4lbOmGiK4WxSIE8GZ1N/gaPykza2R+Km6zh
3HDxiRCkWZyuVAL7qHlOJiAMrbspxgz/M5HviG48McvzKt/D2VlEX6eubJZtvIZr7ocpYiir7bzS
2edbHBVEOTZw5DcXdLODT3gGK7NvIWvqsUdK+XN+9y8fDeyzU1JxXHTdiSqft/7y0Ns344nfnuRu
CSvTUJ3ZCwO5ZOcrQs6bMruDGBgLeB5iECyfYggdC9XCpa3VeJKzi/oLm6xWrbB4DTAvIyTSIuvo
3L7zHSE4nNA0SkPRd5D0f89Yu5xHEE1cpUSre3WWje/8kTueGRMj5qAvOfo7PfNX2TP+qslkgRVr
W7MytDF4UlB46SInGGWuAfdv0BadOhZEnebRjC7UlIZUEvZRTBKKDOqlHwKkV9YCrEaBNx3Lt3Fz
YrFax+G3/QAOpdp5fkIcyhMufJU4NOq91nMt+UfX73KPmzH1oimFIoe3z+JHsjZoa3dHxAZqX/yX
yt2PvFoVvmLUYqe7RVDUOLjCnnl9mbterU9ObtRRDeAPDvD8KvfthYKffqJtCLhK57Bi/wO6dGdo
ZE+YYrnkOrk53dJJJZpXRuoX4O+OwU5HoIVS1YmFb5b8GA+Dcf5iFl2RY2HFmi/qE9fZ3Do+K1SB
KeWfXFlPGTtZ6gjRld/ltyjHQ/TeojW6utacZDf8PGF5NuSFrSHzQEEO7NMfVeKrbJoOBN8+1eiV
ine8GgZNzfZbj1gZbjvNfUaGF9rE0zgZd7hMpQ0XnS1Kc74G6jQPHQLU/AKMRCmNlOD0pcc/iMxE
KscL26Eo/pVcYJFGjnq3ZaOg05z0Z+w0LX0bDUzVKIptJB86T/fky+vCthESrfG4cmN0DhwoWt34
zrSFhuf1uIPIelvDIZSqkC+x7nJWDMZu3fNTNgCGBqBvhBNUks3c6SU+GltgN3FmRJGLfizEdWtH
RhWJ6gj1S1jVHnKr6rSFr3PIqhgkb5qWewNT3U6Fe31I5jJBAjyZKeZMuFhQB8fYgN8lq6n1UgYb
JceHzjpmc1ddmvBSUOkHFeb0RDcZT+YNlwSGR0R1g76gMGbK8fg5r3/nFOJlaCqYiQ1izwCCNoWX
OprHdcu8PjHJ52XKVcxqbYFKrK4aBvArVFwma1KVyKEv47GpeTcsim/tXRpv44Vpcuz+ZSP0zByU
4feI6th8RCuiaolsULfHSVoE129ysfNN+qyW+syVXxEcLWQkk6JSbacidggbzpz3Matcw3O593LA
5vMd+VxKV7c24N8LI/mpYSXFFsjvJE7QFv0zTdnRhbpfMmsITywY7ezAVpev2X+GFchd34FnCSic
0GGI0nnD9w027smAW41Xd8ZsB3BJ1KdBLoF3CSvyuQk7HF/qLfMtEpVtTMqwBSOJ0B+qJ+HeJvLd
3POwmXLtUy7GT6Vfxse7KxAqso53tHOenIgkYVvUXg3+2NwuLsbmQx332A+Xf0Jfe10050myYEO6
C3WKTdVhybGMywcwhBy51f8vwVXbQjUBSY0HvT2jhvVL9LUad6lXlw+P4AomkjEMxWidCsslIBtb
KLAYYt+faWVs1NtgTlWHHdlktDkZxFAp7Sw9hRVPa6eVSkqftH8dT6xq3pPuOSSXb7lNukBokuFV
cS4/86BW6K6obHo2u2v0exTXnXC5E4aWANxC3ACuRvAtsm+PJ/vfFe4FHNhpZBbEt4/Ny+9MGmDd
/snWii7q+ImAhYkAPKp/sNXNkGLfuzdnr/aKsUc5MEP5EHtXTSn5dZ582oET0D7CUMABwaNReaEj
C93U6ntRUJxK0+pkr2Fw6QYZ6KEtDAamkMYC9x+gcdfTQmdaZtaMTrpjOKJjPzNUU469Is7iJiYf
ICrrl5sQLNoX6fgZouYRDqkLD3oQpTJ/nkofiUta1c/4z6FJkrN8mk/SKn3DUAB7Fhco9L44ZExI
7b2kUM74u/qtcqcZPAOe6C1lyFoDL2u26V/wm4ngc3w2yNPphcfrnQ4No7b8WE/5v8+W14KChA3N
FRQGcDoo/er2DQMiS5iE4ud85wexVcMV4lOqmg8NaeXiznyKze3FIHDBT2PtzSVpPfj0EYVNEkM2
FlJ+ocqCNx2z+i39TvF3aGNgFcF8k6DKozDZY68bGbqNQcyvwrC3eYF0C74iSe5OYF4pwa5u1LWl
3ZdsqIy0cfrTUkRM8416JszdosZ58+C5ZVobzQZ5zE4JukYAZwNt552DrSQtLzuGFKe6m5IKV51h
ASDQdC/1jrgdslU9+092IP9o8UwX4c4cl6vV0w6X7lLpQOTcFvxfV6azB8YqGZt7HI2cH8MxUq41
VWd44+RIhwseHbaZQ5Kd7rdgDpAHxp1Ark1KNEHLNt8XpXZwKtuRLakJVxGqlL26pxgvAjn1De2T
hJWZkipap0D7RRzgmm5ei9nNvW17BcG75infKcB7jLX4RDOfLJKc/6mc1UufBpzn22vVni7Z3odg
I7MLe/88Y7NhovKZg6zhRJDBBcN5om6IpqMr4rZAaRWaLqFRFC7UPR8+8ylFN5urPdtW2V9gfEDT
J0zYz3461hdPUGauaNJ5nhs22xdP9+dyzeuuaNKp9Z9R7yLsvisbt+q4P3GuiQXXL1Bwy8jAmyHs
HHutRc1LK+WruC+E0Z6lCqFfHgrw5/XQE2xGL71m3UUaZBDl3mUCe9p+93vxUi5B4+asBakVWqnf
c2or3Ypq5ucv0SApd/ZBdv71ohiYhwUhod+XkksiEsjO66MLNqBgrvxDaXhRzJv3T8TQ6Ujr2LPF
yUBBxnJGr71EMr21oJ38BFpLcJGjsvbJ3rtwW9zwurl+6baf+DX5Nt8wSjk9VoKKtlsSYipaxFE6
j0NFQlb/As5zg0RmbUrcmrwe00lLPPKLBKd7bOU88eVP36loObNzGo/rmtDbuzNU9nhakpALRklj
9erD7wIMqLCLAxr1qAB8oMf841xj0+TQqTQ1Fl1X1kyeHxjL8d2neBD0S3/OIKz1CVYz7qxwC7W8
uwwCrDS732jUeIAt/4+7Vg/DD6hlHBDojBbsfXzQCLQU+uXjF/24ZxGHKRFAG/VtkTVQX43od59I
T9TGttnVTClOFeJDP1lDMeeBbvsX/Ki8RFQjRZ1BNopVH/ifTp2oetTJBZcvm8ZimkkDEvo+UqZe
GibfOHXws1OQ6Cam7uBqIkfggvgFfOrip9rlRgfC3CMUGw55ijj/0O0uJ3hXj/7hyj3fYmoVCXjw
R8vOMOFInX1QxCwxDj/ql8L6FzapL0iIN6ul6NXCZ16r7R894zrUhQmZvXWZYuDOHbjLheOwNiXm
uJSCbOqgEb7VYJ1XXxNPj9mru7PW7YtZgQWXAzbBOIgOML77b+5lVsFK7O0w37x4G74RvmQXzxAh
IQp0CbdubbJfG7F/cp2ObcJi3pS7iBV95ihTAxUVvcTD4wnxxQXwgL9oYifWEXQF8LGUJ6Q173ES
UTMpZczcOgTxgfneSQ/4gWYwPrRNeumVhIeZWQ3OrOIdPG8r+wWIGfjE8940cSgrwgyCtCDoqWku
w4eOhFb2UIGcRecvRptT9mIvJhboV9wD0hPKWo2BiSUzat2fc7yz3NCKVsMHPUdjsH7db9mC3Byv
edkvW5WVWBiAf51CajbQbXrJJZBPjTtx9y8kxZL/pPSeaQDWY8nlWWXsPDUL30izZBvSBuQ4DAqu
Qw92ZKwuglJKCKD8aW6w51tBzC4tQFQYNYtOwa/GfFkQ5DV7vRkmvjD3Fs2/bUAZwLwPreEUcH6S
VWQpmmhMUwS5X6oOVsTipiJ5WTPOywJQOz/gCzF0W8NfXxnEsgpqKqWTw5hvQDEbnmN3563VbwOJ
8c9s67mYBTw3SNndGnQHNvg98rR439ScAsOlh/10SJidoBAD4Bf7Om79CnFUOZs17r7s8a+0QA6d
52iKIBBgvY/Wm8HnxavGa2ttvaIlUe0Ly95R34iTicGrK9+A7oCq4LCcOXAmn2DMLwA1OmbYgX9G
XqzAuiQ8VhKMo/oJW71Axnypdpccas4+h4YU4jcX+d46c+834Gvs/1EtJok6W6PiHHqNgPmjucFI
0Ort9pX+QlmMegcbXCco26lUeBUx1P97To36HAR3AsH1GlCkrkno2wrYZ/VlpZXt4l/91ozpBu5O
koofIHnzTYkf7uxd0YpG81uU/qGUluTLYAhEPSQYJhc32MozkK8GF4Xb4mzP+PkrrOJTRmJtSdhY
Wyq33GO2FiWJr4P0UTSKB57DCypfT/PHUUABGHIdWARtRZUI9bZD8AjwiLr6QEd2aHQS0tWX89qz
h248VKO+irMFmaskNuulYpQgAO48qh+XWVDu2ZL0peL3M18SIXWuRIfcgQ0DHRdSzKIVbmzuIICl
nPZiyU+2Cq0FETk4aFnJcZh2l7YOET8hKHk7l9xLSISARm77NTqgUcSFghASjAR8PPuLWVnRg8ZC
yop1rz4tkhTMFrIWpbhvOnOkeWWD+/w9yDoI7kj3yR1gQKmV5CCNTZMbsihlny+BAEr0PGDdvGYk
joICbqzo+DKF6JVXfwf+PvoVL/RVxYH0pgs+/ihx01/auxIXKOpjwrKcayYMARTWfsMzKb4Fc8i5
84YZLDdUhl5J+myHfOepabggjSNNzmgW8n5sQMQHJj5q+hvagyonpiXjxK9glsueSROHTaFS25ZB
Lm1QB8lvBYEKw2/rw6ZRQtku5dx5ubLdibGQP9IB3ymufeuJhfT4JuCVVnGvzB5YwUiULmvnhVMc
kSt7iOdR+2qqeIfe2aQobGQ3DmyyjoI+UtvBe7N1rWY59Kdg5ks1CRa04ZQMmSF8EDZ316CBxIbs
5Yq0bxt7Ww3LgYH4iMwYjreM/QGJYoJ5KW9+LHR6MPNPoPqX4cXz5h22sgsBeBlKFln21kg+ShuF
hQokK+3kt10UdkaJNccOn+cPN9QjhoUKYNPdUsBykTfOBZ27nF/stVuoy7Spq398FE4me1Jz00+i
dU52xOPyDH9nZ9ZDjRB+mBl2lvUifKHjiYBdD22aJD9ulhTK2Qa+pnJ5uQEFh71bjdvMQ4sAy8or
ZyefndE8YSxeCE67Oiof1yKN7UHzpuko6DVNqc4RXrdbB/O6x8TuJQfwWgvfb3E2/NaWMFbhgFX4
ouysn9EG306Xd7ABhCzJJqqT29f/0uL0fxwn0ZqPSY/mAs/1t8aqwnXHU2cGK5nm6L+kQcbN+YRY
6N6xIMHJ8raNypwYUOtJ6wW6ra2MJUqP5/5M7QGZJseGF7RTTHYqrSdJfuQJL3uQ4SkOHxu0W9jQ
e7yQQKS0zN526GPKYyQdsll1LJy5Z4fLJpo9j/O2t+ubcWIZ+U4Be3j5gLXKSWtCS0WsAHlp8lw0
+FAjlHOTWxIoAU4fYXWC3HbSk9kfIS0A03tNTHkXLQ1v+G7iHNm1V6ijFr462Jp6W+A8LctfPErI
jm1JOOZ3XP7lSRbM53kD9H7gph0m19lW8MvJMNtVEsHkTu17V+ocKwcmiQRQQjQJhF2K0+z9frIJ
IV9ddHLNoyxVEjCvp7m4O99n9X6MunaADCgx2HIilo3pGUIaZMkOr46b6QCQAeuQyMNSi4uyIh5h
sWmtbZSj8hw0N69d03g8XkdLbd0p/6i2HQi2lpGE+eKCuKsi6dQnzFvcq1EzkrG3ZjBFM4pRtmVZ
0SYi4RGuGrK00uGPoT6Ky0XeaC7WbVK3pp32PkfKqKSJ9iVlPCHxM35peoH6Ld1sjfP3WT7DkvoY
0X+8lkRrlFsu66sAJYiYXw+TF1+4TITvXktL8bsoXe/Wnmo4ls2tikkZF+vW110pKPWDvr59gy48
6shwCxj6hYqcggjYqx/X/7p0zQea8fHGh8TWvLCahv2COVypL/lHIiWnuQZU35DFKfZPYeCIc+qz
PAz5iW1ncExpgzCuDKNT+xJKHnb3YaDmuCqY0zMU2eRWGQDR1stXYJEhk37FypQzs952UUMQIbtc
GNdELxOdKZ5aXXrdvX6+o73k4E70Ljq9+4Fn/5Ipar1lgwiUFjMpn59wLJjk5D6mAcM16YqJ+PM6
XR+3WYJygnxKWv8e6Dd4xw6XoXoSy4ncX1mJvGzIVF4hb/G8RyYwaRCVF4uauDe4aUzTm0fHPHsQ
EmbO2woPSLI2Y0hy7j1LaRuxQNyyH/BTVo4FVTQTSYegtTonOh9WI6qUfff+o4cSpStp+scaKEkv
eETmlrVJqiXNwFVdcTLqwybEEO1kxMY/EWhyp9r5+W0vVIhRLTgZI4PtorNnFC5Dk7D1pLnFySS3
L65xwN+3PwaaXovBWRayCOYhz7ImaM3v+tgjCOvpaI05KCwxuyLPmDFvbwHRsqCad3rYgd/RDTdw
KUzgrHjeH7aJBeh2kupLIQ0rqLAapHZkfiv3V9HsJT8droyU2o4cdkrz8Lfms8zhq4fFC+k0tzQG
1DKZRfjtZ97atE07SwWm11h9iU72AWjgsvR23DtfUpaeNd93N/J6JqR52WYr51HVWlPXHl+USjHl
0FhnvchqXpnfX+L0D4rgxdo58msvjjWBCiW8vS/T41EUpkPjgyxOoGe/A2Bo4cX9j44F144ZQpRo
X1a4KPwoyFgGdq9VDV8jFXc3PRqOSK8hBpwPCvngrh4seJp40lRoaktGrNp70HHW6RKOpTg8ekMo
xsaBA+DCLk981UpclG9Zlcs4F2Kij+lwlJXBD+ii5mRPX0NvXQ/EAB4f0AUx+EW1Y+y3QUgcvTTy
GcdBaHDsQP/gkk19/LYh9GPfFbaA+j94ZCQS8okng/EdLn9E5h6eYWGMlQXAjIuqpeY1GA1pkcx7
CiZPrdVCDnF8aIs9Ohs5Wdtu6eiZXaE0haNo12rSJmn5R3TxvGsKTcT/kL07dgCKYBV2FNGR3Ds2
VFRSzXl1EOz84wa+hAC23b3XXjZByc1dZbgV8TAuhqI0XF3YnKxSekxHmqsF2cUgseumD77ADMeP
kocOTZykoaI6v9wtx1PWtX7AdbL2GOpbqQlhrgB+om2uZtPwrd5x/IEYenz5n/ScyJRXYzCEgIs/
5YvyBUg+PkCVscEQpi1dKqM6QI+TNz6KlVQvz6nm+1iBUbJ7Eg5rkmC1RNJugftiVd1QHrUd0Jxk
gHd7nvaAmgOAnPtuTLhFlBEjOAvPdTBxNXHqU+27K6lx23/zvhGCbOidDdZikABwAs2GBq7vyyLz
oy4XSjCAhYit5Ngtun75lAft8dL2+tOJ4sN2Z1IVHxeYpFjHmMXYQSAqd+v9hVRgmXCiywKzdRNz
3uAAwE1UlCXFfvzx0EPJ/VsWcBuIEuSeipdgKfb6L5iGOkudavl4xYXQ4YUrM8AIzysvRfMTg6+m
RBoeN9K2BVZgmxhndjfaF7revK25eIyR/nGqfcrdHsylotLvTuCT5yayY5G3IrXzOW9Zn3DyEzZx
vNqrLQ1CM0UAbbr1s4quX1BXB26huBRPMJ58pRacYn4THAOn2Ntl4ejvcF9NLDUQtfiaItvWJF2G
k8NKJ75CJ1vtw4oq1JWUv9PfatG/z/dL9rcjjF9U52zrC75uObvJFlK8ue/XuszV5VVmJnISAD25
tcxh+po1ZqYdE3vf0QaPuuPmMLkIIHQHfEV+FaC6fAPvx/YUhZgjN+ATXgoYJO4fpdXEe1ZgVVAo
KERxcd46HEki+5Itpa8k5p5X0PPH3C05G1XBERSCAaFN9gZvwIGR7PxM8n6C6KLAVYeiLb7zoweV
Fbp17sBnP9zwQBeVxyvLrZ2Txg0zLHUMnKDRyj/WPhjW8y0cJ1A7UC1xAadxSxhdCstvtx8XOxMa
aCBc8mQtjMLQxmTyzf+Jy1J8Y/AeC1NBX4/rRq6xrhPkY7iHt7lzx22OfTBQsnALiVxcD1CFyJKR
/imNcaf0KuHjgPih57vMA3hu2nod8fjna/HuiWcj0XMIEVYFrKOnIGlfCth9YRVwQysrduyF2JsH
YaKEEeWMjcmhNC4hy2c9/41K+W/JovjCK2TwPqIV8ZQmY88v9ymahDWQT6pFOQHuWvPdEHl6/u7q
e+YMHbIHhWVdhpEAAFM468dCW36aw7k5TBd9S6B4Kzj2FUxnYKN+wUO4ZFN31RQ0Y118s+Zfuus+
clhf1EIWMvP3Xduc9Uodhz3YEQI5phpp76Hc5LKrxTOOueGR7WR/da69z5rQ0alCx5kgJkZoHqOM
DwxCv+I0NkNsTE7tHOZUNAlwqZmg6k3oxUuf5OWmHxfX4hAWtVTnh+lDo5qv7/bt0L1+ptzXvb+1
Tp1oBVw2BaSUddx9tKGmIEWspz5ar/R25nMkumUgvTcUGJrNG3mNWLW6Yvk+K7Tkwn7hmyKgJViS
XzRSJHlE3wj+qIyj4DXmgS40iRH8K+v2qyBIt0ep799bBUYEdF+zk+YxSJRaqFaJ19w/uXyGA/Z9
bf02FZoISLkiAxQkMj3Om2lryznCnj1gKm6cz9Al8J4wG+7xnRe8t7cdFdqfg9fWOFUpJO4sUr55
DBHKjTZa4s4cUBKDlW8RPOABzCwwmaLXKoPYeJf5gsY3qaOq+YvReDPZuEghQ+NxD7dOyTkPMOlY
vZ1CxjEmDh6vpeco+7yDF0hrz3G2YblnLY3tz3N2UW5J9nwS0wfz8c8dQ5Pqln/jMe9GjAjPwDNQ
woid/3vTMMN+PB1t9+fuqDZ6QjPa7s+9o9RGWcSVD026PquHIZxt2r2TEiEcH6SRuOhBpRLcaczd
GvrPnlV/Fe9nbrnoCBit3GNCbNMzNh1crkOTipo/2yOrAD2L3O10ybeFCLKHAx+Wi4BulArYZCiJ
ELFOOGs8Xx+6aqQHeKTqAVuZy44LGel8V0sgExPxeNJV26o0rCzKVlDy82cuyViwk0pPnMhOm/vp
KlzVkcmSlCCUtPfNP8dE67Qlumljo3UObaHdCMTw32j4hEMLqAb0e3cCAchgrpS83DneDQIzL2gY
NCsoJZeR+pm/xi8XPtt1PjPb3ieTT0f9bNzPi5Ns2cdwwm5gVjP6nfcaQZN4Lqz986687ZSdqOOB
LJf2u7535g3OLoWHoRnTmwT5lvz1EUYuXxzzCeyplAVNoBWsPbNAeNmsjR86zK9aU4dkCoP5s8Wk
VbPrSI9P8eEnlHXgi6UtZVDJ5///VEcYtELHgSdkGb5WyJMaXbVRmrhB665exdU1kCOleprcnLxU
HX4Jc91UFfbm1q3RA8WCkg9rEr4G+8pC1JHRSDJZXje8HL92cs4bjeG1OhQmlkEsphrzrK44fdcw
9kMCD5K48in/JSWlayIHw+T0nWfvWKqzHWJ167aSn0vHvlcz3gu4hrZ2hjbDtMl5JWJjGxMDw0c9
pRw48tblfpwbSl5jDH/2btrSzUEUhDkFfkuoIj4UdBXUfz8OchN+I1EQPsg7YKiWBZu03PSDOmEc
cCAAvp+mRBUbrZ1rfzbfVXBRg/lIvNKYsNNlSbucQO8JlQdLNyy2Nw8yhdb3Yg+2PZ+0aaTRUfAa
tWMU7/1MK0UZ/hC937zTtTnF7b8MR8E51//DgV9jR9FoBuTOXbdsQjRitMbm0t+4b6qPYRVvKazv
GKd+KkM4EwWMRXQM8xcifk8F0xlYe0TGoyTQRpPKH1DhZhlAYPHDS+hB0UiipSA7Ha2mwj5JORG2
NVy8To7wSQftHBdH9ZEvqVFdzI21nFEQHWpmvMmOiRvG8NjvkAOOYACwCGkzF0qrivPk3glx2INt
TRPqK6pgXHU8mnVSqpAxqtE8Wb0v/F7qtFJ6wX8WZ18YXcRjYZTZyT4eduZj5Kcs/5K0zKnChfIy
E3ANstabq01n6e8e/2lUM24eaN3G4bvsiLDHOYEbzHhMUgsVmGOunxRUO1Ix4QUUXGXmz7/5vVNS
I2g2rEoELMyCa4fiYFgGlnV6/4BUjGMQLjgWCELloVCqSn/1tnE1u5NMyqcHBlbvDwyTDHuVc69R
vevk2WXhLjiRXlHzDrMgFk4dnv6DHQsvAbW+swunQxsaZ3vpp47Kd1QTRcnvPXFF657KsoQXEouB
a0mtX+dd1M1BG7quRllthsEEYp4+xRthUgsXnvk4IKyeHz7d+h+NGbcHXhlOVBs8V24XSy/9Lnqo
EuLZcyWEXMmGG/RASfct3k5ghD42wMcOn/lNk2wlHHx7LHK0SkawxF25E5tSkso934Z3dzwz7K6S
1yBqyLsQIdVY/K5c2XNbTyxfWk3IPMuY0B+jGQ74x55cEtgFHzR6LWRHIS0B+uStL9Ca5WqH2HVL
oWELnhrgX9U2X2bVAcHmEPFPZo/c4P98mKILkkOleB15RwIwaqYiQew1UN85QnerpaI5maGqX7Tz
o7DTViXWlA1psVorScgXZi0YXsakjgJXpthLt45YrBjDbFVaXCJ00SxPJt6KZFXJAzVMZCe4NxtQ
F+/a+CglnBDAzTK5f0mt4tnitcpnIY69ofljmgvYVQ5jRusKTUOuoxNVYYaW+zlURZV7hklJ1gr9
ykpBU+4STubeDGFX5eaPHXRpLT5pJa9fhW5tM7za/3cHKQ5IcA7qStyEjvuzeO3RtPF+R0uxubzA
dxhOcoq1HQC3/w1FOv/g9G+xbs8DH7uzmlGNWGqRxafJ9sP1j6DALo7o/ecW774clOMdUA9f3yYB
lb1v+LuECBLVLbn31hlVKk0ItG+ibh0G7k5MIZa/LEbfl+tVy6whKh21LYk22SVW0Xq9ABIsiUnd
0u6jKqaLSQNUmXgjtnTMXJZ/P/kaOWLfcQDRXtF0Rqum2h+TUP7lwtcWb63JUoAGokZAlXZeVr98
3sIvMcUiWVLKmM2EdF0yj6u0zZzg1Ksg4iSDTyastXx2OBBHdU6nP+MYI7By/kfaopcmFv5iv768
yrj1X3ucJX9iEDSuyswg9/y+RFjjLbCpXv/1G62bQUQ0M7BQaWYNBgaJu0nf3b/wQAiak9k8QAdJ
YE9kiGqCTsWRIdd5kkSgrTLy/gT/hNMQ16nnQ/HmP+FcnptSGIYZqHikk+6mboG7ZFXfI4uG9Zo9
4keXYhfP5DYBnlKqCcl3s8L4MbPHAceDekSn7jraEUVUknjpy6i8wQfLBKkqyYkV1oKvlYoDBfTS
goOkhUo8V9QicZH21pRJ7j0J0iNVU5knk0X0o48HdT5vHWzTqa015Yr9LzobjJ1TUkWb+63xWaEc
NtKDFNR3ENEO9ztPqhL0H81sx+rGH9a48RBRqQnfovQft+z8HIUScuc69NCw4f31K/Asm61sRUCe
1VxmdhrRpY3M0QN07k7Tq8LK4nnVQN+cGE2CF6Ml5Emchx8eKqpdkzFe5WIxGZaamYkTmIkIMxhD
NNpW1Ry5HNx6BN+uw3ibi25EMjY3ceMHDC6iuTpJ/KlZmenYiIkwtwkRC96D0+iVhYpjZiSMF6tP
ZU4dWuHFJn5ggfOoZ+XRxVzYSM3ZsGreS33UpCFG5sihFB+4LweHQZ1Di6E0d+MFlPdnxQhlDytW
khiweKab4l7BBzrKkc7+ud0Oj7+KGDBL+6XYgwfkgVc/d1dAdSHoVCwJgWeIEpmQxccz7ofqmwVI
bhjs44g1iQzrjXQO3Cx4v8lxxt/ysvu/UnkXMiQhE7q4m6vzLfPtBRNAz62uSTqOJOOy4HNc33aD
pEzrGKVJ6KHEr3e4C2hU2HYwxv6yE2ShikznWgxVGWCZrXxk88SaTsGvDjOw0Q2jxIusWx+3XZIl
/Af3HyR4mleNWHrcA+wf9lK2gFXK/yYcF0ojiZWoh6yIaP2NSJUqqkBdmSJVP4rYrQZ0suqb+ptT
LYxnDXYQDunxRQK6cErfB1NRPJ5DCpaZ48Qohdl6q2gPfnsI2HwMAb1ta9ZSLLjgZOWDxHY/crcL
kyrtKr2Q95Y3HWFE2nn6XWWz+tEdej3E3ubrt0viCQKZyyhblQRHngTtGfH0EmZGypfPyJwPL6Tc
onnuHwBfwa0FHtu06kLukIJ9Mv6ewIzD1iqGx6KeUUDcDjdlNe1pLM8Xd2qf1JCWqSsfPPyV4gaq
OX7x74gX1zPYMe7LN6mnhfoOVL+pWSGO+96AhYcwuE+tWK7mvFwSu0CxmCgh12r8AMLvaIqEgwCK
32zr76+LPAxuyzdL0NN6T/DInJlVlHzEtcb+X1xPPYjBVb2eLOjxS8YBu/YjuYiX8Wgmci2bf9zu
37S0xI1D9/jRYo0mYopjCNJJGFjPJDR0U/TXP0Y7o/Pat4AvaZGnbjGcD15K+duIRc3KLlsABHKz
+YBQEIK7R1hbwKvE5btV+lgH3/rtnihtRMfnlwkK+HwAHJEzfzptBy6OFrfyacDIqJ6H3NAlZzcM
RmALl+642UQvIQ5GFydnhzyC6SmrMfZbBfDeyxyBe3mTTH1kk3EEawwrB/R4WURHhX9sSw10SG7P
HHS9vRc802x7lAsSSGnXVtCAq8uAghNzmGYFq5qQzqR/BKunqSE1sMm+DgcSaVPUQT5HKwPLLpmR
NeeSARWgt7wCMeH6g+FMp/bUPcL56kn4HogjzpPp3QQY0p5/Z+DYj+N1CIxEn0t6xQb3ZIwgf8Tz
QQegZVvcv0rcu3mgd8KsZZ7y+bity1YAZJ4oFiIe89zjGj7Oukc7fMCBZgWWw/MH0rxkjEc0fUVc
QEpAcnD1pxLMOqew+8BbNx53A7Hy/MMmlLunDuDW3cFDrS4qsJqsYaBdPwOLfUUchQdch7GukMqy
fEAo1K9M4rjmqNbc97X1XkxVN4pwf7prrFwrVOod1mSj3C/A50sIuf0zRuUElvwKhHWN94ddwNqx
e/7N04BrwboOuKlFXa4x1GHBa7tBvPRmJcXFpa4XtnL8S2Jtn5jNHkvPshoEtLXdlU4I0ohMnJY5
AKGodZgdiv71wQx75LJZmVmSs8PwxatuFMUHIUOTvyGmYyIv6cquSmlfbZ0YXDH3F4KVspLPIri+
9uasmG1pp+xHKElHWuToGqRD2iuNyeRL2mrsPCnnE60q/VitP+P2FbvV8jXJgghl8hm3eRiv3ecu
gp5EKi2op/MwMTcsVbMvejssdEe+ZrNQK9JDFbxzlNSJYT53Dd3SisFvxGcCMcNzg5bqREiBKmNL
h8LQzG4cUBzXYQvTJoEKjtlbM5/UqbsCobTuKVd96MRw9vd6aQVFqhPUNOpQ+z6j9Y5rdXAYWvu1
3duHjicod4fZArmeRfdG8cV/xgObifUb0NFy8GwWtPLxD0v30AGAShqzc5y7w5KkAB56sU/+ZDk1
onsqfpAb+ijp/5S7EGsoudBjtsRWrbMQA3sTCgE1o4s1v1tvwyV3l/5kac4JbwqjQ/iL320ePWxI
WvN2Gy/PQ1Jt4G8sVbutMU4Hi5gV0fp57cGD7tV+8jsfRC8Y0L/IYRBFMWjlncXZBl9yRG8h62TG
TmaM1dJHReBmRZqq7H+UZ8hm5iPVxC0nnqJoNosydNXzCtmWrjGiZNgRdPTgsR2mf4EJmsIr97Kx
84k1z5I5FO43gEQF2+j6FCgJ+JPAJ8zCF+blzwt4X97k2TMvNkxMBzcnmXYRm8seYY2YYaEewxQg
uvuRD5XjXBM0IimnDWy7p+lg49YQI+4sHjNX5FqFw27wuuXWNtJD8CRUS3VUOnGODcJ5HjWGaCea
a7mvtnPEexGGreO3JGoaseIqqauGeaypbrxIiuURfNHlGMt7I9C+5zTbVqPI7V+la68Z7wZ1jn1p
USXSHBXnapC+xszWrrXGzYy5rX8K5ElKHsyuTmQbMQ9sFszrRUSG/zM5z57QTYGkLW+ncKKraSfq
lqlLcuO15mVcLTc+CckgE3ZtYmR1VqllEB3ZHXdpBaNROmbYotcuZTraBCH8ZtF0D5xdmzy+55Pi
mjyo787fH6aSVZvlCWxr5bAK2BapXVaPdalCp5Vk91CGaK0nDvBSk83eLe45tS+UVKxTop22svDY
MqX1tcFSoP05bjYrBqqnXmDyjeJgQHv0OmN1Gzt33EFEOUM40YdO4+jbaHMBVCfUayn/5i2dAX9F
4HziSFEMlVzveBhsLzePJFmq7e6ir2m+AoEwuSwpfbQrqjATKgHyOGGTK9/kY6KhJ2VXdz58cj4u
Cf7MKan9WoAJNEAj9cPPmjJYR/C7uCwBa/K0o+12JLoIaWLEJa3DMC76ZKmVHgvP7F+VysxHtHa0
NoCgnnrG/eHlPMgJgAHly2K7YXhhlGFGuIDDs2FopUAJ+b9oRD7TbMTXZfS0wBnBHi/b6ZPL5sYk
dYsajgIuRf4F1S/QMD5RYRyhpgi2urnBTz1BosuqFR3WiXnT99TBZNd9z+JAOMqQyXzkvOUF0D3R
561mHLhmNAKJdzjMkpVJXts6u2AVGEeWFAqFAik2pUhxCRuqa+gPA+z2fx/+fkFuydC64hLf215I
E0BqzDKdF6guCUh8R086feqn16yhYK/CV7R04CJ0Qt/ipFHYNgYZ3VU56fCcBt+Ud0Xj11FaVVHS
J+oz+RaUSynM70Yb5mB+nfzp8+ebh86b60vsszpxgriqs54RekGyQUyxxWLHZ4u84S7bWOejXCEg
f+8hB83LKw5ZnkUDCH7OIT8VTdadSrPFauCtofM+iw0+m5RbA/y8F0ctKZqpoGj7QxeDgTG2+qCk
utaiyD82QrqzAQxxJezNY5hoZ3V5xV6FRv6R9Rn8VxM5k0QqcRZaq/2bp26L4HFKR67nrcg3YYFz
krhlycSL1Vn78Sxpg03gAYznDiNBuwYB68U/GF4jXIepE/ekHd40cEqWQA7Awvkt51oj2DRquH+k
dXVHRjidn8RL8erpksng8JvAIriomkCAg+FggJZSGQTrzXv3xy4lWT4E4PLnErBiZ8pO4imvnKen
E/rga8S13zNRf+jxO/5CZLO7cHFDb1xXXWsEdgOUbhrQPMKfx0kCfxCVVdZdBTInGCV7Lgsh9Mcn
nvJYtXeE8LEiAqgMVPkPeOn05qpoBzo0UICuBFNBHLklICDNQo78rD9YN+1K7fdf0VVaytxnustY
4+BUrUgsEfj8F0BLBEP3CBl97VSeHbSSWCUqvfmeRrXgOLDrvmhvWNb/SxQOiTVNo1xfhHdSlH9C
YWxmurIeo7fC3KbS3EzmR0eq24AUqNYJEyDnOhg0ektYmqeAmm4KVxL7T8nC9Adx6OQjlhtoUE2O
Z8yHmLQDx1VEi6tmH4dppm3Vn36hKh46RVoiBGMf3pAoideV8h3A+JGtOf6AzZVP8dDfW4878/Zg
dZTd+YybAMfVTZiR7dhqTN12kj71FVqy0z462HMUobwB1FCjqyxpDbsFzScN9QuipZIcCgNgC9TS
oskRb7d3GaELv30ntnc5lQHY53biTlV6haILYwJuwlXmo/+/QEsA47TXQI0JW8LOP4TO8Kz80n9/
f1kmV4MzX+vO6rgghECuAZxzZ9sSJ4VzoeJUfLTv0DY82kNrGSFEuGTSIiucRG9ONaHw30+ft6Xe
/CTuW8Lh0JinR4n/qc+UQNtvjncVv33Ww125p3mIZ0/m3VKcSn8SVF9D9Uplja0agtpJDRLi151L
xP3RXOfjn02U/xdxd39ZkAQmvrCVTv+xDJkWktx8GZ0whHAsxyhzloxlZrG6ZTXPor20L978+Z5Y
lmvm1jwoe+TFTbGWDFp1LxLDH78hFM7VzaVVUFbQ4DlnIEj73moWAZnGiEnNWcdwvAKgIw7X2L6K
DIQLZSMQWLuwjb6XLK02fX8qo4KncJboWMM4wg1JpMKc0htkZwuoh+FdZwVEULg2DN0ZrZLH8RRE
eHKuaNjNInQL5kBcoWztyDBLMXmbQVPzhD+eJhqWboHWO4XUjunZECI/eMl2Q3IY+IaFtFJsjNLk
JFmCut79p4etG0PUF+iTioMlApJOfXG7xc7pFKS+JXjdAA4WIUNr8pGB//+ir36hT9hRqPerOTuW
BidKNmzLuexZq3wpyNrpnyD13t5myj+fE8nLDOmmQLOs3qHuTOLlkz8UHTb0wzrx+3vZS+Vzq9xf
NvVoExrP9Py6qvA0g2jVSv0N094vyJ07KQfuJzoANLgeur9nRnAZTx5ZLO8XWTEQfqPLmWSpX30l
z6Le+Ubt3eZFy3MdB0GSsrsI8v/4T4C6c92R0febDYylvilcLJdFBvWyKpORqd0V5viGzbvE6JfS
DJMTnNN65fGkntO4/wl1MLLLoU45UwpQF1w7rtfWEZuYd/6JY5XaJBng4HwKTN4v2sJgJ5+UgG1r
eAUAdtMJey39458oTEj02Z4fYBf1a0ZhMptDuuPFR9uQcvOSMu0H9NfN6D/f7ieNCUp8IjCaCOAt
8OMQXXXTIAdRZ9C+oSSV9yoxnJtzM011G520ZeVa6p7I7EUhNZzOZsLi6WZxcg3GoUqdSBPewzc0
0ONldjIBA1X7Y1IzACBUdjY1GW4ofLVjq/m+wXlnvzgN+X91R2agz1akjeGx6BnUuXpksG+RizJc
V5c+1ScTjqex+yOtWOFGPW+rdqmmhwHgUP1AB+JPfg+bacd5EBFaIJLjZv5I1iwDM4HDsEXbU3/X
HhCGdBPKa6uAWNXbImOiTqnJYvGlWfsPbybFB6aBXFHs3qpIr1tEfhFkLcMABkyyQ98Xp8Y+5gFj
fZNTZqsWp/X/odOiAyhD197mUzfkiDbhOAWAl0L7JyN7uFCCEF+X+no94XeRD72FNQGRbSEegO4V
sMiCLRGDLgGIZzgIwsaC6RvBhKqIfrrC6LQbesd3yoZh2KvLQ4Xr5pGG/75YtPAKJ1ptxJy6WorX
YqgzX1iJJSRWQ/uTPrU9X/uuPehLl3p8dZ2hiu4ph2K6veTgFSwOM7k18ZNQDzm9bT6zKTH37ksm
tKpGJvUfwgEBhLLI2Aj7BIqYRhq20Yv6WSNBGRpuxCafzY+Dgq4I9hxkDdGdi/Z7Ie2QKmh7uxwM
ICxbxgoaODg6GbRiCSqhoDxJesfk4SUsX7BRjRXfJpO9cJ7ZzE41V3CIKTsT7lDRL7lA5dEKSj0e
3FZz+shj8Odfd7KnUOK90CodbDKAJuaj+ln1DGQakD/uD2Er3/Buy0aSemVN79aGexiXPNHDqyWI
Axmd67Nxte+Y4XkduYtlF1m2x+qwDJIjCeOs4faBr37EvYsxmyL/pxIfaNRe5fKGimLKQmC5I/Z8
D1xbEbLZdJTEXUIPjlELESwglB73Paa6PKBPgLg3MAk/H4iIreMY9yNCOGbTuHlm5libR/hJ+865
j8gKFcO5rgWdBZq+q6W25bje4oQ/xbSl8h+9vgkDv9LSVdKoyfhE4a7xUKe2xx/OCSM3cpPiXRWd
VsurlbYVVclHYY1TlKTGN870TUYfb7VYoZwgGLZdhklEUu9MDW3kHRTSxdW4fOnzrKk5PzlpZYzc
dKLMBJUMqCcOHrhPll6EhgIGGS71wkUReC/iijRzhP1MsDy47/BUwcBbvOBurppHMscv/Me00fnI
GstILMuiMC06fY5GWCHtnFH8Z1yTtmxo8GxHWoL0emE4ExXj7lrNZ0LBIop4E6nmH7OCevrGJsr4
GoCf9tEoHyXMiYSxxaOcUq7OMdvuEp/vA18b+Td5CjzWL55L3FfQ7G0H9uwSUsyIaIe7woymHzjl
t1fPe2oeYUUtREF9DadY8yU+q4/JmSSCeecL3cJa5y3Y3O+nrUTp1JFhTfa4rvZHHshyHVSVGvU2
tgn4pYadSXvMr/XNP6QAIxE9zCekra7TMY+O3qV/s9cz8uBCRoGKjCAi6sgXOkLJUrFyCFScP7S9
RXkNB2zhg2dkznCrdGpTYVtyFYw+XlbaX1R0c9GNKudAgRqqt5otCYBhcMxFPLRZq7LbHtl1JvT2
SvMv5QJIBefKG+OzTJ0A5G0SfzhXEbh0+To79AFTenU+TimWSVb66lGBmXvV3Aimmsaj0yQ6YBX9
D++yIuHbiZwX3kKm5lZVFXEb50AF0nFEkEa1jiVornKCcVWdLoHVRT6b5sIfCHzIOdSEehm5SD2L
cxpDnV7zb5PzgdRpDgU4LAj5zAsa7ZCP6QuOTJfd2bvdkfkxE5Hf5dFq18lJkRjsGWj9fZqLJmSJ
7J37w7ahvZBWNfXT93HVKylLCzgGiLlVVry9OdZJcsa6PrVCgS8WjB6a0HqBj5pNnwvEISeXSbhg
19OOM1Qv6p1hm7m7xMi2inxBWpWuj0oo1WwL924LFuZF7Kv3I3X4LPMaFW9j0X0mKaJkQRbekZTc
5IF1s00A+wxZdCBxdV+S61D2hAIuF/ljrZz4eTZuNPuNwoDv4KrkeNyBhbTuNdsLPoyVSlWh5iCa
m5xbFGDlJrRzfXH692hHP/jncICrCV4NbzOQ++FnefRURW9/VtE4TdO5P5Wmazh5aYyBXTZIKsF5
yHwgC8dED6LVe/33kKJOwwoyMmookSqF+cgV5ZA8tJ4UOyS64tSOiHY+1bXv9VLjvIYe7TUQTdM1
Aq/BmNovMpsdJu1YPA+pIVTjMyUVcOv8uOtWKEFoLHCETNfgZnHkUsO+1gu4G9P70uqYwyMDrs3q
BCmpwM/BggrP8IuhtganhlrSYgNYKGJ6dLDX+TFoTv+h8sTFwiN0kEF40KJocNSEJ6aXWv0zkDAZ
02T0VoE/K8+4Xwcxeun3s1DN+KjfD/TjrraJPO0adABH+HmjgECjOUZNmFxqsaRzgtvIKHjeOL7l
TqeCpr7D5jv0xiRyim2cZiyhGU+e62gkzsrU1wWi9FH7YAxvah05H+G/IN5GQS2XrL50+LENpj5t
r6DLpwbR+yIceukvCDiiRcm+beL6Y+ii+7ohc0X4u47zYZ0uftXtEChb0bUDRmO0ET7gaRLhRiPl
eLmj99QwxCO88uhWAsHCRPOmeEz7BGVR4uqP3dv3KaP3XgyrROJ00B+p2hGDM4Qu7Sv7jP+lPwGJ
9ljgVQ63Mxg87CiQF0ljKXhjOH1AgFm9nX0g9k6ZfH2IRlzpSIGI7ZZbiiTAILRisjikN8hyYVij
TSe/7Fz0p5p64y0krDOLwA6GsULkuTJUbhevW3S3LmjDiBWEKlnBxNucCs3THs3d2dz5nvmLyHMK
8UmLGCv3E80rHu72Rh14udU1jkRM3X1RbFXKy58kTgVKxhU2ypZ1mej16pJKpP7KtNVZ9roZr6HG
CmfQzlqZNJ38RP9o9v9cllZgl9ZqxzVBCqUNl1irsnvORddf0QR9YdcMC5yDIMC1d+88glnIaHgk
SiUmGo5+g99BNanO/B2ZjntXDPguZ4XMrAXq5REGz+Fy3pza3aZgWAiCbEQpSmn69hSkwmzU8xmp
a7Q5QorlZXy+OM1JqndwTCkBM5avTK9YlvwiELpjw1R/Qb3fdlan2sBYDxz8AT14pFLqyX5RQuDl
pOfPfR3aknzxUAcdZf/rxSjLVXcOV1fhTco8RFa/Q/CQHRyta+6sNFISJERbA7hK6t+pIhBQ8JSR
LvsRU5DhsIYvfunOCIUlNGckCJAZX4RBk7NW7A7mo/b/46OQDp/jghUAuj//sbzBs1NH97lSe1hv
fH/HXUl5z+RRDIGPd0V0PWbkgNq18vS0f5wpJM1rrtmdeQnTZI6h35XYcyKKew9vOlhEBPbAGZiQ
PLXnh1CYcSA8F0zhWSDPcXl4tX2V9qFFgwJfaJM+rfqNl5IhLDuJAUVYD29uxTMFFZRmzvvaBA/C
E4uX4vIqk4MS0mZBBj+I/Iwq+CdggNbOSzByE2IM8RSJAP/Ov3kDzzFnUh5RargguX4OAr+yYnjJ
ZLsroITYDcmeZ1FwPGNfZBi514ACVoGtZrvgWbFrUpXxZ4ywJrZIQDkQ47YAmBgJ9AwN/dIcRRd9
CnC4lSJeTzRKR4PQlcOwRsnbv5E+YXkPB97yIwA26gyMGJUdoycE9/MY+Vuvlns6Q+1yt1kFKgqC
ds5GIS5HMWfWjq/V6athaeuwlSs7ovmkdTX3B/YioliRrjNbbT9CKVsXwBnHw1WR228Xs//L1Vzd
o2sNhpFGX/b3aTJ+GpyvbGZ+x8IYFZHF1DpfaFGI7St79Z80KfLDkPj5x29QWpmulXxQKq7fJZSR
T9OMqHjSiXruEKzNFreyMhDH85XfPpHKhRziCgtDXA9xslBZM5Iz4qDcgiz3/PE1gCs0lA4UW4Nm
Mysg8eosVUGbtHRRJ5YOYMDFEJtiDQs2QS2chLI8J+PemWe7RK4+xhNpyJYHAhEEs4vgXWYD5pNK
CWxBtNVLdJXvJj3ja/ur+BPj/nJw/08cMa+qIpN4kggOExSf4FWtn4UfDdnt/56aRE7A+gWP599p
bIANTjtVieVh7nfF+V/F5r6Tice2NdpvKwVG09kIxejZNe5/j30zmlX4AAlKeO68Vdbke2lEcZ+F
B9kJQMCLGNrZcGExOyBC6KwnmgmWKH9f/OgPnJgGOqY93mdVGNTRtmFChMl9dbPYw1zouPqp1Hp0
eOJh287eB4e/A6ZAsVgPEK0tVpS2WOuftv0AXketN7xiP9JwtLh5j6PF6Y9/5xGuBqMT3t6VlsHJ
d6buEwkI2gYp7oqH52YYPwJd1yHILpsr82ZWnFqXHZCMgNVMJdOkUojWjlxSusPxhumeFnouXCK1
0uL5NcU+/309nGHSZsadGubtgeSciZH/SFLboqsAR251bwsbXqmA5Of61Go9pV0piCqEHi8i34hk
RhWd1MursIOECPk1H1xGOtGpZVmRB1FfvPj1h/dh2rBHhhg23doG27FcLkBJomnrxcD3aKfFBvDI
N3uKvMbxyDkerIjVvX3C8VTAafo6j1hAn35U4dqxkY5oCSp83q+OkT7Qn9WVpw4gurORK7jr1Ya9
Pg/xJYdZRCaxJuLS+Tnk6mzXGmkkMqGbGPjA38sGXmhn64so9bh56obSGhOVGW6zcsItf3VZprWF
rr42ONi6d33sqcrdQ4Yz3myBn/SqyhYDrETa7heD3cMrIdcBFyaPVcBpRR+q16Rwy1FF0HKpRL74
wxR9GoaluLrv6nqdkGoT5BgGXEpwAaWOzpjcOlAhCVU6t/3Z4taV4qJ0BBzLI0ymwklde32LCF0N
8117P5MVLcBdvgfJCfahxSBYdy8UXRZ0LCpZBsUsr3LNrpBn0Ivr/6wUYmuuor4bRXzjs1thvfBk
RshDxb9yefi3OIPweLaoRLJSRk+0aV0Jj1ONj4Dj7T0chOxmFOOtw77mPJhxCWVfspmiBbkeW5yf
zSRwuqsrc4wOS8wG4yQ56d0djrN/OapV7fj3em72RBCIKU97uee8Sz6z+xcnw+NdUpQHf2BaMHwS
OYN/5pQcu+WisEU7C8VtkgDxDgJ6XJSHUMUOEC/chrfHe8nWO/4k9RnofjD4dAO9o/F/ii1erW63
vnjfgoRI7WuqRcvng1yzKghSuj22EJSnKpvuJfcL6GS8BIOU5Ni7veLfjKga1yZyYB6mhn+4HaZu
aAbSziqHxySUPDJUfRpJk7BC766jF6uogGlM1qXGTcfsT+gFhapdqvbZFlJAgRQNevabIVMb62i2
z9VSowwrEkCeQi+eWV4x3jyxqtJ3Jc9td+cvSpbzk9IKHLqVtLefmu1YzATP7fZSP9ijKeHNcGsp
wgSyvUqziR3pJIuLK2KHJYIaCEw7bvWCoYDIVXIe9FytksHs61HgOe2sy+UYgnj2y/D0OiExXUDu
Bb9WjBpXb5wPNMVh0jMHUfH3jKUsmLAfQKCGbDE6PI7LeI/bjgV8lcmzNv5uSnw8iwS8rg/ntudN
w5fotx0R+fr1XStPahLZzxZAFwA6rAbfrqpt8QGduY3h12QDiYTr1kIRVg/xc/NuIFN02Kdk/L7P
B5XMQFPJ/KuK53T5neRKF1mD6JyEELziVzv/YMxlQ2ulkH3X7IhfMJdSaNtnOTZNho1Uy+Xi/1Fx
Rznnr27HY7D0sTi4BwSSB/7e1gXS+ry/kbKCuR8XKzGbrAO0WnxVx8sBQg3KfvsohgN0QZ3fXYzu
vz24A7QcjEGXukbnRBA1xaqe4ZSGm4e3DSd8z9uCVZEuFI04tTvm3rkgvQnLjShyEdy2XZQz2DPW
zUKJmPHGN46L2452pM71KoX7oTurQ6BOk4IKqy3RG37ZE8p7qStUGZRxBiDKpibYkAC2T1Afq4xo
uUnWU0wyrIGvdUBs6ciHqQt4EybDtQ9cMAfq+5qsqsc1tTBh1nFAZtzbkIJEPFX0+ZOBnACI5AQf
atL2cBHlVO+SoRy99R4yLL43BR0Blg+xqwdQMikq6xLslcFTQriowzRiCV5jH6MuA4D3fgHiLVhL
7zVjHj0lcYgbEn7eLQE9xx8Wps8rpjEesJVBOqODSsLMB9rUB3iO3C42hpEOO/LkDVdcumpY/Q/v
fQOfpMGf1PkQd0q0CrEIl5ANu+HCEPdHk2hLs1qZsyiPZJ5mo2sevVB5U0rxdKkon+b3s5Jqmm47
7oQBUQyv5rd0IcDHEj+YmCN+hlEf+xNawT4XQn4xT37otfcL15AY/1w1sWbYWJEfE/IHHml0i/LL
LwrJ9JwKqkJ2XeZmD4Hg1TN1V9w98mdoghV1JhVv3WOZrhJR32Gmr7OorXGIGURTQQqXslh9UXP9
mAUA6PpgYI4vMV4XEUB34CTyGZXAvHbuAKcX19VK7s8LwBqGfzeH8/UPAtFx6T/xvOjBfIa9/zNX
T4raprC0uP2MVQWEAFPUlcGy3gF6nyMV7r75yb5t939ZnR9moT5XhxKv+lEsPY4MOVU1HQHh4Deg
zeGZ/sBk/CwATwb4X1HxIg09v9IDNL5JvzATY7mjSbTzEBvSYFaKZ/cMBozsxldWFH6y/7uqsKbz
ODcTrFUvuYewq8b+OmdnlGDLyCodS2tAS4Wg1nF8hP7YeUb+ubmSmPZeztuZldTenNtYJlOYBzhj
pAbqdLnyKuQQgPLv/7Kyxg0U1sWs6kvm9NF64TTEGWSW7nFfZcy6A8b8dAwnFrAsKT5fVRLX4sL5
fB73w5SmRKK0wxjzsv7x7gItXHq6QO8YzGHgNxS0iyjpFpogwOkYyBVvE7H1Uv84rtqRw2/78RRW
BhlmoKc6ARkut/OGzALOXrg+KGXE7aXyiA/5YxM40+PFEDx4ujyQwXELfXm/8df8IxzacB7b+ULC
qmuba78C6te5JbXGrXK2Mzmtze9cKZbzHte48jCW86BejGQ594429OGJOBjQoW/X4qxdAiEctosv
Aj1mJwTj4LGmsm5WzKuuPrbORkgPDYH8yumNgeYad3dsu8iQpx0r0pE1VA/FDTd0I0MCnoUeeA6h
epKcpM91o3vDoSS00NjemrhlqJNAk0QdJqmytdOMgp8ooRdDjMkvO+ZhCeFHS0Z9/ZFQ1Z2ZCWto
HHhz+NkWMiuuG8hTtWqpcvdSCQ9aLnjcevGdRzsoAydqzKAjcqliVsXQ1PmXdzkASst1760e1Dv5
smOzu7BtQDoRhcFozcfMMXbxPH5+gKIdqCw/qE1AiOcYxDC/0Hr7R2TJkL51CzRQF6ghryKW7r2L
ZkcPVup0KoFTvwQHv7tKUMZduluWqFkqvMJSy/X3JAww7YuQDcEm0pGnljvix3xpiaVxp9zmGiG/
+f6AJPsawX31/bFXJJjBTZKfbDzPWMDGMRpBV9DBahj4GHi8XNE2AueAjkSVYNnuKVsBsqPa8p2U
1TCBWRzynfIZhkx/gUq30vMGoQMBmO4Bsno90vEvBRbz/Ng4waRzp0rht7I9OLCaE+wFlYqwswZI
zylrjLNGxPkwY8yrStYkAV08tadxAAZttsXcuMilfX8wipfTuMPfYoi6Vwcmnx+61Q66QwWmiB2j
cnYPBlOwpySRidxrbhwV7URYn/e/D2hWs33uCHZW+98W/Bp9n3d/zerJ0Knk/7H5hYD72OAeSbb2
MMk1W3NJwn2zixxREBj1MtKKiyTfmruebiQoGDh4TN2ftQnhZyyodaEo46zuJ05YeWDpLtl0PjMm
T0Diexo28QnqKlZ4AnH3yrIIFbJAASRc0waUA9ojHjHc0YKVxr5wUVo45J/6DDyEvSlIAZ2HtIjy
xtwrwNZQIMICV7aHmVUKACesxYNJHlOJ/2D+glkLp1CMcipY3R2LRTKOKpirpAzHt5hQc2Y5Ztl9
FSu1JvbyoUqrcDOUYih0NucFJMhT3Wmz4UI2s7fhSvR32RZBZTY6ZCPjgl+wAZF1E1Mbvf1djOwU
6jVu/glfnRL5i/nMgJzxvr6RCPCJWQVR0rYs/5h6IqRbrViZJBhTZaQQVUSKRgbugjaqHNxShqpU
nDc9aGdTPs8g8Z/L0WFoHLtJiVKn45fxIFtYbT9Tp0abILCyzbwXR1HWkxNPk6sMVGRxdOFH556i
tjgyO+ijN5/EnNxHKazwqMWY5HQjxbR8RooQhA1QGhr3ziT1lae4fx9nU9J6ZMquahMq2tCYgsI9
FnqoHoadVgxIS17Yy9/F0s/rVyls/k3LPJ2Ieq0b8RTnPWZEOUSDiigoNIOFI/DOI0jpC0FwhA12
LtuR9GHBqJO4LYPktrCNLIXEM1z7pi8xsOlrdZfLVhppxS6RG/6Sf4FiIhZ28/0Zh9Swk1SP9kMw
N+UEsZ1YB+vq8SwwuwRDROtNgiCFH+7Apb+Ft9Qv5tHZAVvyzP4eU1F+XdL78KUM2hpOUvSVSdn+
pxhNS813C8GgCSzHb1eEJYmVOAI5QLxfS/oMUOpKTAPQzkJLqS+dyrMixWkBbe1xL3dToWEd8hIL
54sQMBvczO1tzFgOUlQ96XTcDGnGoN2jjeT+zuMm7k+S4hEkAmGYt8aW0JUSBMYWdX+NCUZqCf0T
jOj8qCFjFciFsMTc1PXWJOqEHbcloLTczTcANWeDv/Gtu0To6V+vxNsQEFuCCgxwfeLIEYuDseaK
iibAhTN7oDqYQFyqX0DWRsLN2xF42FqVbbolvJs8RU319yyduLwTZbpVuuivV79J36XicGAkmIEu
3wNu3XClCPl8fFCmToP3TvrhBXeiY8O8GLwvhWY9Df0y5YOJDMZ50/AMozMSiKuOlIl+v1Zxo+Ng
RN9ETGIfJpncWe2AeN8dCIs0Wlj1IQqwKAqD1GClYhNKimR8+Ngj9Eu/zNYfTUSL4eAtaTfO8Eos
tPwIfezocdMil3wbQucnIxhDATYfylHD7+IB2W7AR8yLVE28upTNWdSOjH1WzdQkKM34b5iQujr8
cDi658WAC037ZldC+RPwAI4/fyjJg793osajx9YNG7SQgz/ZdvGfGjvxomqx0Qptdn4GnW+LBdGN
RYpqPiD07AROa+tdxIkPd/sZX0kVPzhZTaXe2crUVBa+r6ObdyxMwAyQil/7vbcJBp6zefY8fvqX
zsoRVaUtWIIcKYRsPkLHHlcqz7yZn7E7aD63UxevYOqjDQzNLp6iW7tWOAk6QmwiDS77Vxr0kHFm
IwqvIbLfRcvjXjNIQirKTJ3r7Q8f0cy7TArgRMMy4cifNLbKqf3AZZn0CQ3hoTpn2rCsM+u9UWYX
3cjae8TNd44F+lzhMS1ZtOwZrm+AVAyemvMdMAtwFSN5+wumiHyRg7qIebfWBUNSD7BBtSti+1VM
MCGzAPXhTByQxy4W1Fp5qcW777sftnWbUu6YIUY7NqMiNMJsSCmH/UZPC454xC0KvmAvtA4Qmcxm
6AnyxlQQouF5HANdzNHL8kfL2S/xCKF6VK69sUu50T2QdXPA9cur6krUTD+uQq1tKGCucKRla3tp
htApcVnY53HQs4LxlXZG19/6C9BCyKplNce90AMXeV0uPxKUUNoUSudDG21sIUanKywrLd7lzdMn
PpZ7hL6Qi/HgvnfSYx0RxWU6UVwyyHSYBIMd8O0XDF6EXR4EXmjkrplS+sp3aAyEqYeDV8qVco5w
kL01EJb2TXStCNY694l6WZJZdW4AzQ5ljYq9yVxsvlWDy/4GQhdKl+57GPtEKDEJOOK8gm1TEBV1
8sYopAVPe9/IyMQCHfWE3egdQA4FLrz8VQwYxYhe/b3IbhnIpuOsvJ10Twxkz0fnzrYGplJmRAvi
u18AJfYhDW6P5ABOcJaOVg19dUgBiR3nKP1OzFT1T3Az4MK8wEsJrFTBpEFLGstgYxRdr6ClO9Ej
Co6/6fY8Vn3iysJSmfEsU61DenK0CegTjmv5hLbQARe/5S/389B7qdaBAzROGNzudGEiVHf7ej2x
cAvLJ4L+nwtb0Yu6j6Ile4a7ZDuqiLTanYtaLnBvHdgMyh1BVQMUG+0qyU/4QI1w5BinpY7hmo9h
wL988MFyPPgqrbyDGBq+srG5k4S/PHUd4tT7Ss5AyBPTMdAF9iW8/6bKASoBoPn4XXvVUcr9JPMD
mV4E0BjRQIUdaGeiozKe9CpGe2e7ZJirc49hPD0rGuCBp7Gv465pDgnSBx+fzeevKDtR7bY2XyBZ
WpZhygdbR4oPUdj3mRHEvNYy6XNoCMl/e18an6Y4+/eYYM17zZtVl5TcNbWRRFKtV+uraR4y005r
DTTSDDNaVL2RwrlKLgKYeCsicnDeqa7ZlfoK8xDKicGgEN2NGe3AXXgEUPhUvYHBHmW6rKMBq7Yl
M/RYFUjIYtdplEt2qLjwy2w9m1PPSnKXmEyh7BrZLYkF3fzqvx3Zi6TrJXDbkZa5i+t1YiRo1YXg
+OZBNeBkZ8TKEbnVUaI5XXpwGnvSehkOmksh78MsLvq3X7qXoUNkhJcMbf+3LW+YCzEogoS+mw89
F7ip+IDnmFE0Vo/MzJKWLszYceM9HeLefWgSnXHpaGJnuP//Ett7YGI30YGm5QunDwMdJsT5Cu6y
VL3BrFrNb9KQT2XxRf1jhoI6hPCBBTZT8lCJg8dj7tgl5K5jUEIncnG2aYm0SnEe/oXJZmVIl2ki
UYhurnv+jO0wlSuQD3NIqy+KKJ/TjZxrA0vMRgxZm1GFMJMBu+RNeGKu5WXlqZs8c4GY943knGte
qu4Cjfd6ik8U4PIFCU5zvrj9h6IpAwzna+nnrl94AFmBOzt9mpfofkvHMUFLUXAvUu9ZDsH59XQl
o7m4mmg2BkZbHgwUT1wrnCtzy/qtyy43QaeEXo37hOPLrqkHxtsplZrFJJYT0EcOUKgnfaweiyzW
RU3+ZV8ypPQCOfF5wycu/XDz5WaW6VXSBrAPrc2Y2tx8Y1YQAQ97caRFFpIewgn8z2G6VR8GMm21
cVknZzwm5MCqbAPEkdXU4WGVxEATROiY4xtmlih1WaH11psU/TjXslAN2NVOnPHv/D+8SBjGNWYq
k3krdg7Fgin9TOpk3BWTkNsycDr/sYbN9JexzRqS6OWrhrNsFegN+WmcuXnaLPUwUwkrjUpPzCv6
wsDWS7akFEW5GKibopw+e4C7NALY+VQNpwQ1BKUueEtjPVO1+SUWNcg0Hn0JqaMVbisECQHSGBcF
IytBH4O7JBZxwe9kPwbRh3venoyL7IWjsSNEH64XeKJqetoMtaAxLXBisljNO83LXnFTvKHqZwFo
1kntURWSLmNk5teWWCu/u/8JP21yWbzwhjH+noR2h7AQ0SN2ToU4pixqhJFLYNdb64Gjm8vGTcTq
CIt6OK5T5Pep5Q3RSmhTK+tQcy1pQGFPPIyIodUrQ9+yc9ypelwkhn84QxfoEx+ZqjmllRVYjIB5
Pd8x9PvEGQqmqXieuGW1wMx74AGwHruphKgnsX60qFrzU6q8oI+NaLEYiCB5WcemcM/yG5h52hU6
Qf5jKz43opj7/FbEX95DmJeN1mcZ7s4Z7I1siwI1c5BgFaeWcOXopDXhmKKTIDvWs4JrnIUCN3kf
De4ZFKLEp+BAtoYWW2Mg80Zi4tMK4DP50QD2OFj/kBagp1J5GvbDh7pep1kfJeA2Tk7t2yu6lNuV
4U++0zIdQ6pVc9P9S8v2evdzujxIZzwNgJ+gqb631D7GHoVW/YeGBbc1pYLuWbGKN0b3gFH3vJgT
8Ou1r/pHtzzzmVI3ey/rcxBS8EwyPzxKjRtfj0uwJYxhsth/l5uHT4+QMTq3kqMQ9ywZ2xS3B9nF
sj5TPpCWQ7QcSlu2VoJ2cXTWwkzPw7yh2aEmDO10H2mx4Zaeq6/yWje5no63jLP71Am0AO6ybK5T
N/Q8P/O/jcf2XdczCUZEFsMukthFFAXAuSHEc5xyYnKkb3ApphlWAJK82dS5M7Ucq+2+LwITAd3C
zMSKMLlwFxkdrxxrDQyJU1IK7q9hqkuveTE8DS3sWvx4ZMJ8FQ1CTbLTB05OZCfxRDA3VSHPfgaS
16ENVzXLlb6PndQEKq6b15rmtUDdyDS3+f0t5bZa79Mglk1Us620BarlSBKKV5ZIkS3uhaE4Ql6t
tqYc9Kq34pSBUXjnhvLZrfcdeDyzY+K5+v22hBoXxLypnnnDtmkQ1mMUOqDzjPTjL3lXW5VUO+x/
XH8T9TfhnNanyoy/fufFXSchZan5a9tDcWaUaCuNI/4iOTfOdYtv7y3uucd6jEFpf8ZGMzfiJsXW
rd4O8E8LU9sYaGNc2W7kZclKXmhlUxfAs0um85M/HP3F+UWhw7SEwxJyHCeghPsnm102zjR82/xu
HKOHZeG8+V/jy2wLtKq21t1djCaDQAg6uoJ6TV+1t/YWJFkWu88xQZwK3oF+grXNt52FbsL4ifTU
JY2vFitf8XcA6jQcXqz17p1+RcSq1FX+0bZ9qX/Ejj+SCSOHBLTU675rBuUkjl6yAAX4SweQ4Kyn
PLfV+jlHqTb+NkyZ+L/CXABMzC9gLE7GHEw+pWF+9g7fK1goF76T+UdpTt1TMzXn3gPRCYaNHyIL
CE7CbACmDyE2Cr2MKEmE1tNu8i0xSOC2KF+6VOeX0tstJdf+TnkFINFZvDah5taihsEq21lYpqVI
VHhDCGAAj/RR1rnTgq33fg/gCCXvWX79xRXJJSgAroTUgnr4APB4MBoHmw0g4kJvD6nrQ18l1Nve
zVuIKa6t3CBoJ4lUdemFsIWaGf6XEiIQeeXY/8UvThpd1M/aJW4K3ay/dcdNOMvVTHFy5NbnRX4d
pL1JZpf8oUw2PeJS8t+igLtJ/wu4SFUdG1xrg6ZTTjyBgf2yYDf0D3HwkoW2vsxT22Kq1/5nrVrA
7vgp9dVhgZ00LDyKaOA4RtkfLjPXuMaP77mBDoMtj/pyBTOSA+zcGoEXEbgtL8uDBBWEde68tdwU
gSUqrI2RqEZJZFEDFyq4V/2Mlmwp9qrSn+3vipogo4qtTWO9/SeH7voZ0fvZuh0k73PuCA/tqcQe
KiUoKqldJbV6RS99tqlI8stp1rq3W2gdBZ8HOC726wo543fzCNvjXquUjlDUORNXtZYvaAIEz9r/
YlKt29l/nZLBjJlsWs2wWcEFTHfgFkH1SBYo98hVCuNHV8PcyKvOCbyyzblqd1qA/5DjCFbKohH0
iWVov25Bel/yMrL8GUSZQErx5Nqck1j2P64OeKZe4727l+4dGbgMYjdnC776yUVoe1FIRCm8FVfe
aj56fYmMp56rJAK+7mYKomHMTgvz7tZ1Jz9vGN5N9PaBErseln4BT7IIKrEzu5DXmxHPG1NOmqjA
4LG+mmK5xSRuIFEJvFgvN5ZPOJSp0TAZ8/GP0GYcaf2fW5L+K9t7zGTQCtp9Mie2f1pb1PdFrJy+
7klsTXj15f/yltC6XxR+18M//UdAux/M1if1aYp0sNzPSs2R9tfWYOm+0+wcsXHsvsB3fgpnwmOp
ipXIRxkE7BiTQ1ci8c0P12RUgb0oQZ73Dc28LGPueXVYoW0CtcVB29LUGG+9/me4Cpd4IGw7udJ2
YxL6j+iHeqmSmNEfz2v8qVCdnyYMEHJ9gk0bnyAK9PpXi8MAPYNj4rFaPTCEkXQtQFpAzFzeG3ky
2vhUKWs0TurZVNAUyXFP80JCLX28+5xBjRAnXqCm7NNPR8+DTjk5ms8oYA367bEJm9d2QBGNeb0p
ubKnrX4kZ8JHCdDRcdxVuMNWovQMhvePObqqi78lvcEFEyQAigipv8xnWRQaH1H3z8OK2wKM3mF0
/o1DanpwPwW5/7uORnOqX+z33xnR5Ub7fAqekulXz2DdfhClbXxqYIAOCa3mE1xNxW0YrkBtfCmn
rdrtLV8EYNC60ReIo4csffThu24DwZQIS4FU1CHkZVobPl43CV4Qjdrfy8eZS/Z93I7gjZGh9Qpq
5lTsNIT5axpqbalaMhc3+j72wIjc1cmWlRZkUcHgORbjP3DlAqUUIDTOonj7WiehdKzXM4Dtit0F
Cnbb0pHYxSwibyd+/6+JDv8LCiSympgT9GGoxJkUQql/ODbLHDFWKSjyxMNFzq0IdZElxJnoDIcJ
SA/1BHF5TYjLf4Eu+LnbB+jovO0ArbpolpilgBUlfttib1OuNEuvojS1dGGJRRwhwTElYxzRvfCh
5c1jedbUTy6o831uT7ENgCuWvwV5VIHsvEBNy7hS52ufLsEObf57ZfyDi8NLCDGgFLAOrxDXJQOc
m1MqGpjCzeNJighomNa5nDIVPhccm0Qk2KcQ2alI8Ptz50bmZVGi4PPgNUP0TWjjPWrikO73gAf2
oituPVyw+036CZiF9s7dGD8JfapWabjxIRfOJMkeXDkzRsgaz06nEbXKmsqvkURohV9RQuQ0//A6
7PXwP/Rp3+zOXt9XbSk3L3Dd7M+UEeZcIf2yNyqKWwODHla/ks3QlZGQT/6VsFHZ1seqFew6X8Qq
f432OS9xZ87fS4DRXB9BkNZDKXXgYJqu/tjMI5R8FyzlaSHGhwek3cn3lb5BYLXgoQWmWBq/4rL5
Ju67ZDfj9zVtu3UDtbKrNoSGG4fe66sGZQaKl2Sm40RjXtDWUdc5IiGDBlQppL/N0C/ys/oonh+s
hd41f3B0WEt9jaaIRJCoiUZBftwafm7abhjUt4+fgBbMN81Vs9CbneygFqLqtpqntmLp5sfa9+D+
vD8zloLDRkiD+m7msq1ooNVScUmFBypdbfZDDJyquShKEJ2dLLXVoq+H/s13BwuVmjh0FtUYSgG6
CQsaPDhO6kFZfXvKeE3IEyA9oZGVWeMvDYnapXaY6xl6iPztmwqhEc/TGgErFUpUyn77tB+cZM7T
oPM1lM8zH2+NMMzTDXvmZ9iNEGdqLk29D6l6XshbxeY7m7dKGzGOTBSWu76U2c2pVyN+gSB7r4VA
kqXP6+TFpRjdPaurCZh8LkDBLPrn+IqmsF8fbljxpTZO2bifYtiLJgi2EXFZl8dBQd7o5VoBUal5
2xaw5pDvvamh57gg62WgxuelgR2WVksZnB9HHPXg4vA9Ek3RTWzCW2clvbHMSi53Qfbos4uWsj3W
KcCNmXb0IJ9hrcF0/BTo4JBJVjOw3UjTU3si8aM8APgQMEUWKRQD92gbcNrW+5zTGsn7IgnmGCP0
t7TXv+QcEi8OseoWjVDzQeOQ0RsuZlJ+yOcOvOg1zuHtgwhurwMsaK4110OyeOgLDUHLo22abIb0
6LY+iyB6uaDjx9R/JErQUHp3XJhOeFBCe7HX5BZ0fxiBqObj2SrhvRwO5tpYAgNIzm4Q0yL33s69
CnpP/bmeCKspmrSrrYaArQWbfil1/c1PlHJVNEqlmppqyuij8TkOUTjQGW5UwLMruJJGQ7wGIkGg
rTYUD4BtnbAtDktF1LaTV+7pbJdDnfswA/Ylqbq3FnnTsd9CICMDQ5ptUAiC5YBPI48TF3LxeFdC
IHiiaXb4/OTS1LQxjzpOgsEZSN5g18VxgmD6evqPOfdAHvpLyRxCIRIDR2g0gOEAwfMzycCIR3b0
BnH8AJ7Qzzi5BaCtSlrN5BG3rk9ZEd47CmDneKuGJFpS2hiSMIICTXggVedm/APk09t+Cj365Yql
f4b1OXPyYrDgaoWP1skOqtI24qRWZ+mgBSdPMaUIcMo044224AJCYKKQpk46/aDyu8knopEULvZk
jzXUh9H5ks7nIf/7CnFP7iQt+CYioT4+dTegMdyP/9T2rqnDL8yUaT6L8cq9YzPkpS/P8om2HSoG
NSnlz3hlBuIE5S18tlSM8JNRRoBpdNVoSb6oHORPwjZlfqCjohWCxQ3iasIprrmZNGAa8ZkvWTcR
b9cP+jLnzuXkRyENJ5zH9Dfcy2mI1IVu1oxELrBRg+FvaUBKEvtlvPb4bAHPjctiG8oz6t1H6vMg
DllItyrPyiRPNjJPJCbbT7THOamZce5xIYp8gb6lJgzwjRk09IlsfuAlrOegmPf1P4CgkzLYKhKt
y8CezrnrkJhhN1dqoFnpwd6ngnqJLA2uyuwutXCv0Zgq6FGOzCfjDRiuLBdm7YtfCB9NBObTFanw
YhrVkRka5MdJQLmpb4IyoOsgbSy/HcOYPBaTmFk64YT4WG7FTG2Kbx6HsZV32/oMpe7CQLBKcgkS
D4XOAHp0aMO/jc3/cbdMAjyxNfR/MSD06a2wpIDofRcYyW+jmVKNsWJDsQkInYTr7aMx+FhDiU6s
tFFSxiHslWbZBpq3QXZDC483dypeCgsS/o8CBN9iNV+o4ZWo7to6UIssxOdiARqC/kiwhG9cBEPo
MoCcC1oX0BICuWOaBiS5VDZa5/RXjqcqGaOJ2eDD+fbG/z28CqB1F+xc2vNtJ4HztzhOJZw1EjtM
H8PpWAp9/tSDkr+byjm41liIJxiQJ5aCZKXZoDRaK0/Oq+WYLJ1jquBAZEEemUplIeZaTQlpD1fa
XFnRzMjXo325RyuR9iP9ldbaD9xOyNm35AFiuByGhN7Z/LMjk+kZlxT4yWyxk2wdDwWFCi1Xkgu+
0FBJYz98iSc6aYChZDGN/vl60J3dLocKbVI+fR7WUg4N14IbQH96yx/qi/Ufw64cFJhCTE6s0xgx
ybFHY6Jq3yhlXDGBeoUyTj1Z8q9snrc7giDhijQhBQpNN9riNrbmGwCQLLXeDc3dG0wjL60drRvR
c3jVkssPkt+kiCeGMGU4//beZmKv6LvttkdPtcJ5UNO9GfA2PkgQIhdeNN4xgnnpcZrG97+9OqZO
WVMNLHEAZ33s3Q0iMi9PedKUPAqcr6laLmoL5iwp1nRa9xqI59vQVZk35sy+P7LRxfEQ6QU6obC3
cID7ELs+jalYeBw5iUqPi8ED80dg30JD6+ibov45bwnkXfEAz6aOVUDUscqYTGNnmByCyEZF+QPx
zE8ieZDYKwPC2H36bizUZhtwjkBEj170bPUQ3qXGlHcNZq4zYT0igB+xmpIAIUGfS8csCD7oXQMo
YHt67aYCd2fqUyKUlyxcUnFbje60zagWMU3ecx39YjaPRNB4bFBcbrWp/PZNAMjgjYvy6boYxm9f
Eobcrxe8xF6tB8XGalJmmn2yJGTUQUFhnM8p4pTbOOyttsvSE2r32ILCbTW0DAVkU7/bcXTYCCS2
BeJewum+jvq13ia54fHS8s9GgWZjTxcO2Nuz3n/HFnmOKRmUAw0UOg10EFFCj4j+FtB9gjEjy/J5
GeuQDzv6jhQCGl+sK9QUXfNrpu6ors0nKnWZv1qViFyrY9GIZIMiMKy4s3xP2guQhciEJFKR6D1Y
CH9w2XXzWNqZApxM0s0RH7OaJ9h9u97NzZCK/yWFxQF+dT1anLygFthb6eiSSe7J5gYmFDZs45ge
fzZD+WVKtQFK8URLVvBydXWv47ZBuc+XYstzf2fVIWHLaCaoxCq3WTMj90lSPOafL2IOh43xQKMO
InA+qCPQmON4A9xpjNsKNTqUYLa4svQWJb3oAo2tpZy0a1GyrRPuYd4wWKYtWvWCpRZV1hWd7wdm
f/5O33Twt/ODjTq1EZeQvvToqTaAJO3StTVLpetg+6/t8vJ8RQs8rq/iMU9fFM46BkQ0DWrmrhZs
vBfwoip/dzFkycBYSLI7/rciN7qmr/zTo28A+Agvgy6POq4aZexW3jDKg4bFlYWWnuiRY6AneJJH
oVZIna5Y2OTpDlSZPusxar+9wilgUXcUTq1HFbKd0VdpNLphLlDSNWhAttFm6aNTsfEiXYb0BTKK
t8ZVbQeIHsnd8AFq8jUPwrc3CghwKu6tR0uYfBTVDYtmAL3/NGMgNj0odXLPqDuGXhOVm2fVRFbl
pL82DLPEAqBo+9EhaiI4BoFD+2kEki8m+44D2OF/zNoG3P4sPXwF46RFREvud68T0ZJSevIxcHHD
7ny7Re/Ncvq4dMBxiq1FQpfa7vUtZk05dEA1yeX6LxxnBZfi52aXhE0fy9B/ciKcbmOnDCfn71bj
ncyNgfAebKFKVV1W8XHB+ud3LYkANUCYhqo0FJGILPMdELo7QO+PS+zHE4JEnSisuyr7frd+5tCx
CmKYwZG1/FpETV/mUpJkO/XO0H7PPHCQNtX6stnpaHjtI2zRZjzebhK6Y1c0rCMp3T/xa29YQmGb
WwdpgNNQYYeZ4o+UknZCM3BFVh3AdFnqAbRoRUQWSpktDBD3Uiq0IWaf8GtKRiR0zclrraFYBG8x
7K+sayZRMTTa1LwW1lTrHZskehRZaQxskdzTVx401NjF/ldeWLoKoJheuKQp3x/9ObRktSweHW7w
P0QLPAQ9ZzbZuyjZ7QjbgzDTydYjce6QjXOMvZg8OabXdCpZxpwIYlubuE6ptOQpWsb4UwbfNW/x
zISHnNp5Sjmk3EBR1wZKxmSeo0mR1x0nEks9DTzanEVlMXP59RxiL+smuo5sjq0zgtwpqabs2/8s
EJm9mIvDmagvdFVyiCkqInOfJJeQDgR/yncGIP2gUzNGFch914donZhCptODIzB++Afj4XWw8oKx
5NJGFQyCLVvzLrQbf8VzZwtwcG3qeON/8klwrPeCNqZTuBg892nGAeCe+ubEbsQpH4U46AesGX55
gwYxLiZ+4lO9DdSdynF/yH5o+lXrQLDgq97K56Kqjw8LK4LfirBGj+og0RndJXfyjK7ut/4l++kr
Q+tmEKjF+TykGoNg5gsklhvVSS/iD4ie+WMZn2vGWnR5KRPO/rRkHHKSUMd5xlW5+cN74EzQ+yOi
gZPDyLQhPq/BfPt8U9HlyoozZh7MWwV9ax66gxUaklkEq599pRrAwFRE2E1mXITqepuNbvui+UOk
ny7W//kiParvoUvE9Ae6gk91PeA/v5RY3UZ1d2AwHetc6aE+X8bNqJc/HkBe5vPpvRU9yNpuGNeY
UrKeaCrbp400Ux1xgxUos1+OUrVqEZqGKTZ9ipa+xK9Py/iPt+aE0oW1eHU2h7tahKa06ZfjVnKR
JDwJbT6PaMH80Wf/jBs4VijETqqRExJut5LvrLK2XA/mSILFyMZmS8nrqGSoBIjK4SeYjwZRxn7u
IW/Wfe4+ZNEcS5M7iqBZCDrUb41sgWYXG9HEiA24z7gR0TQtMal6DSx//S5QF+OsC8osn1uJIu7a
0ukSTTAROLhV2YFJyfTcws04h8JjUWMM+4Eka7IfF3m6OiNM6M4PuOHFmy02m/kfSDUdvRfGkadW
3buBRf9KHyUZojymXsLU0QYI3HBPIyBzjvfbweGhH3IVtRmfJn+DfWENKti24rfmGJIlp1+xCWbj
VPzYqRc45qjf/7ESAnqXjL7FNUAIOg2au2T5hc479Ag/p068GGcVrkp2UghX7Qwc7rO/aVUkBnFX
8O6BN1mpSDWGPnOgCrFkgzQ9/91wsJppNF2XZUleIwUTmHOxufLbTlSH9AhDNBkgMNMUekkNmTru
72ik2jpFFh6dUohCOVz2y2P5OQBURIja/u0LHNEqxMtvYAXSwZGC50ApV/Zujex91NmuYG0mHWF7
VUKLUoskIQ2DVBFX0UTXUHgQPWCnLlZKhgB4yq0ciNqYGMY33xXRYTkZ1Yl9myCYeM3azeJH3Ek4
pypl5q/+AE8A56VEBWt2QbvNKuy0tGxASdwPk+9UitfM9aGii0Ql9CZSghUpApGWeDn3KWKuCAT/
l1YrH1XcqbAy2vT/RzCdg6Xl4pF4LU2UAe6ca1HcD5nY7NYlsn5klUxA1ebD56hLC3dKX0kHOwqO
ykVMX6In9CLzvXmZEtvp1bsooADLk/uSpNoshNh3P+HLVb+30BVOhk9gKSi648FtKx89uTxnaxJo
yo65DPCw8r/zZRKteOdK3VtMYfGDGK1Z7kO/sdM104Tr+Z4sivkSZAncglyw+19nynPOIWkxiecZ
nFefw3of/e2up1tejQzzWP/Nznorl0xDzEjDGmfevYMLYrf/Hwaw9wLUnV70spYZ5h/yOmE+HP7m
RAsAnrLRIiJtSfDAjCPt9j2l6mdZRAy1U5ogf9Mq8W1J7HQzvdf+k0+b6xLmOqHjyOc95DmYCyZg
3wya5peVbNmk8yAxrdsX66ZAr5W6vGf7InmKMJXNVo1PbCMU2fVlnjamooHeufgWxTxl7T8jT69G
NGnJjCqbHXazctzDCRtmpi+hl9rG0VKb5r1BT0K4WM9822pWTaKbKqjPR+PTCm61Ygj33CtUlLQk
d3dWsBM3EWKUsPhhDMuEOHQm8WPgF/lm7SLq3DhXqIYL4cCWed58pcx5oZMkRka8cuYi7GET+9nk
G6YA9Cg9vY38kXPWqqYDJppFLwk3jywILJICvct7qLtrQshY0Jbfo3YzntRNO0yEN0CtdB0db7sY
rvBUclIkLpmNDwQUMBFIre9/ccRG9Gb75WO+N8VyqOGil/6/MpY3UZgLq7+zxrtJ887+pMSEI8Ak
E4vK2uutAwXYqgnCok0hPbSinP08x7hw4laxmKJFFjMoYVpdZBW/hG66RdPJ4Y9MpC4NZF24oQNg
+0QxaCMLsNlKwkaLOeQMt/nLgiVRD7vify7Qoern8QpJmYDyLn/4+VFqtDJVDQLLFU/41Oaayqa+
QVahzQrEG8NdQ4dpdcEdJHrVH62FAgxrwemxkerT59EWk0JC/enGaYPT3t2QEyVTGr+LLJ3cfWtM
7PasMKDyzBq1hfNYanM+xYzwM0aPmT8zOlztDlEKDrIqYIOwt7H+qn6y9LNoURfQhJvq496bca31
5hpfqqzz/SwCkcCEg5fmLZrNN3iW4t9xbf06tNtAspOHLZcgKP4COJkRDbJj271uq7pVcMGX3T4V
8rZP3fqArZ2K2TbmrgaXtdfpEVh7b7zumu5b6liPFm/mVXLhJC5encQvmG6wGw9+JCW0/SW7Kmtj
jGIXawim5cnY72z1spBO3RhQWUcTqAcLTwdv2ZCNkuPU4ImMWbWv1pGMdCNDZtgdTcy+kJEDlkI0
k4NexMAanWKFlwty2g0w1/uee9xB4c1ZBkbYRK6BWLR+d0zfUMwoNjfhEjahapA6I6QdLlVPAPz8
9pttM8upnyNR7pb+bX8gyFkv/jLNMzge66NniNblzMbNPO9UDr5B9uTsDz6ykADu98MSqaEslvS5
eBOOjSIuVZJdR2VOg62k0+ys9t/m3DyrjqfuzY3zyg9QuIL+iqG9K/uHQcLNaBffgBALqoPfRFXv
FoWGCCSt422cW5fAXNTSFKX+ZTpW9GFW9HnsZ/8DyuwH2Pgm2kD5GHRmSTgR4An6yageM4pV2vaB
Ow1xn4o+PZoZji24uP8jFLB8ZHt5w4khr3Gft4exFggUg0yT+dYvL9N93oLL8IBvEGIWfGB7QViN
Gr/bXHQ6NlS+OGELhJGDHP5xlNvnksU2KkesjfL00ECHUCN6u2jKqaMDNeWymQ2JPHDpvNP5lVYA
3cABKdjC1QPGNUuBQKcDwMBm2iGageGi/CfFeNlK8Ie6MnqiqyFDy8YvgVbC0r6AniqcYXKGwtqY
gX9umLIUU9FmEbcqSxZUW2+QeM42YsNPaPhPlI9bxMzJ2pZ1JIRvbNzAfiBnDhZlpGCV6/oU8Xlv
ACEWbwuRE2JUtQ1RTMWePDIWFEwFWn5ZmOnu6H50P/HL5LGLWPHHSF2xdZZddw+luDyGvCGlYB43
Ny74G1Mq1ch+m+iVihCU8aTj+dY99UfMAIoOLWLVStnxMM1Lhk8bsKj/g5xE1+4ttruYMm5d4DRt
5A5UjZUO9XffeItBmMY3lzCpBNaxECcVLW+A6GrCz+tMkJEBxzGSmut/Q3clgMdcw1h/WVUMim1X
+Y1hmNkW7hUESiYdm0aERR/CsbhyIc3Kks4UOk2S2N1/mE+daCVUd5afe4mpUopij9a5P4xBVXZ+
MyCBQJuIT+DR9Wyx2pI2PjG/mYoGN4N23awRjclWnbesrw2W5LsXGBsM6RQzpFdzElqIVQdV4++8
GEZ3W27A7PQr6MyGsrNDpwGbBYlDibapHv+LWHLExGrqqLUVAPnocQVOkqXGCBsvoqZ2XeHEovRr
xGpJIkf8j0F0Y9TTphLL2Odnpv1ozSgdQLahEwipwgBO4siQsc0R9Ju69k7V6VrN58JRfRfRLxQ7
4W0haNpfBJZyZwzsRC+0cvz0MBQyIaXPrcMDOTsAjVBxseL7H/DXZbNJWUpOClRZoNfcXt2COHWO
kXRVaKkBa21NfOGVnnPynsBK03HpxuRo9zSSQZO6V3co/Q4KvOR8eTCYgtJgB5cFF/g3ZcdTh4DH
jqRu0DQs7YRSAkLUBlxFiWnFzV5tTMVwufsKchYB4n57IHrMLbTQ//dyoYiA961R+aA/ODJuAyaL
NotBd4XxIyJe5x5XXC9xlDNEyyxR2ZMnwzaRGFKoI5Fn8eDOFodJqKXMOHXmHuN2z1lPyk0Y5U4c
Wxi3QDngQe2vwY1rRxFV1X0+2WIinUoBuU3ZltVtDsZRkjFWIInvONLQj+xmP0y+Ie37axKztYKZ
dC6ebtkjxgLL8qsjLcdA05q3CEIYViMGXJVqDSVhtpkAATJNmYl0AyvFvqhg+0bTkSaKSh7m0b1v
72X8FCdlXX+hCSpqHi22L5UZyWpv2pbe+hcr3wweVUbBLih3q73g/OGpgqM7dzD8enxoLPGMOs3n
ykAdpZP+d/x0aqZl9eRbMZdK72sNLItCikqwjeWxgireb8n3GsOesRwQKWMXcqXYXkAlSOy2DTIS
xTvJ3J7wIqt2PhKPJlcDSeTKG+VcauxxwL/eMc4gjpM2fXjYsSaqHueU30qmCOh53ob0+nEt29tG
hrppXy7QyM/ErFACSPHc57Mw0uQhL1fU2HdYr8Ad7d1gdZCUaSJYY3Fi+hcP/7Uey/gyZyxV2uln
wTiRbhgPkpcgvqr9uFghFdResFmPkTzRRdCehgzszzdVRdg6vggP+P4YFJsoC0q9kkdb+tNNyt+U
4ffiMVL+vlLdO7C15WW9fj9w0XRWdsbd8floqj3k6dIeF8w6mukXGlvwe0XJWFMCw1awaalEwmsW
2fT6uy0V2CTMedyidWEvQCayWLcl3EaEJaBLTlvdZFFXHp/jymFVceWyFj4dAhmroZbdWRfo/EiY
3R/N6tjXcbED1iuF25RI5Us2NS1IppaidBGwVocrHEgHwfD9QJbtH4ZHanhSx05+GL+wfqhKfnvl
qwiLgfs7ftemWgYVAG5UuVS3dMq3cQKzwtdGNxsHFy+ckORdnN0VgyqL8U+ztnZfi+wBLFVX4kzi
LKiU057NTVp3SXVrzP/wdcYI57kc/ZJ0Ht/siQQsTNj5zSpunIPCU6qqXIwnt8sxDcD1jOoucUhs
MA8hrCx35xjRVlDMr3nRj/wdAQtPJpDQaXkB1X8zf6XA2iA+EcuOEjXxNOTqLFn16RB9KCWekQI8
FGDKOkNADtwP8Hw3mcw5MU1RQvLJM22DuI7Bp279GCik0BG1nBZ9hP9PbIF82HFcg4hTcxhSdr0U
gXFuic/atLFZ6siTxJJbRzrNUNIUSNMBgR9oViqjLHJeACuhBWNek8sthtq5CoHgyv5PSfsAKYrc
yy5D/PGjxWl13WdhfOf/3Sovrovuqrlxu3taL4SRodC5ScLURPwt9pTTe0ZIF+uVqjfzyy7PpS2X
gcekMM60iPjih0pKIL/RRTAWuRQ4Pbgjiolh4G3I+K3TmU4amKhNFQ9u/e3laoIyUhosNz9Wm13M
u6N/rcbSZMlO2AznWPQJpi19WoEmdwfZYLmYRdU2QC5qLEDwLhkKfvnlU0LoqSPdwO2a+Yd59vSH
Ve9m8Meh/YJDwV9BSS6niaJeqOhr6dJkELePWyxocQC2QksT7L629r9lfENh0tMoqrhT29I6P9D7
+vQM6bRWJeUcNA9mTnAYh16NEZ2lwveJrtPwjzDV8QbfPujRIJQ7XI7ZFAgAlZlexKRLfJVkqiU0
oeUX+uhmDrlMW4Dl8ld9CwUZbY1IDVuCn8SBdOm0otC5G3KVANoaN/yzi2VF84/AovdR+IfwAwpe
vHu4b3R2Dw1j6ieS3A8fVZU9SubaiL+1C7tclgdl/69B0qL8xijzT3PCcwRePAEecUoWSgJR38Tn
FuQj8P7w1+xHARyqCKD1mcNMZ5rr3wbs+T19SNMhvjHmdJSZk+BMiajklImzQGPrzAy/RagPOm8a
vKF7x7HXLdqTV3fcgju9kGL0KUmZOkH6h4ofHlpdMKAABnN6U8xzoQceCZ7ZWn+uOcJdi0tlNJOp
BHG/D3wpY4B2wgvft6wZDv84xrPYoHkaKlnJE3zn/w04PRsJFcXJ588SFW1LqDCtHNVs2sbwm4+H
m/wQDCTHdg35nK9vWWVeRg/ySDtaDVieaDe1eAG4LsbD/geqeTALqXXPZAF4Q8Ti/uFu/C5Mntgn
ELyUsNeYlVxGproXN+N8mHlqoFXpttj9MphIn73RitZNV8HEkAU4ucYmh0iqs3tyvG5+mZ26pnTg
FlovOKakjmumBDVI1ezGSvvRmt9wws8OG0/UCfUrCcDKQF5febvA32rsGuH1kELUs0npUcQgmRYu
eWcKfrewxs6kKPayFINooKVa04Plc6mVrOVNTwNXgD82N9n6zHZce0yvUqk5Yha7296ezyKWqmKb
y+E+OSKgWeOK2f1v+MEkemiEdt2qkEeZFTAYydz9AvZ6NddcC50I81jC8NIzGPUwOfVTZHqPxn/+
xzfm2gxgirVK0j912XyJYvxU+plVIIloNybazEPkG52iMzP70suv7illeK10m/zugC7V2peuuMAL
YitGyLgJ7ALZeGsH+ptE3isjlRnggbQL04HHU2M3kJ0YMsy376kIOkw/vsn19Bu68gEib4/MWmNj
MglFzT7WB7tHkck9KWV/EQjM0D3di9ffaeHITPv5+rabRaMcRndIk0L/BAHajDVppCSAUleB9yuA
LWhL64MD0GJaBTXlEg4SvrI/9KBWVt1DoCSzGxRQHxGShgsJ0AXjGkYlD92cmJfAY6Mxk8oHD49F
Y/1hJ3Hu6evPsyG40bRMVVj/Q+tRLDdWwNKZBMWmban22Kfr8BgetsW8QUOtquwnU1accQFdx+kQ
6YWF+7usWdWIdrEC4bgNxBhgShXKRwO+w//NgSO+B/1aAHJhfNNhV+zqZy6iTxFcDu+fziPV9QLz
iCyi79vZOW65l/qvnkc/JwWMSE0rdZ/Sk47rNradRiWMt4gQoctoaQc+Tn15uTiGt8fxVoTrHedb
qp9eKi+tjJUDveMVYsaJy8H35aFqXgEx4n5U7BBhItkX/v674UxaaQzTZ0vFt+p6IxOMNc47iNeZ
Q7KVwSAxaNIvh5W/A59Ebk7CjC2mYAg9LCsjj4XoTPT0WbFn48FGJ5GKOK01PS7gFoECGH6pDl3r
2wbT9DCfnz0UvLPpDTRHPN2eCnRtmsS0IOv6m/Xttx45UOqAlOBFXToqonoSgkJlKVwBj0yxVH3n
sGYzHND4nW+0NcPiZ+eHHI7IIobLR1k8GdqdENt/gm2M/e1sY7q/oNccGbU/gXCHOIWOdZ7ufEsP
Qc5CbgZHiYpg0lZaVpHCjyoTUPiACaDeiXboq6uMiGDL8W1MRqbg8EN/NesQ0Lr768dB2uKQfSw3
9124OSySfpzeanw6kCqLShMbmCd7HM4/D+zlzLGUkkPsjO0Uuv6mn3PlyHG8M+cDjZJc8+sykAHn
8O23dl85rrenxXtiuTSKo/sm27uh7gMU/vDQeigIjPioVfFWlsusIX3YSavOVQ7Euqvlvcez78bG
jsmUmOvnxDOWagMRWlde5jIvGuMU7ZAmmrEMRU1pedd1038XDxB0XV69pf7eJqNVqfRezJ9nYJOv
h4cxChbxgbMfDNmpfnYvGyX3iep214IKs7gOHHzKubhdVKb/FBDZh/NLeJB4SHbofrKoNwFsgsZc
1hl9FEo6LrOgvMcPlw6IxstFo8xY6wzLRTvsaZmaHX8Wg3eVPTmG/Tnwku7ctEEfHoLr2SlnucQ4
07OJaQ+nMxfRIb2fRk22dxFVAbzODMxQB3GmlEVqry35FpXFs05nwtThsFqayhwAq15LEF1h8qhH
jH3uSOQv4xNIpB4/9qhMrsg2TdHAoKGg0sMrLGVsEK0EYU2iGyAe1t6qAj4C37ofhBezMMKmN4IF
bx1B+VjA1ttzDbZzgSqyiUPmsYDX92fKFxdYHnodl3z9JSOirI5yqJ2/acW2/8irLbr0gMY5D3C0
PX/+r0rNGJLBftTp4pUfuwgz2x9Meo8qLTfhVunUmuzFq7ls10+lrhKkeUPbbwWcCVnTZ6PRw3ue
XUFpX0a4J6aew/8cUBWBOWA7l+EBWi1Z1j/hlDXYEyr5BS/V9t/+1edogkkaOCwu2Nw0pNhQSPyh
LmTm+cvoD+kVbHuQvi1Gp6LbL3xLetv+7IoXY8odaTnoZ+48KOskdiVMtDnaot9t5RgJm2McOmeg
le2OzBEwasfFrewXNsjB+uduZR1e995YZg1ImCTLLofD5/X2DRFXTT2UbfnPkOXeMlLQGYXpqkMm
gThIb8ioAVnu22GlMEV2D59vnYT659Ph+3Fi69mLg71pMMsN71cncuWimu/K293oMszheUPb+Q3f
VB+4VztFe7kYVoSoKndML/8RXD4eRbt0CHagL0hLDX3HpHK+lH5kcSLEzaknduRA4ZSwqwKsusVa
+Mg1s/YIr72SNcONfZHR+sGFLGNzgt35oMbfL1KgZ5OzJgwoyHAx+7MPhhn4nInfaYSBc7kWxcTy
G11ZwgybZ2+9dxYVsCKoxgKS0NDeW2Ot0tfiTRQEdZcZIChv4s5uPQl5qhUOZFUiCFRTW30VgXc/
YaAnoRhEDJ0oERmd/EOVoYSjnh0y5vOXhHLv+8sgJFMX9iYoYW0fYiscgh8LlFEy2bCx4AnamfjI
sMsC9u63ziMbZl5ZBAuxdyHFlM83jCN6yQY8/UqGNT56zWTjPKZK+0GBW1pWWNb0q3iTWLOQOckJ
/axBPALGb7J0EUBazaOmCSIdMpIBqKtlxVx+p5zy0yKEnhvu0JUmLLX/rhCj5uC+nZOb7iOnqpiy
8owjZslqpyNeqz3qRklGQDzLIJR6H1nmNEBYgGVFiOjF129qwPh1d7ImfOZ/xB4IslQ2kFhkb6Ca
QsF9eFWwU8kClHmInOjVE9W1dVCmo4N4mmNEcrdRGgrBI73dl3ykzeAi25dqhYGy7KPmfx3cxh23
TqEwt4go4lbhEtT4NyKyGb8lbus4F8mMl7PYMmaODWNRc11uQttlqktyi45e1++0TO6+2jT2YA6/
Iqx1pwBrfbefJ+uEtdKcjIPGkVJf+H5vrVzkxzT600MnhAqkzKXB8sELpMCo2GBlo8/YUr7xIWbU
Nk34UIA9KTQa/VYqToXEV+8gbCKisVqawx9LoP+H2c+YXWVSqqfDqQfmSNpuqjseT5jWNuVwyr+F
aax1KRhuyHBLN22BYEUHm3Hb5bzoDalWYntopINH+0nMSqfBPgTovR78DnZZ7VyXLK6PG2tFaWMx
J+SE+VsXmlMyU9Wbu6tIjsVbZRifVYFPk/F8tsCUCVYsQsl3o60Bum3uUQQphEf4LcJf99J+9Yr4
8cE2usZ/TQBd9Y8pvQmXXRpn6g/AQx0bWp7ehuoBEwVH8SItM2cD+gVF5/6ut4JKToIksZg9XbGP
ntSGKBRgrRUQZNd4GekPEJjBMcj1ES1FBTpkA7t4Nn1fbqOa6mUy27RG7mg4N5vT4VJtmwS9EtNi
5Outqh+7BsZaVmZ7lgDjLLwyldppBpw/BNod9Jny8wbKTyXqFYcQUIyw7Pk0013o66gCClXuYGEz
tVDdIqKTwj0jzVoBlwKshByGb7gQUXdrH5GEpWN7UWTKHQgnywucRw28VxY3HWg1XVW1eLMB4vgA
VdSyuDCowve9lvyBhkAfYpM71qbYWFK5aurRQLJ5Yz9NW3YT0k71ae8s45GEMfMMkIdWIHz8Sqnc
WaEqgT9ZGBfFuHqImQDTJvdbsswcf0IU8LkSOdxKshKweLQnox1hhSfr3W+i6VCSAkllMcx754sK
d7cXdLI58yM0oVgY4cdJXF5tJ4KxJ2TeedIEtO4quylj3QQD8RKs6dVDjC1oeZDM+8XZvMPcm4aI
ZGAMocMoPmidJJrrrQVxDPMeyOPNpOBGkXkIfgkJBh6eQdTwj9YQCIPLe6CfpI3b+Z9Stq9Z8x9Z
4ivDVRzAwa4wcvlJSWh6nGhqbZ5q8RrJvz6yBjoyQ1ZvZnBgHXZwz0c/aDJGmsEJRpfYcLbRXfWA
U682MbdJxGBhkVTPNr9+HHSCL+XW3smeTTLiAsiQZAtAIU1/KfFStuyOwYX7G0ZSpqiZ2gTL4JV7
CKxtUP79YKG6WXqIvvhUBVVijDuDDLMaXgKw5ze36585q7aWa7AgkUMumA06+wuXzYSBstvtN0E4
PXeXBCPqak41umzFICato6lkMhRYPEckL+9CK2t7OaBukoBKTRGbr4PkG5b94i3+SB+l18jqkQSr
BGr4EVkHaTmzse+E2I5xmJsPTSiFUbu2ms6wCj2+6ZyBwWShBK5o7AjLrL/2JSNkwxBfXiPZ7Bqm
MgOiDI+p/yIOdHlgjEFYS1sQ1nGc8EkBx2wxu+zm/zkTp+/ivu7JzDa+kah0W2Nh0I9L5zSGjass
I+S1tDNWLaGboV5pv4eCq4AJ1TzIXrakMjPmxAt61WbeHkaqj54ZnZgVa5nvJ5OQ+3sCs3VNJ/Ht
BDTsVExYY8WL8DtrmLd4fl4o2QU/wi6bijuGp0cFPgWQN7Z0b6ztrLyj6cEBd+0ERUX7A//QPzIc
Rrsxd9uqchgh3DuOsLeTxdh4LbQg0ndf6Gxj9DvYxdC9ebtnEMYSMglFstUoqua6Td4TGTY/407O
s1WqawQ33/U4rWHkNXcYz9hCTJVXMB6qQwhfTSlkhWF0o0WjrQjSwR6QqFSy8bhsPdw4iVf5dS3N
x7XPOZNMxmjqV3HKNx03YDGseGfAoSl/FXulJbyOXMPYBd92p4yTxsjkeG9IB3o2/xwL6igt08wX
Tcvce7iH8pniWdL5GMhSViyYe2cQ1W6vSzw9v+feFZffR1gUFDHyim5w3g8cBaCIWa19ILiwaAdu
b6n81I0AnfZdb3mkB0z3stwacoCHR60ErmKUzz+kmcujKl3IFRGnvRqnD2Q1VuOVFHtgTrQXZY2e
/rGn7NpHR/KwSjwbXvwdNm4ZBzvmwWjdKzzHmPBZE8d8FlDuXlDCmVnGYbdpibNYW2dSE/x1XW96
SKfd469VFYU9HD4jVjKVe6BLZAGPx88cL/gXMiFoZXE5O60r7lc1wRQIZUJEQgnof6oxREzecbvq
5W3RwFwXzPWuNT5REd8tkTOl2AIO0cfhpVev5PpKG96MbwReMKi5tD/DyDDpKAMlpeTArSPyEHwf
kETmuQOVOazMT9zjEaBP3OC4EPVHa2o8sHIDsz03LhPBgyr2Uhiisy5ytBNRe609qQMMc1Z7NXs5
pqSoNb5tmpjmdWxTA9Ybd94QoDdbbUKK8NDOJg6kOZ7rR8fVc7OwtPEdA4v0pGNcUe8QbJ8CoK51
13Y4MpN9+h5Ni4sC5QWV1zA9UPAIL6ZSVhEgEN/b8xrKr0nKwhOpVqGsV+4oaGmWgO2K/NuaAzBT
ULMT7/V4xvn0iKW1N3UG0UyFCRe84BGLWWc1NKcduQCabtvyCt/3+ztToYv2fvLgJi2pITuaDCJg
B30ZFk9gbLVHiHtlQgzALlPIk1aQJPtNz+Db97BQA0E8LctVFdOUOXEj6kIVe2J2E9mkattHbS6f
tO9ZL4e8U4hne+GiHEGe2NfyFspd+RSpx9ADYbsHhKawavcgjMmc9DgPDCGzpaPWozHxzBmI5dsi
WuBc7+JJBzSoszNzoWUtesaOJNIZL+etqCxYWmU+u8KZjbQ8ViJwUXc8A6Qh7cWWcXGff6bDWZi4
T19tqtf/MkQJGuWqadxj/cGb/TnIyRMFmyOIaRwMkpufBaQU+HpQLKZWgcWV2CVDjLQTlGLj/wWn
7tV9s5dx6XdPC37UTfVGMp+QgWmwLlRXXtZLqOEUk0rk/F8sfN58cMLyUcz4nCMQczYdR4+U1PFR
HbpfALE7YT/S3PyB59f/PbK3IM8vp+5SSQ4TtjClRLjH/v7J0Y3v5mM+AfTiJFrF7S0iINRTFf3Q
BXQGCI00m/g7HZh3tmGHme8H2Fde7SeFaPCGAkWXPo3mBR4wla/Ev6I2AtWFSUa5GVcDTpoHZEDp
dEm0FwFF5kZhSB275VKzTy9RYh3qA9CNAEJSZQouovd9SJzxQrtvAyCIW2ASt9v/zkHbLwT1r+Hk
KQuR0MV5Ya9BvxjhSbzxRDyWB2e7VQmSLNMj7p87BZC9re8QdhHKgPYX0quINqhyeeuCN+bSdiZW
jQmm51hfHkA0/Y1/6y8iqL8ZATcu4t/5x0QIyPHrdiBMUJxu1BBnQWABlExCqiedH/tiMiFdyme1
3GGKyYVUgdNowoLN+hWFpLx6f2lw3EAVN4XkfVuFAB+fpVd5Af/sR85jN+PAR1hjzSKM8GqP1a43
e+C9K4YdzktTbUiVunt6MdwfE1jDFtKyIF8L76kTZDwBWcJR8LyQdU/W1OCLubdd2UFlUCqNzNXP
gBn3fz2W4kXH5ioOniqT+5zV47QePxv2LMInNGDMQE79US4EMa9Y7O+plPwNyMv/+G4w92n8CUGO
/NM4Y9BxWh/Xig1+E557LTXRZZ0yo0ml4iIyGmFqYN0LW2BPi+qgEfrGnxTbLegDk2FjIRto3YHO
9d7QqmD7YdhhOOoz5PfDrRiFq1FWBNpKC0vINBQWgiE9D6eHzrmgk2nsVVy3HD164INstKjQM/xR
0DbhYpaEas+4QA/INpWJvXhuz9x6UH2RGzPwdJ+PRHL6tWt2i3/1/pYenvx7wfNVuXW62nY106Ia
s89oaiC8PTzDezxhhELInvnY24Z2XFoT5oF+//Ua2jbRSfMQplwAV7HXFux80Xk9s7JlFyEZ24or
48zl7QfHEOilvU0Kw7cpqEs1Z0EuQrMk3Vl0kWOMBBWaLIDl7PI9BCW2vOBuu56vFaan1uOLnNPS
ZrifjL835efgVIzocr/f+BLuyVNLoFV5tmR6peuBOGZVPAPPIgc5RWMs6v8PE8i91MeXebTa53At
jWxDjtCfk83jsyfEObVoqSwSstOv22tVLBoCiYZydmPcR0JPw3H5SqxoHpyqX74I5+zdFMfqkAHX
O2lLJXfQyWVqsuPoRchBHMComKiTm9wZaZuyVLJimjRWJGWwEuuPGFfVka/AYntmcfbsPz6X/DFu
MXw7EDFVHOcQov21Chx93rTIS8Jc3kxtUxFSCJwZU4U/W9ommiYxJlTNmoUvSc1IWssNzQ3pJpTB
d6A5rpyW5yJmqKBFGQBk0d8JIe9M1QwK3B1ejhhyZw1dWGbKC0B1oBuquUsfCdTJOWOROOnkHGwi
pcg31W/XmyHnj9PWywKFZVT4W23fhlX+/P/lFUWwJacXDzkRl0vDqPwCVXjUp0lY/zt5VsPWzIfz
TZ/pQSTSPUAvbboAyJhw+ECBWcZUT2RQB6ej0kpDNzl/HPcmJuUSOOO52qRH0vWABtdXR5j9DUom
ZrY5ebmDNJMP1CZKVTOrvv+GCfqh3ieeT01quZE+rRyMYoKlF4sOCnQbf8Ji+7eqaO3DoDbFhck/
3PU5Y99jhyfY3e/tbXeBaK313vnjjp5AHCQUc3LfSUH6bFDYTaWUKFRFFZtuV+iEk/FX6YmRuy/f
wp9Avpk8Zb35AdM3r1Ew212JY3Z8eiZh9JVkGjYxBK9C2sEOPblws50I+CA9wkIt9fx9JwzHHwC9
3sy4GExcPtlmotBa+zWpdTHw/yBqeDGtcTp5fi0JYexHCkGtsRlOBaHdhMedltq99ABKVw3FR4uL
Ivz/pCQyBoNK7PvE84vl4o7pgPiFfO3LszK9bvB1wNR8xUbgP2ghByRX/C8Di9I5zTa30XhN2+pG
tTSG7yM/cHfuFwG8e4bbrB1vz4c1FiL+Q8y0cnerE2Xxgrx3+8OTXdGG3Yfc+UA8ytKT27qdI5z+
+vIC2Omuu7qTFRt4Z6dhwKC3sfkYVoiRrPJlr3FTU1X9eKuVJgWgrquSZPkGsvRsDhZoGJrIp2Fv
7Mt+G83JasmuUwQWr3RcyZNAuDXrVnMHi5OANQzMaLupa6YpNR+5qarFiMVZQaZHz2plUQk7/mTe
rnMoNztmzKB+G/d7MmPihWRXkyefr6wRL4CWOypKedRAu7M6crvr3IbQrvXDKtTuqKFG02ZSGtJ/
RCbRSjtV0f99gfuaTXaD4BZ3zE/1eyf5r4t196PaVjlUm6AkZ61ULN5CKJl6fgjPaiuAdZeG/wv8
FTz2LwjbYaaXqjq9sBgMg1PYXCUcNTUbe9el9ZLOkFNjD7vNOZ6zjEc6iivZZ05jKUY8vVWFLvX3
kvA7wPccNMlhJWz+dODIr/BlLBxzafWBU7EYGOAbrc2uB7VgDak19Y2sXJgCZLvn1sVF0Z9lZOsw
gPFG3wlD3bkJw520Jf0hobzbRIHroUQ7JtFnY58yHurnkV/Ca6bBfQjFVHvSu1rninSkyS1r/3f3
DBEW0EsjlRb5ICamV6IOEieCsnGB5RMm8PQ69SsmqAf9//HCSFV5nA6yASkoqJPKEeUQwzhZK+QG
8yO12oZUWgHof2SKbGRO2S+rSIf9BRBciyeoqyemIzvGuSCpOmBBhh4gB2RsvShMn2VsiKNBmD+M
WYdPZfZrDR9GBcDRxD7OtDVESBDJnJHsQTQBZaDUKS6SuywwfqBbTb8VTqifreNTyFh/oCi1wWb/
n2yjsaTfpwF6tNZ3z9RLQkfHcT18jZUWlpIWAwCnHvJH4N+kqC3jNDi1MmWEL63AguX+jKqnhrq/
BQCvTIcZ9eEyCMJvQcGybLTiTlwLIMF4ZTabIzX57404/qcleIOtlpuTFVf259Whz95BklpBXkyu
8EIIcpF+wPcW4NwqtXG3r9jixQNv4U6yRxlguhAEHE7xJApJx40NgwSxhif/n0q9ab8A9KhJv9LE
TQQ4k/epR270vBhyhKdVdmsfnd2VvdGippfdZS/phf1f23tcowq0Kn3gQ6/akUZX9UiX5hlTw4q5
LkBYJIUDkDubHylIXFPvq+v3Ts0KR/le75csEqNPE22qk0mL4tEfQ6oadlXZIdoyUZk66lZfBsrZ
gXhykTBmj7IDhMaoejjrBbJBTKEMUzMRf6moW8tTxBxRmkZBwyMg6R7a52acF2F3+wt/TOzxlaUb
8dhFzCwbbbZak4OUK0C9SsgKqGWx+u1mCL15aOokfpOP836BOyHlSWfAINcAGGp97tRYlSH2HsI8
VHktkV5wDaXtI1FaL27UF3UTsmt9xm5zTlrFXjLDzQklL9551+QpPyZ6pp7whoPnle9rrwVCM8rD
sf5oWKLS3hlHE7uF0GEEkLDKGHh4EwiofWuNj4EtaTAaLglvSmmVyozAAS0ydJNHvNH8zQJ6a8TE
ZGCdrLvzIcnPO6ivqAg7KLofBmcasqDtAro583SpNz2IWgRno4jso9v9anWdY5zImUe5WYSCeWCm
H3Ktste4jek/NrQf6FYdejp4hDdu2CUO2zpBPd8fUDkUXeWnwb9fgYqnF8nOscDNsnjIvfkC7ZFb
9bRn0f3El5SvbomX8/atruGNKC6T1p5q5wLUxXTOOFQfFt9tSdpJAJJPhPdZdZ4D/d6Wz/X8WJbL
8IHpEXUfNxB5JXCcyhelOH6qVkcz+jQ9kZ32W2dR7jVb63aaU+2mvyZsdeQrVppY8Ab+W8UJRxOm
9qRDBGb1WLgZbDVYkkhO5+z5XbaOOX+161YACU3KAcgxPquFjFFghH88ZJOnW3AZW8hQAO4isSDV
sbr7woTuxw1HhHPGIt93QbH5Ua03+k4wkr7xMF+dYLm2LuylfIy8n4+Y8pcOg3QFoBJXKhTi0yaQ
17yDbZOgQ4tksNH40xrt281oJS07w+H1nW8gZPqu/TY6Bh8HlOP4iFAhrTHnDLu6/AvuzZ3Ky3AE
klbIgQg8tInikePozlHvVwTLC530y0/4tJNC8AbVBYk4gbQqg3wbhxkYWbUqoVAL8wV8cRzaU/wl
8hF/DDsYKwVzrpkLvTAXzCV+e9GAcl9MucyPkff6+dh/9LSmIx7gABt6np5ycXcEwhIhqxxRK38R
VbXECtX/Qm17APA1zJh+0a4VsweJiDhDOg5ZMjki9S90OBKwg1Pwvg7+WyNLvbinawJddJmf4wlD
p9qtzTLs1WBPs0cyNG0RjX50kc8mP1n3uBRyrHU6q/Z51QjadX+KxkROYDBzfv5XXsOqZJSwZ1hR
1FSQ/YNNbCEaP2e2cBvvhTbZfq+r8esHuqaXL7oM065ldEhb9J7IBHX43kY30eT+9TQos0iMsBPT
gWL6SWycdTmZTpj+cCE+aVFN6J4gXdzC0i4CboOVhZA24V1jFiPGAoDOhW01z0k6MMye8GaMTMfl
aT+r+B91PH/qva11y/4anInsVwK2N+ldtsyl2rAY8BfS/dK+WIzUpHcHYMtkGnpfzsNv1q/U0ZFe
PmqZgHImWpMhVSwkqsUK7x/YhKRNFEbnYjt/3DmhdBstRb6ZDaVftPSj90YJsnZGOlcwXK+Nfu2B
CLcNCpKwD8ZDnG0DCKTBes0fRnIFN3/5fbbkGMGPqfsxu1piWK+nLKhoLWl8MaHKGsAx8CEGng+7
y9VBTfj1jBIakDhmDQBeyrQ7EGjkmMr4kwhO/d8FxmCwYw6tWWPpfDJABlWr3VyFQ+kHKoWchIY0
5kFjzWgIPc75c+fP+zXOIaF94TBQHGQTzLffJc4qDcBENvPxk03H0iqhb2jQDklBhY0lHagC69B4
ytLkIWYkygQB9QshyKPaRzHWoGj34aUOBlCriAGFkrh66SpIHxliAPn9UvjuP1HGtjUCCYOFKsmz
gF8IeA77DE/IVqbRNSb5RjCtpn9fgQt7PXHSGTdHeGn6xNU9NxsQruK7PuBCUB1/D7qOu2kPhThk
1pz71/866Vr31PHfNK2j7wZowGJHViAcFNHe5uhzhCPAff5jc7kMmWmARQsnowQ3U4A/3NUGyPkL
/fTbqNuFsANB7k+r3jcWojYTRhsmAChkoNf+0UzywXI2Hkw30v9LL1h8XHQQYYH1wDVhgnYf63Zt
jZpm+1dVz0s7nhmmaKIjR5TtUJq+PD90XueYwwlXlM8Fp6/taez/UybfdVsGlF9QRwBgudDJ0XEb
JOkHdhkzTKMOCpW6RhyXI+L6v5yaVsyKgr+xqKv5BdCUU7BhYsutgxqm8DgZ3TtvTOxYz0rGIqxk
7hwcM+g0K0KGhKgiL6u18iGeMeJmaVtaABdFygdatqnaVYY6iY0dID+3J/UynHw0vCaxsYkjpZBg
WklsHPnTfCeUYCiIkYToTqzTHj0gjW3+I9WYdVcm0M0CVRR+aEtUseMOIAly6XmMWf2VetAL9AGu
lisfcWsCTmnX45ERwZmGPWZsbC1yZExJXhMyj1L8OxNE+mz4858GWjr6o5dW+ewNHAq6peN/bJPg
4WoyoN+BtSwjyGt4c4bn5n2AjG6DdsNBISJTmeYOiUrvHBnx8hwmFvMoZaciWBqO+Gd9nTsOZil9
CpE3iqiJ7WJ5IWRNx1jCeLx3heAYNzvQMJRQr4GRb0WHQuHGKPlaB097RmPy4z8pK/udufK1K5vy
S161mxuOmZMqe5rBsBaPA6McMjgD93d6kHWCFb5eF2NA28StuMfzbRY+O3GfSzgmxxz2lqRDHNl+
FHRXtpm33Pg8A5u6eHAuc55QoYMGW3qBLQeBtoPQSI4FEsL030J/t819f+6lUmEzVCXVxMDV1d6o
zGEjuct/ntoPui/4zCqP0iepRC5JIUXHz1mc/cb1EwUIOX9bmKVk5FoZPKX9un05QOfnCjIeWTEQ
S7Dv3LkzqTf/uTwCl8MPtNrQxxa2IcMm2DPjfa8Czk7d9OcLP5/jMVvRRsaiV9M6uWBeXcuf9yz2
vRsfxGIvxljqtjhPMXfmuuxniBsEXd/Oy1UxPHWt0iV8Q5mvbUbbwPTFzUe/q2lWuV98PlXIGPn3
V4tnRYLfMO/96MZK2hHbu1s45FJa1/ijW1wRSykfHxfsMTYGo6ehrhkZyH2S8Qxy7j/avXbBE9BS
pTUcp93jQ5x+zhmnNQdLmgpi147J6Q5iBopUr5G5uOlX+8fzRlw+BcTO0UpeSMizCqFanv7GKJRo
JTB2JaWGO0jVGW6F0gvAQUBqRR8LPcYIfUqMg6ckxp7w7N0Qh6wub2YxNMa8cXcORuFHdxEQYiuD
RvKSFur4RxyAyoKpcFg6HES++VBv0C8ZO7cSjgFWDxGJSxh3CJ98Rfrn6b6F1fHSAMm2VnhEeg2V
jrjixmsLholyKge922pam2AtfGYu5TV3Fjc6Yvu3UGDG6Ihwkhhz62phtFUTVEH66okjP6hvsyJT
SQml8OFRq3S5Wog53tMYTjMHxq0pMHUJncyYaMkW7oInkkdAdwCdFJcgIgdmPQlEK0RVKkPDWbEN
ABB9oNIJu8/PBk/Q4ZSZI3MtZGZcEtPXryzWyKQxmrx23WbUZ7iAnCOIIYUhvnRWLFHGY1GlDkSz
NPgyqV0ZhvhMHAYsk/+X7fDOa0WhDuRcv4MN8AEzjdF4IKOYQ7CeoShTgSNfz9WwjBLDaEYzQ0Vr
li6dS4tyqmn5wbZZc7RfGzpC5K9eWegbKdPhnFZMvlp+pvTvitYUf1J4SkoAkggyzh+w7vGqM8x0
YjUeOBLacsXCXBeotATbdqqL9bea1d1cnfeU8qnBYrdIJmVfZWfJdILY4fdl+Mn+Liqrgw32zzXv
l4TPj1cmozErmFmuJPCFlzTKMnUfEk76PPt1jhhXa2iBoRWDKAmv9ccaBgirkShxL7l423LgKWwK
7l6sQm8HUnCqy4ENSBtCKJZ1NDpPG+MgW7VsgZmXRzR7YEWg5im9/Lyzzyjf0mgq71DkcHCmkG1t
tEVHnghKW1ZADLDZwIyOUXAkq9Y7jhOc6Nuolz5cnZqR94lnJmmLFqtnHHi7+6gpHyf8oIRUNAcM
qg+o4iLfSMQFKLN8tCSxB3R6izsMQzv8AAifznnlCW7bVsqJQReg+9SgPvB2Se/Eg3X81vtYS5Vq
CfoAHSixAqOtrkMy3dPJ+mHj3wI/lUWF2bqb4yfhiJQijUXTYALuu2Y2Jx7kQyyLFQzyzilSRlKn
89ZIDmmUI0b9andQW/NBB1aHpp8g38hnL7SEZN5KgzAXWcBVg8TiS1BY33iUTxhzezWGZ1XNPNmf
8V77OPGsyLT+Sa72Zc++FN7ffG+9L2G7gHb5GxxzgWdUzo1W1L+gEhlZcJzYZU5LENNS4omDFGZ7
TfgG1z2qJZKcaVSSrooN5A3Jj6fevYVP6LRXBuU+2/nStMvkE6ZMM1Nfbv2X1YCTarjX3WfwbLPv
2KZfBSOGCrVme9i0NHRTAK5mySTc69gHK5a88GiIrXxnPbo+FOsVJStIoae9l/LJ8I/h4T5eC4T3
4g6QWFkeMCTcjxROJHVuc8wT/Qiy1VKHqfhvUAft/WwyVnBi5L1U/gitGrvgAHaJJq2ZN7wx3mYO
9DY0Q3YgSjqALoOgCjhKIOd8675cYJdBts3Ae2t4JiW8x1U0MqWqcjfp+n/7UfnuZv0974u4Ydrc
eb9qzSEBZj8OlpkjuLFSvBIjluya8miuwPZK/TBkIcIkQRzYVDjOBE/l3f+W3f5wb5d7P5rS2XJC
YIknDijxGwRkAWs/e4GeMxsAREOcgtQdlGgcFup25qUz35bPqbOro3/LvEe4McOjq7RdhquoU3jV
c3FONrSGV+xB+6mH+H/1T+d4wnuO/dYVQgIOJOlutvJWYZH5JbfL2BhOCevBi09MC8KOP9n13PiA
qs3N9TC0013qd1SA/huhdlRVZoypS7TrrC6jn3vwK7eeZGwuyi2KZolA0Is7fOT1KT/6Xi0parVB
hrvpN6kmlPzRQET5cdkuI9OS+VvsUGdJz9pewbN+432HmmBlocCkBhN1qeN+9027lGEeUflsO0hG
Sd5+CP4hA80A5uxD3rNpwLiPGL2z8e7p/8qbAdv7ggWlEMWrUtTr+WEhNCBAOhwLytHhlzHTMMF/
9RxmrFpyqRaKZGHze02XjyTh/nEOK2WCB/tYaG5GMV7rBCX0MgNyjDS3mkmCjYLlt27S+rE0kBxK
Drb+enUSo8C8/85AoIqQ5uzr6IcMXExcpRnEsfa7yLdhnmUTutJlwAYF0QMYFxs7uABYql+0g4nx
cgW9/+eSjClcIcQEHStrPMAVj27f+ZN33bhrL5LZRxMbxMgVjZHVg/h1SQYm0aUvMLuUyjaIwfvP
SdpjuGsaM+Xv7QDEPF2eqrI/m5ZHTnJOeVM0SQX28rmZUSpV9tKd2RtOjfqVgwfhHwJ9oTSLDt11
IBr1e4c2IjgkAdNunFCwusuM+nPUThwV/z+CRuighsJ2Q2vA2nk3aMMGggr1lD5fd30oFzK7hwZz
iTel+erUGuBl1Q8Vfx4SjokDLu/NteK3fIeASQvicgAVjhQeDvhh2R5k9HPCJzfzv7AaIxUOFsSD
IqeUp76ZJgIWBUYfVmthr3TmCqk4ev6PSjPlfPQ21mGd6N7OkGz9jm8j/sR+rXDdLW7rWDKm4quO
WwqDajITsEuPmwo2SXh4xaJzahlpt4oAYcd/FjspF6OKKIyToooRn5+W5YUPlCKimmGD1lOpfpF9
VyEJzfoCirV2V8VeTdhbUmTSfQVXCTRKWqwlcHlDcdgtflELcZPexF5Om2id2ax26mJJ2evM4Ygd
SgVJ9vhePa7TKrZ2n7X5Mb+vrsiCTTVmPECXdxmoEJRvMwbwu5m//vVQxA5vsuCTYPorbdQDzQMh
N5c9d7sRaNumj+DefBJtF94y6TzCCrYNg5JOuBJfheNF0rjIxQI7YXyhbdEn+SzImUYm0lJBHNdq
X42kyRLdUGRTbEEF925+gTIejMkPAn3jt9ySSaw0qro2PvOmwT0IstXHTHlpFlDWrP/YL0SmOo8Y
7kK4pU8pgLrm7w2I/t8BdVQQtYWufpwPxrF0eqbtyGwsIEt7GI2YKVAIwLBlyHLlYv6VES3gMsv9
23LGejAPjAgRcHGtKCbmJ8lQQRAOvr2PNrFYI8r7P7B6UN6214Cs+cIlJiSpiJcvM58xNIkA9QtZ
EYD9S7VZ84dNcrj5DzMWzOfqkxXeYpnHB/mhqWxEekwVXxkakMWf936aiAv07Ujs9wXQ0wxQ5hNZ
VG7e+vXZTCAAcRI8RzZT1yptCRm2URBHOIHIxGtV+8q7DxJaikM/n7NdT9eFpA2GxN89aMN+lvJF
aoi1VMfuq3syM20WvJZNFVmRZimkPl6WRjhilw0TiI6z6h35deI3wr07BXBfO+GinszUpPMFaDR4
oct6pmSUJFMpuJnC10wjtLP2GiO+4coWRvKWZ2J8Mx0OfoyRlDd/1gS/r1jqQfHmuEr4EFILrqLp
JBZDjOy1LqLWlgy9K8pqfjaVRwykxF8pfSDEe9Yuy8f4TTsZa/Wwx4mkyDKMh3JJ9ZcOLkNPUjzR
5fxE5C2hPaiwb1n9D7HUy9u4PyMfKV8uoUGPC3ZTL8E4EAYjR6GWM+iQHEo4HYZNmX6qMqGR/Lq/
hSYl3O7tjF01Bho4+wXW8omZl3TtpO830cCzhWp1VZa87StfCqNKZOwpLTmVO945Y/JlS+UzfpZu
uMn1xXtlmSTJoseBm+/A42SIuAOHP9mIyHp7PRFocgKMDdjrUgsL+X0Q4yaZjSYOjMz2AmsqioH5
gPAX7SHfTGDRtOyjUcNoa/5PVRSCOgMLc50n42gGLKnfATTR1QuW5xmXlfScLcQWy8t5yEb/sOl2
W63d4IjLh6LkvDRKJWKC3cLmx7whU0ku4ZiXx+jQaJGcj4VYk3XNkHrRvIPSvu7KLTvltQmlsDBk
hMZBDBGzTg5q0HbPVXeNBkyqNlL1Nj4q3qKFx3iVAF5uspPFeCBaK/B63r6h4SCGR7c6TYgG81Mi
+hMhJg1SEGaGwpnRJnLYU4DYFzCk9b7JEnrWphf7wELiM3tEA1HQPf8ox/tjKrB8QpW0kCoJ7zmy
kARaMdQ8/WETok/Ik/ekSnhT7oVqKlftbgNlZSSSAlxx3oxII6OPrqsFH8nYauFPEXgg5Qrz/WO+
sxCcGE8OPRHwCsXEcAsZlZ/6k0jbAhpNhtgQH1wdsx9NAwRSgfLKPA6oqGMY+HLOdbIzh/+oj8S0
jXwzJSrisVXuIvueCDjAWmROiD1vwLdbvmbYLpQC+Z0go3rWHlSVbIjj2ex2IjkV8L7fb0Z68WPD
q1UPs0JOAIYNj0L/wr5i06nQQ7CCM80Cr6Gv7+ylKk4jWuLg5ltAdfL2mHbhArlXCQslwViJV5xw
QoDSkb+Iln0XmeZbvngbn5RLPAyuBeRWRadvlA9bP8ypf/mHmH88EhW/ZUOWbhW8LE4tiOFVbyAt
FQH5P7fK6kDxZQAvDeEytKjcQ7OBec+a/D95eeycpaA5rnQ8BGUEsLnnkLRaflKwsDh9Zf55NfsP
Nlnz0UT1Ba+L0njA9Dtak80fv3ohUVxF9Cjqpy4R5PFFac+wkFm8B3485x/N6cQfMT2UFypQNoEm
bspRWsmk4s4RknkQCCKJiFQYC2eFNDE3fHHysTUgq5D0jdSqu4AREDEWwb/ki76cso/Im0tlzliF
HmavhglyB/3ELEch9pY/cDD4XJehwXPJyJFjNE2Cyig6Ixe9OXsstq3akgui+ah7V61quQV5VCjY
+D9jvfMIFMlhrDweHi5QJ2ID3peV6igfBEDJz+FxMON7W0Azy4t1BIKSGkuyfnQGwpRoF3Uyibvg
eXRaQW5Eqi2GlmaAzkJMCGJJ+atz5hR8XTHBzvTazOXJXrG4y11u91RyjFrpFXEI8L91ew1RZoeg
GLkRhEKGNxDtUCSviTGjFH3uAYVYaPojSOfVBJ9nADmby/JBHyGFlSigRIioYYf5mzTTGtDynnCZ
Yso+i7xaJSfhVt0Osn091cXhRixWM/HitAkawyDMnAGUm5Jg/9qwz8OTFnzX3F8gIwsNENGHi+/O
YZClXO/AkCjgj79soQWsWYvUEEnM2xOo8A6dAQL384bYNhY7J1gOYKUniAqxte+sCilTKgEeSdkv
M1ScdQxVSVJznB+kfblo5xFhCkLM27M6b+GyzglHfogpxZGL9eUhzI2y6F8mO5IoYroxOwMgX9ph
nYDe/NbETmXc+Sr3eZPQ1HPpoZKa5PcVLdmhj5nBEG7f7uTdEv3CIYDPhIEC32hKbSsc8s4RmnCH
EvVTQqzveBJ2AoVaDxXmu47i/ZpsQf3kv0oRp4aECnKObugBxmHZGKRdnycVyCyYkqU7s0CnsvQH
AJJbpOuDgTA4GmH9Jm3vDqMiJ8ey8MTUxAHXxqoixT9XtxhUZ+bsoc9YcZeP/ImSWjMs1Z2NWW+1
N2DvHBhzCMi3x5tcUcaWd6s1P3+CYyNC85gX5SivUTcUE71CrxQDcfQmyEngDjRyc54VtHku/qgr
inMz12Xq8FVRsPuJFc2qBpkJJSAugzDpwSFXeUwCH5meOilNb7YX3aEy7//ZYpifct2G2FEu6Ynn
E8JhF33BWhUhCT4/Yu+JxaB/IBGwAzprBh3w05vVqjbwdZ9zn+m3zMrJs5ojLfq1Ce0u3xTIE119
L6d+X0k9lJ1VMx2KtFjbJHVxdfJUyp2KsYRBPp3xWrIMs8TEwOzMBDJFpumUCHnlqNQ5avmkv688
ZiJk67N3NeFreF/CW52/tRsepnOBKtFKXO9mfdHDIvPwMdq290fuD20zZRrqtnAEJcIly3s3AT4K
9aArw15pc7etKkafk5wWSB8X1NFgVUygoxVQTx9lL2gJGAq+A13nszPBdTObnSFdGn/leOsJ7PzR
edde1SLuIP6cM13DH+uNqW9fAvMQXv836A3NyMenxYheYoZ6979kCZRkXGPJBXQAKF1hhDRy4LJB
VLot3pgXKY4yMW+ialXOdeZgvpQen8psCOCk79cjzDMvc2ebpGrcCizMAjQJhpGE3+Kgp1hr+XWn
rzfoqOak08Xkdm9l3d1IpXDjBf1vGBJIOnzTxPmzGiGaeAyqKu3TiPw53mjFn4+bkqxQ5HI6vFE9
YYq/3mPV7q86uSGfUFWE4iIYvzdjV/ZV+iZaA/URfyzTnsCKmfxLXK7/f2yPODfbflrwDce2Jhea
9jt9H2myhr7nWf5Yg2llLRCl43kvAM8Lf8qhDVGKjCKuKbQcDDmVZNry26ctZRPMCYBAeeuO8XM/
rV7VsCHHwcT1kzVNCQslER0RX/H4N3E8p3vmlIJHLu4v/Yzr7W6uUSwmThMejaByFubi1pypAZKe
fTbE1eoE/OamdDyeTSxdaF6k5+WWjVd4OOp9kAnTdOS5SZXlUs3h6Z5UW1wlWAKURHh0qvGVdla4
bfyeoLiWPsvdI81DiN+mIEwTQU32xB8yy97JD06hc+PlXsLzLr4Ci65OY4YhEdKEn/NqgHAmJWyd
9K6xoIVJJILC6jT/UOaf33dJtOLqAlGBzLIWmsrKnMFELyS+2xrqt3U04YpsvUcDh2mNYE5D5drZ
gyaaBFsHnjXFKJwb2yBPEMMwD6ylu1iqAPeWeFxTXdJenBGxdHy77rhTN0xfxWi1lC7OYLpStbdm
LhYHKin/6FQZapS8yZl7MdSZ3ZEAjQzo4hHSQyUELFN0a/oWR+syumEcKGqe2+TVHzFC25ZVO66+
rKOmOj/n6uzhQ4Bk1LheYAA5ompADun0yBi0gnxtVkLS0YsmFJMK1OSaVunVA7bi0ZwfpipMOAEO
9CR3MIcxSX9EX2Z1BouRFQWgFCGe7WIzNL7udTkHUowxn8LVoOkxBNnvgTyhLX65jsFZ11UonkhG
XtjocE2zxY4WV3gqyyuacQjHsgDemtgUP2T/bWVPCukYIf3+pOXagO/rfGEmpUYU0xBf+MyCQbnh
xxAdNXnwZi4LW4tphZWkxRcvybpiUq1th1ya2pB7wo+twXJRthU1AfmQMG1RNq4ngPnQQS5mypV8
4eJcEYT0LLa1z8FC9wFnt8mswUJFYnYvb0j5EVyJ60u7sjxmNJ+fVnhKTsrmNrnB2LZH+9Yc0fMB
jADzsCCLD5aSFwD6a3XNFnGKDDIN9PFWayb2Ya6cIa0/9Z4p2V7QXi+tCOZCn40l0L/oTGlmfv6z
N3XkEzYlX+nFtHM6JV/Xu5qmLVruTc/qWdZ5AmxG6rg1Frqt5aVrNCqrjOQY69x8uONlgBzUzK5a
ScMSTikLc7+jkYrBbxub74cbX4VjhxseuBGvrPdo/taWHC3DgYVuyKBuw4i/y6zqU/kaPfL3RLIS
DdxHfbvFf5aS46gKXRTszzu8NsqXAaLOxU2TCte6we4G7wjkPiXZHBj1GGbWau23ngPlT5GYImwV
972gfryo52zBjOPrFxfi1t7YON01H708+JQU52Wn1R6gs/Fjjb0jafBIaH9ZmfRkA1gY060yhuFd
x97QIWwksv7NG8mGx4aFowNwOWq9jI831YnEk1NkjBu0dXn6oT3k3LwosY/e8j7vJ3TS1Sy6bqeq
G8IUQH2Bb9fQjkJ9rs0LQ0tvQxxEDyai1O29BJdRMf2aUy32QS5AUD1uX8YnmT3GfjM7GL6Hu9OB
nZryG9Il/obpmJds3kyR3MD9s12DtgXeKgVfd2JE06l3TX/hcBO5FlYRKWY6+GhXWp2uzE6e72pp
aDUmE4n/WcHs5GRagO3KZQvYju0eHyKedYSrHITplFFb/Qd9F64svvyPGf1tBj47j1iAPmBxj5nE
M3R6KQRXiymdzHTPVIZMOwA7YiC6E/YaXKXJQ3qBa1k5fC2EqeyOH2Tkl2yGjt3X4WPIa7ppsW4T
l94oXpAX6wCfJTZGaPcQ9rSvKrC2E2V2ipjNB7RS9CI49ycslndP9ReEe5uQ8tcRKEYltbbhLyVt
MdbkN39l26+TKgb770sW0IeavfNg0G7e4XpyFyezmfnEdnIYjsjgHGpogXBfAAVeFisEuWuLo0ap
k2c/TRVneIOOU748dcyJdKN5TdoIxWra3FDK/TzrmZ5AJqqphNh8YhrG7/Z3dKL6RyEUhEyv47vv
mRW+w9/DS9sUVUdOBQ8J+KT+3jRWSds6icXXhbteZI6TK540pEBkje8AknzGCWb0V2/hhsQ+3BX0
+6bccKB6ZPrwjMuJAHh887c1rjrwGCSSTHLcEANTuTdo4OXvIdOeMkVxb8j5GAfTOzERWA+X2dY2
eOaqJnfe5B2C7HHcxzxIbu3ub7S6qpBiAFwW4YtcFlZGtTJnZ4DKxzZDEsMMtV/vKytZ1b5+t/zt
ZVfl6MSGdbQspKTg0tU14sa52I+iPXzFdZERVUT+mo0xPUzdygltdha7hrjt4BKc+isPgTgLO8Uv
36P3CZ6vLFxnafWQGuk1yEzXlZhlahKVv6dG61E39GvHNQD123zfuEshEr6nwhpBczbLRBCv0ny1
gON2aOmmG92BuCsxMWsvj72tbdwHCLonbyLtVwRHdeU5pg/WwPm1xf9wOpkT3laTtVvaA5A8gqER
20+pBBzJnrUwUft/RtIXSGRZc/z70b/Y2Wa5GTJO1++bzyIIFPZNrari7xL/9/w/33/ppk+qJeB8
h5a4GE/kkUB5WhoED69SMGnpKMD7sso5HkGhGan0vnW+CHCzNgd9LRfeEjgBSefz1SuPcUJ1C8lW
3VX1iDNlS+cJIb0CA9UZ7ulGNmx9WHG1aQmm2kbZEennxsIFe2qOlzm57O0v7kUF88BLQQt0Y3qR
O9DtGVEd3JNwvvje9cKCEOOaKIhirYxNudqOYnICSgxJBNuuQ3uOBkCYNleEbHDLFDElg11RneTM
xx1MpBGsOSGQAXZJJVbFCSuN63g1bEvjoxugxqADj/5RCABQLl2zN75mhgMd6Fg/NvprEwpbvvxp
KM+pj6nP3OjMAHa9siEQnWQhCRgfwMDsxk3J412B0IKuFScI7csOb4Lc4eITj9oxG006ltMubY7E
+EGsWih5QsD5Skl/hwvJeHsxTqtOGrS+k4EMdPZatoduPEU1GgujbhGMv2dgUKP0tLe5Zhior3Dl
8kftSYBPoMl5pLTPZkqG7PsXydrbHEK3B6Su7h4qkxnJysxgqY3GJOEb9bFE0ZcKPqzBlNP/YH8D
mdEnOP8VHHcooUBQ4Gd/8zPZPmkHsJVpBGHwJKTCrxN7dZfStkuyqmLssWoTbXt1iD0Mu1s+HwvV
AspzeqU7zyG0CM5d2h1gApGMxBeCiTuS2tqt5MUtx48Ps4LyKxBduYqhaHIqhXJK3R7VDohNRegU
Aegqwe3wC/0Djf9HZuX8wAbHOCKTYE66GNAV/eRyhTHuBcrBhJm56w9Ghvsm/m9en9EoTFuVN3A2
QcSpGHAt/Zc1qeHcHqp3X+/ERmL0fUTn8xHUn3UMy+jF6zhvNj7nz4JdZFh0kKphpyMfjJXI2Teh
yrQXyp29tsGISWXksyH0VD66zBau+7XTr9INr6AusszZZ9D1iJxK0+XnWUys4zjlLGoPdNQtQ976
UgCY1vey4cgNIytFp1YnG4HsSeueCfIRjh5r1tn1ocB5IP5Dx/aFKMkjehGhq1YuoxB3bqsdvpSu
nLmw9tiI2qJI0SYjjjHDgKKObiVzSMH+8KS6S0GSOjEhjM6JIIBwz2rsIJHIt7tK3YUD9XpUFsqm
mhZFyfKhl8rtktVVtMp0ulQtbEriN8jC19LniqKKmGF8AKznw5qkmtGRp9h9YDp77jgY2y+Sl7zB
8s60yCQ9vWYDMn67+CD+SbRdeHJRhgbTtTQbsh3LMTjrd1WV8puScV8Z6dO7S06os/UGqGBJFsGC
RJcJt8Q511EJh0djpa2h9p9kmKF1Q0xf88kUOiSX30bEzOZm7z1wfyvtMBLEUolLmhnJJ+oeM+Sc
XgH4yynPPAsO1Lf9IUXJzyIWXpQv8R/DwBzENRh8owBq2LoDiLE5RkwaD58u7MjlrQi/bK/yIbtw
7wnMmNXWM69X0ye4m/9BeWJHbhi2fdO1oAdcKK+xE4mhGhhTxa+/TR1SOiE+TdsbTnSwic8VF9YJ
8k+qPeDrbIu9gXw20sJNAgnWAs1oTlfpe3fobEQDvqH+sHdaXn0wlwu08KCAEEYaEnq+yS48xfgh
GkpxYIccStKHIYOhQOUotYdiVEevHLJtD9LUfWnP28/DlTZqoUhQbp3kuaG+VDHTLBo+kdq7pWQQ
TUvxTicvO/HRQ2iKCKbiUdSDvIwijGK9N5lc2fZE1mdsmzAtrW5G2+/ShkQJJ/M86LaQWf8CoAgG
57QkM+Q/tWxAy3RI5rwrcDFWWHru1TTNktf8kyyHJ0s0xDi9IoHqz7SSZq98l6uGhE2KHt4x8BWK
ds0GcePFdgfG1GXCFNRzgCzc2FDNTecQ1dXezheXZ7uknqMjupcDwc+6ANWy0akh9jCB/2Sq9x4z
wyme+GzxoFej2WR6rbwmXOtq96DKoJl5eVa/7d8Vffi7IOqcWPWXPFUNz79F8wonHrDFHt3yKvi3
79nnHx39SAsqbc6SY7iEjg9iGkxMoqDAA4N+WYgINhzNMvdCQLdnGUlR1iw0cW6oBCQEjUpGf0NU
hqziGU/1600yf/1GAEoZILMetaviwrW7HjPqMm6ej8eFd98/G6R2YlO3RS8GI8n6/Ts+QWdNOjWR
Z3NvqyHzKkduzjwlp9s7XpeiLQry798d0bsawWKkvWcvXneiEchbJq3ZrBiokBfOAsrqSydeW3Iy
pcet+0svY2U55/9tnqb9sJVCwxpG/v4R30Rf0jkRZ0pSBjg7V3P2ym/B+q5B157XeIS0mNR4cz4i
KwnjVWMCNW4qhD/OtwCl4iyAmMeJ71Pe9WQXBLPFH/hINzYNq1dLXbad0MpzqvIvYKIXqdM1hiBA
6DZS7n8X+GkW1kYU/yi1uekeeksDJZGgcBEgkSPqUI2Fm3dJbVOcepSsVf/rQAzPxpvte6Yx7vfs
QP9D7xITbhO5ejEYlwRqo65HkEQF4l280sf3TlsW3yt/rwYXZwxZonHjPiIuRG2IYMD7ceWZtF9z
P4Hk8/oOM7j43yeAwQQOi26hTZP79fgf5CS8A8MqW/JxmnNv6LyOb40DFDiYO7E5Agzcx2aVQ/Q5
D6OeN/g0lXXU+OwsKS5fbhehILL6GXvbSFRVs4jyo9kOe63dUe5oYEkc5EzTp3CRrBcxKXWzv/T+
PlNBV+Ugs8Th4CLa/ltVhTrEePQGUd/ZjmnmDUg0RKMJ1xdbg8lY8HuMRIpDRZS3AnMcC4TMj5GJ
WLcopYG1Srh6FcYG6wUAWVZzA2QoyB9dlqc+3Q21pxXxbC7bVPtIA5nMYbYX3f5FD4HQjZySbQU8
i87yLv7Cf2ObKqNoKd64dDq2fum/6vz0swYOmhnDv3n8bglGJIA0CxM7TLsrM/bEHhtJDIr5vGow
35EPFYW8VnFiGIuOTSuYtbVKeCQx3RJQVn8pTN+4+MFQWbWViuXuI2PgtFgttmtFlUUaduWOeUbC
OVMri4BYWgvU6299GmuJ9Qv71vDfJgkmHdO+S63pvYuIk/58a934oA/2I1paNTLgS/U/ZkLB0+dU
kbl3fMaVs7ihjhifnC0QZAIraIZBYXsychPTWdEvjXMHWd04k/GKpPe+CyIAyfE7bJxXVDzkWM61
yreniOGNwQm/EmltRe047pL5WqjsYweggZSxigzx5/8wVJ7IQiQngQLt2DQK6QoXUg9T6q2E9ecz
fQ1HZt6O5zPZ0x/5oL2ki/bIdFBEPqw68SpCtkoqx5bfcKnf0RF2Mtq36ZSTcq4rDenuiuEycjkI
QVjjerWMP3Y7O+B3VcGOlzfxawweSGJwuJGRCvFHyJYV/RIvlB48+oioQsidtyvSW8q/Kn/d317v
TPtUDZQHDEp9SzwFCxknevsFQN5q/fBBcff5gkjfu+CbPqzwZ97WpTJTYV7EAPbr/KvcsHzENsgg
XWwz1ClkVqNmOBXbYt/0592CGc/+pOf+1IbLFrUDxj/juoUDxJt+Hx2HaNq3UOYLlMqU5fVp9eE3
XZaH+khbvckvR0Aq+czi5LOvAYj/WqOXTB8GFBgs+oQerpXhSMyz+84/PUH2QAvxDnA6wJTAQlMi
TP5PRpRwlTOygGW3jFpGryV0dIt95GZRkvxODURNlpvC1kvbKJsNBtxWelzvmET4qnT3NHTAbuh8
5PJy2o6hnqNBvNDPLcaDYBukhHeaGst2Us9/JZvjSrSamR4LP5GNlPXYJyiz+yJJRchRx2kLy6eA
y8QWKPKfuPPLltLaY5rFJWUd2khkxuKXeGgyL15Z03e5+25+UV6vOkICZ0mkwuUsXwpCcyW6JXwt
fnugRgLgKh2wavTOwE7Gov4Tbt2e8F+Ot50L1Ey7RICFDLS1hanRJEmcpwZ3hYND6Quj5WOosBDu
cijg0JMUmst5JDVSA16tHfd/NVO8wttWlgP8NshHDdwqGlikFNbzrPvcEcxPte9Bqxw7gMwO6sEj
HUh26jtZ+0NlUwxpQ3fre46/n6GbUusWnUNq/72/ZwXC8f22d8chptHfzKg9kkP+t/+bbs3x79X2
91StFNYG33KIr5POQXerpXXz92au2DlQDlLXgrOix34I/tTntMey/Ra04qXz9OyQHi3bXBxZhdB8
HnJ8AlrEuQAJFtk+SUmVgg+6pQY4BOBBXGmnXEaZR5zSb1a4mRYeAUaoJoZcsnrZTfM8nvpNueTK
w7r1j3jm5h/VoZd3EkiP7B8Pq9oEco6sXyj+kloRQIAu4YSYqkOKhl779hnCDXwUTaiPngHymL0T
MJ2GYFDjzngdsoF0pIqu+uoo3FtuXbL+nir5nteEvUgINLB3BvH3VtnVhQmhFPc7MBKe99QFPDyM
oioX+BtLXw/0mER5I3dgZvutAl3SDUhPTAwb4Yh61bPgYGTxS0M9EUJTUnvCRPyrWmO9pvr7mwXy
v2xx4+UVYc9Do662MR6ZN7G5vTvZN6oGc/Ns+w51qgvof6VnuRbyg0muO552x5nyayIzSzKJXpVk
9elZ6pbAmMffKtuuEwOr0nDxrQ/x7asraxgpvS2Tef8T3fO9jPMRk0l8PDyVePIiL9/9mCUQp9AX
SuLxh48g0Hl+mvb5JYo27IZyhw9N9vn8itwWcDYfBeL9ct+4hk4If6iHvhLFKpdr7hO9Na6ryjsW
0JAHrum8uMcFpLnQX8NLiSb6ooQoFUcR1MiaMO1vsoQIUdybdlezVgAgAjJcUYnHKBfsgq6fKXU8
PbNsYILVDZ45HTTIQtu5fPl5T+TbeAU157cTs5Gsw+ga1lth8yHZ8PkOtD/zJkR+ReruT7e49Qvc
5jb47gveKJUymduQ/nCiaJnPyGEUdmm4X7vHnoJKwaku18qQznF8ZZ1VFvZt4G8auCGHqdkMWdgJ
GT0XI+5vr92QJyhXZ2MAFvbUbXXD9NgCQtbNmvTAJjWmVNaN94S3NXQjNWVM4ExbbUtxAzUM1vKV
VvMv0vJk1OoA3RG2HAD7M15GioQ41NV4Qfd7LSbjvuHC8RzXFx6YrkExN3pDRdk3GTgEFiHLJTYC
pYQACgy7JDpGZWc3lrBP8TL9Fb/c+JDHXIkJ56XkNUvVTPRJY+1nu632/TkQsodPN0KiWkNWX7vp
m05zvxSaQ6IVBSr1OSySX9L+MfwYSxGpI/zbp6wjtP7Ow2OAxWQCow+5Pf6TJxPY+oTu8bAYh8Fe
fozXBLlQaeeCcuxEojJWHGGSWJjjS1zTCY5Do8DrXW/DLjfm46SeBYCjW8xYrBOX7ga2TsZOn/g7
42k8UKbmNFeGSoY3hkY4QRXoIeXIO+eNiydqvAfX9kR18FeZFYj0eOASwjjWal1Un8VjoQLF5oZH
3aNhJyhjAbW/bxeQqyFpKh8IgmAQmh/dIkzStYbi9pRfjOpVx7YBSVo0uSYS87zvmhQ7ThZGmlFf
nAKORqshguXof5OQrFxGWtD9HEOfbSB9M5nzlUGpOW7tvh/rzK6+ra2ElvJywpeLQvJENHUYXtTG
SDPVOaSkZDfQj1ezM6kTX8ZQY+WQ6PhjLDz8tN8cyQURIZigh3tWTyOrKeffqiFwgIh6PgnjOHfZ
sozmMVcYjV37FMHTsuzA997ooWaV4upgKBaXzn2x8GsbjbFTR7EL/c4sWIJHVYW419LTEQ4ewVn8
QfklcFWvPmjVaA3hWNgjU9OkBNJh+XPJc/CaVwz4Hp0AS4upQB0D5eWGYFfkThuXCJkqLbTkoZtq
/tWG8IMJq3Yn6lo4AruQCR8D/IQLpXZza3pS+I9cbvPuXRf9PCeTDFYgFEWjbUwSyfeMZK6AIEl0
r1IL1u5aF0Dri/xuYHoTYgfwWX9HOvhr7wQ2v1a9perbFlQrn5b1XmBBTQsav6lo8rld0nRj9VKU
LxipcFbZ77MPTPKIoOnkuh1FT87wtXLiWqtSNrQcMDZUeWd5I9H/K64Wa9oNcmAEBjF/16P31a4L
wpUq0rFTrtxGFN930K8Z4mPAxvjyiOmyj6F6Hz9UJAyXk8Xzh1oH9BrG4pBrHV79vzATGRKfTh5f
zvhD/+M3HkeoR636IyDxCJvhotZrXKejmM8oV8pBYDkK1KPzaV/7PPg22fnGjAXfLXlTkGPGhqmF
XAxBdV1a2bIOEOg0JjwiWgXAxrULeGV6riDX7rUgXvLTo6VqQPGeUYSfmPXpmTTtkLfL5BH7nekb
mA4igkL9iblOcRY0Vl/dLiGygT26OqYZbGplLb6+euQXhtR7B02qmsMU2bjiVclYwBMHnOsrrE1X
6+Tm2HoKMlzh2kFoN9yNG7IU5zIVXnqol1mxFjG+mBKEe+wjY6bxIwwCpzSqa/K5EjQoG6NVY837
2n2WNBq6fhC/A2J0B7wYXOZa1XsAMDUSGD3SGbuK4iRSx1tcS7xbe1Z90GceDMMlytdLHq0g04JU
g5NJut8zPCm064d4GG4NXJl+Iefrhm+niEkLPEZa2mpEAIRd2DiaDo4Pl9AR7fyyUkw11CUcsM0S
8JA9s5BtUFTCIH9AryBJpxEyNgaQGaa8GjF5DuZBnU59FMUa8YbrlChvrlcs0WLEjx+2XiaLLL+e
O6opTeNA9Bx0KdWCk3XICdP0sK1btwBQObrDCXMtYjPbqswSJIVnDHWJoisWbAgRYT6QcIba7fmZ
jTSyDuYPgsSuzkX2vLx1+lTRbUTPhnHxtcddHNe2kdE2tvRjblHKuXUs2jmG/wIocyfUL6Vusbty
Gb5+OWqR6I1+v62kjcctB9cKIDyBdudFJi7zuWMPm1qJvUxUgAu9oOabZsJoq/mb9eeffJmxgrd3
nAoxlkMK3XW1OSAokN2d/amDHOsWtsoPabdB1lXTBFbnv4TyEei0E9TaObp+2z1S4vyregvc+sJN
HjAZHcJwbTsbpJVJvXJUgZDzd9rdEiFOQSWqsjLDt2Nm52iGarLSNe4p4IVJ5/4QxsN+Itm1xhS8
GYw1D4lAmG0saH7d3tt3heurEt97Kf57MHyuAmdjhN8/lveGIBwxYyi1W19xOc72d1rLzizF21Gl
6iaa9XpIPSiCoqQr4joS/i0+BocYtBfKnw5tFyid2uvhujqkxEX4Ro9GSFOYOyu7278iwJeKKwuk
4+syA+NbqEFJ7VglynpmXXMhIIVUy/yWANLgAChkl1FK8XbJg7vrPPvZphtAw5tD1ksa0JkvhxFE
pPijvgBaHHez6j2PctZXLtp4D1PhnxM60l7CAOuOoQrlTxlwahvR82k+tFfyndP2c1yTI/gkP1HQ
W4EsI3+2gODS+TZOadLgb4Lrep3sLvNDT4jGO9cep7chRaqtGngaO7JaGOhc6vsxfCPU/iSW2eA0
qsPzjIBH0vTB1nZzX/qxTNWnIDuyTgjVjcNV7Fz8gR8Y6kfJkyThxHv9P/ckstZXECOXwOqWDrYh
lTIXUrN6eg0aD7mjJc3Xh+l51ESjMvMYl5vNhuEjl2Lwx2N2qJLAaS3aPs1HtC6QqpB7m/+CmUYF
Nc1ueemheIghEWpkeIy7PBBQ3Xkw0Lo/e0iE7W6gdptrqa8FzQlxNkBTQFvg4SMKcWty8kgvSi2A
DxALt5IBpitcOuJg7s7VnzPCTxuKpvn3vqT9vu5yVzH0wbaop1Vjk/zJfBmb//yuxuTg+Qj0Vp9y
ajVQ8Zm8okLnaFTA43rygWz5//T3GIwGD7lqrrd+T6rXne0/0TNgf+ldDKNpjHG7DwSIMNNKpeoZ
4LcMlG1VJ6fZEz05g2MRHxVMD5ZycnNP84pULjwTw/upLuo657U2YbnNfwrDz2RAqSwRRzmeD8rQ
wed27A8FK1HvC3iQM315yUWB9y/KUgqupm5kEMtUEdVvH9E8Fqv415r02DmiXG8qzS2xUHMUJwLX
25h/vMRTueyfaDx07LudqfCtyZTV7TsTrTHub2qAGe5c82Fx/aTUIiYM7bFMfYBX+pl0ZFBNghg9
6ObseiwW0pk+3ihQaeei0ez8E3YJWBv7OM6+x+i8F1ae/DOGbqLMyBf1o1e84CrYnqTYgt1ViFr7
nASFdos53sM5GsVRRLa5HySJbEmQBlv08eeC6zhW6JSE/+Gu8YpUxPDF/eW0c9dH+/3m39oPJUTf
PVpguD7C+FceTxQS8zWsJNLQppWSeAQq2yqKlp7srk285K1URRwn4qtQunZheM+l9hHFM5XnYCjK
RYa/8FsT4aWQ08D8yIlTF+yDa017c+CG5JCq47tbqS+2XhLnNFXUa68LnWGmeBaCBhbJWZ8uEhvd
vb+RtgCPwIwso2q/YhsC4+f2bvYmSetgSfzAx0En40HSzhA2Wrjsit1JfEJfBHTEqmHPSGWybRXf
4YfMg5zre2x6i9RZyF1Tbnfh1WrRSJWaWkDH/p3u+fD0UWn8dmpKw+I4RB4pS8LEOJT/lNovkKjU
ljGhuuOeTo6walh+gxdQG0i2IXHKWLAcxlO7sYu80TCCEA5KzsQUGuPk5eOBt3igVzww7V0XSIP3
omAXI+QNFeqAJwqrF2xvkSNF3MZDiMMpiZTHxmEC2dDYTv0IHI0MStSO928OUo7nDuiqIt22S9PS
T7wUCsO/myhsmtRpH3TIiC5fyc3Zf2mWGT+pLjtNKYrzNO9oSZ1uwDoazfU9P3XVb1KJN7Ghl0R3
aO8dHELUXzPqkhcfunJvAoRG74u960zu3DuEc540wxC7vCmZ0XBeUH3T+Cy6MXcX9zVioJuwxHkz
GZJ1H7rYyffwKsFB3TTj/mqx06MIBr128LmtBhyS0y/EFsWVgGpnkugYq+3QN+1YT5g32ynj4Rux
fysvimDWP+vYIuZdmXXc4dq0+r1hIo+b3nHo3cAX/QoKecX1Y0n+WuFXp0FvWCeaQpfOkCw4MvEn
1ThX00rx0a8INP1WT+WN3sDiDzSfLZ/avMLGps1eOgU6r64eM0qjrH5FQaeOr23v7irw72AfEgjD
Uve0Z+I72CaoDbFFM5vs4Uvip7xKCcEjnStXOfOp9Uxw2SdSXZvMDGcuxia/2YRVXPlao80HeXWR
NLWaL8sGVcKlDbfE0DzdlkOq7nTEQC4RO9AcZDbQDuOZ9PdzDllh8gF2xzOn8mOmRvvtm4b11yeK
qyzkLPCtnM3Q2Qx7vCP6WKImQi8qtd4M/cwBG5ageCZMcvlR7uXJJRWABkUbkiXEg0w6725IpMNG
sLAiuQ7RSbMkDk5bNBWSlr/BtdUIB0Ce9dhA/7f8ICA+cwiTkKvK3FSuJWK+p5fsmgGH8K/Oa8Fr
2luo29Xkq5eHxs95y+DVzJCoxi+xcI96D1g7xSonxqeT2909YisDqvI3dB/gfiCJ7CIu322u+Z/8
Q3EvBmK6hlhM4i0UoFYadTyI6XLx67ZhzuAoQiO2SLYUP2DVHS0ZBK58aCdAlTEqHa0aWVtOYgHk
gYBymZvEoRr+5EW3uxM8c/c0n6kdGE7kvQE1BulewrXdn6pZIpyqdDm5ok+6/zY3XwVcdzJ20pSY
wBi5J+Xi06U4WH1CNEngxkFLmytCRl4hOpyz4DzUULJ1SHsZ4D7Gv7q0Zw4gh+s5z99+VJZv24S5
3TBXeDD2HWvbzMThmRhc+eoh/RnPGBU8JxSeWpjFe8UnoIdIeTZs23fPo6N2NnKeHGmsxmtP5GOq
wzMNv2xymZzXWMZyWjTxE3s/d2eh3ZkkIEkFMCa0pjD8iJy5MMmlVyH2DzbgYSZLj676Nlmh4ZfN
OXHsTRKLxPD2hoCVITvpj1FxtnfXrQJwmmyGz2n3fL1x0O/X1p3dpxBqcD8/Qw2yBqHijVKqK5ai
cO5gY8PuODmPx5GOgHtw9Ock1Fhzeb7IaDbOJFrNOQJm8mv5LEAQXnWmZt0naVu0j7Kbv2Lju8Sm
rH5x3lHB06fPN+9trC7BLCvLDmpY7TZB3WHTg5fLJT6MMP8IDxuwYEceyupfB08qtnWYboPiQMDU
YN7BtMqGszCDH14bhRgJWf9aYf0+dsOcmW7FbvHnmC+gfZWkVRu1HIs2WfUlQ79TG9fPDdPQk12m
FuaFCLJSUQDqzDkg6EE7G5CJXim6H55Z/VdAId0/ZFfKVRJBEc33gpZFKJfrKtYHx31A4vl965Fx
chrGXcrfBIuJNU7Mi5QcPser7td+x+ohmRVBG53azPScFsk9j8kUnLgN9PspXap93TWDMRLcjsin
eWUUWhOvYUSIUt2IjksLlyzn7xOFCNAYT/bx2BFAsviMD9C24zXf5dilGXnewL3sbW2e0cdyAzgq
//S9u/UiZMDfRn8sv50KLgzUTAm5RrtGnBGtI88ZjidCUW8McFscxd0qzs9MmKKFyxqLAp6hpBMd
EwLWgr23FqBm0H+sF+QpcZyhJXTwEP7D1d3SX1w+yLZoS2t0e66c2Cp3hEeOxKWJWxbhyP2o7Pn6
/S16QjuGvPfBAHAQiTbVgJ9fv4wiaSaPCEOtC915TvkPL4yKJb6pYdFgXvQvkAzJFGqYA20bb3JJ
8xJtOzq7pv1k5iTdrI9J/sKPdqo7MzsjGqSKyNI9/rRSbCIZhXD9tfAwnW4qGW4/bwYKtktD5L20
FxuN/YmATLRWyWIxhOB1/X1HeYocqxnXgoIZ31bw9P4YjUCxWG0ubreuTnjB8pWdBbI8CvU+Q9Uo
cTszuIK0hc9r+RydYPqo/qugTZd7uSVAyJIKU/e3lvxgmpbRDzaBzyU7SsQNdOqBynJ0O83JVT1s
Yyx+VvQmgh+PXfKO9Nthk6u+JgjbPqCYbVDcvVtABZo7j38wyr7gBXN+TT6Voutf6unpxVBzXB/V
o55G2uDGMnFSkHTWzs699+5nJ3GutDAISbK/Nnh73i4odwBGLHlkxBDdMEhUUzREmDOPMQ/vaJVS
oLIUMM7As65RV6aJTApVFEglRqgSdYp0QgHspZ++iw0IvvDH85t+aSKbTfZ/Qj/jm2IBQohJYzrT
w5jFpjoFhSlYKoIAtyP2mGz8IKFyKNadM2C3w+YzQboqfaV6U47HCUOzKidYKFQJEYbQUIqwzJZ5
O1CMkjcmCqh0mf8wbanLyxeIUFqtsCtPjEEd6KvJfmI+22zbAHHYbWdJitsFV1KLZh1sbz+sjSOQ
QsHYJow5Ie0rxYlpmG2fQvMsgHwt+TW1dJI+A5hjc8/H2+lMeMfWgUzVERLYteIBrsy8y2D7Usfa
aC1LKkfXU/E05miP+7ngZ253m8AhEg5GBRr9Ja4CkXuWYxPosaLjySI0FSmqk0rEtht5XKYJ+cjk
JkH/Ap09Ky89SFt24evMT104oIN3SXFvejCnqmuj8/lFEieSUbht3koDC16MAgrykrCzu+0ZkjhV
sJ5stzEKQHt1v54xelZkg3pWc8g2Z/hUtRvjLCnACzrzBfyxP9REteJnmK2T5ZKOHttRbIZI+VGc
i+tslyxWRTbcYzwV5zzT45RIilNtM6XVqXsApPEhLLNAc5wAkfVyhCuwdAle79Ae74oEsBA+ibW+
QzzLTRGvagetwd5kRaOgefMkTTI5wDnE50sYTFrkTeqZSukZVblzbcbQm1C0pTqdzeN8YYS44n8x
HG1A3dZy5C6gB+ACaS50N4awtf4IBumwxcjemKPffnGU6d7zzOSEKVP9Lg0dNlOSoOYP/WIvHC8c
uP8VMv3hpIxwl4k5m8VocKmaeIpbEOJrq0KYeAq9oM2pKAdb6MZUBKWaJfoQmGMxzG16Wkt7wggi
LpDlSmUngiQ+51/Bb6+EB14vvtfL84MgLh0yTMC3EE0BaIWAkW9K2qNuyeAdBuzcTlwngCl4ib/7
qpH42pnT5ePLkhx4v3ZX5MxR5lqjwDDn9Ra+XrzaX5eLj6E6OpVubBRAAk/OiBGQsqmKTcEH6dd1
nlv7MHoIXqUOQZim/3bYJcf2oy9JG+ETrQyWQ6t8bb3ygbTrGUOWhoK68+/9aoTqUd++xzT5wec2
p7OD4cbnfkYypJc+hdCLJ7qF7BVsajiaudKGdovK26Ls9neIYfj9FwaunWLDk/pqfIGNVMxeKZtR
9mv+L9gHh7ec7hGf82y8qfkqqeBg2om9jmRMvvnZfGvnr6D3WIcG1nyBaXb9ZIexV6k33YHH7Aeh
DiqWFJjqcGz6Ncdg+wVc7isOD8uiQE//OLXm/YFbg+ctTltBmU3VI3Vti1SpZ745msiyKcIj3o+R
p2Idg87PxGg9ECkRnIoXBnwle8hsxEFOfG6wwUQSyCY+0lkg3zWXuQNBEpMUQ0HxwUdyVtixWO2m
ija7T1CEmGhCOwmM73Zxe7Mh0XogZmI4B1zYsMT3ShX1DDuQrJkFIaHiqjY5ERDoz4sLMfAJwtjJ
qnN+omukF7s2XNdLmx9HWqQdTMI8B/LLWwEJL7P3pNXbJ5lCx5SuJFOIJL69yYSppsGxJpnUs4rf
vR+5GK03kUcvdS/lW3L5/oEvvnP9CuLKCQtqJpYnbzEvEEPcXZNELAvHYTnx3/pxSxg4pEL4QCEN
F3wvx5V2Gc/PpCjeMn5jTQGoRPFZEy5V5aT6tjwdHR7MLwTjZJK/Iu4eZqb7KM0nMjcVC3sJCkMu
1c2hZyI5RYEMjKL6wHJkxN8PQU7L/IdCiVA1b8WbYwo7f1QbfXbuD85c1xC5OBGSaCvtZV2tTO5i
Rn1CAei+gwmD/sKxWdkWnF0Uito13ZK9El65wcrbqdAiN7CDpkVAIrXG0HByfRd6PH/WQ81F973I
6OoIwVHYqpa9sYbhraTgCFBVWNxqJB12c7CZ1R5vzLXUxYmnrZMLQEHw8aRC7fNvX8CZP5bKZVlk
w0O7YfEAs0KtXoL5K9J1scVElRDHMArJeHK9EsIJcw7EWi2lfkqgVIx0AvUvBHj+A8sXUOyV9LSz
5GGok8YF8iGVVKM0sCOJaxnGj6F65Ma7VncacfmtpL93+4GjXNAT2EtpOgwEv3c6UFoRGO+822A2
CGprM/LQN5/EAlmv463eZTrsQgcPwmI/RNS/YSOPIrsaU/lpjQnM3CiWSj9IhpnGDTVUpmxgWj6G
QwTAM1sjTxKSQoYaXMD8wgpH8X1BAiJfGtS4MkfoTFy3npKjiWSufakxuNFRYrzHG8WjaFfUTcha
gCs674yCT2aTi0Q7yy3EC9y2ihntUZvIm5bBfVNDLhmT48Fzv4B0VNsSS4GxjUbUMkdbJtsNZWBd
NdzHYzMNKfh44rr1c2wKjVSphzMHE9pgvzCYFKMbLLIlVmpBk8U3NmNNX84G2koloWkNJLPkkBm3
J5nqPT16UD+IEoY5cf3U8zFX2wOgDEU8sOTwA1xfmikpp9mwQZLuhPtRXEvDV77AchuvI+4EV8Lp
lYLcsuo79Y3NTEDBXhCHeNI16v9ukCHlBnx9YyZOQKsuavETX/neprn3YWcAr4S07rNRTTbkzsyC
X5d3m5vlNuhtsIf2oFRBAzyDBSXXg871XE2KelFWyBwAOZesbv2Nai4KsZ0zyjBhCYMBISLMra+N
yK5o95OIECe3lisBSogQC8zYamQMMh12dFk4nN2tb+1F3QYCnK2EZAjk7/L1+atT5AhN+U5KOYPg
w/LzDgR0CX50aNFeHUHmEPOUdLXmpGepbUnGIG7eevJPZuT0AWbROrYWcbQTbrpZFSIQqsaP6Gj+
0uJzVk2YJMqy/QUYEWw71KlZcqTe+huAznFFBdM4isAuTpHpbydgk8o1CcmzRoyFqDnoQkjNYmsG
v/aQ6KlKr5pvPaoPr8flXKrFvxW7Htsw8MChs5bN5jhtzyHunmKNolBCUwQ983E0iVodLXCw4GcW
c3K3V+4AqeuGZ/VRJUfUkgLirNCabo1UqnfB/RfAVzEHBufzatHyDJOjPV2ed7v1H6qfMiL7GmnK
wq7I3ieYL4ooH7vufQlx0ZS1SU0xzMIWu/tsVaUTOxBuGk2MvPuMUHZkUM4mxTSSsbtcrmcRbkJn
X0MZ09VwLFhyoyGVYyYiitmZuVIPYcYqLYlJrBrVxgqzNLtmpQWnAHk1I0yCx3lgo4XPdPn6mnzU
sQTb4SLO6OhqmRYc36ue/5FISzLctgq86IqKnv/CT1cJmb5kqBCWH9bGq+d6j/K5W5bySTIq/rbg
8/Neoco7fEmICT5TILvmqLw36lGB1TUcg/3YByXam30nwNN5Yn8MNY+B4a3kahZIXgSnwL0RQR4+
GHy1811QiaSqwxomEDenaxqpK1xwvXo7CeiRdioIZLqMjrYp3Gv3FdRGpiIOC2QFDZJmKP5sWCXR
VxGpi1+0hMBuseXdhI9C+7A17/ZPXqZJiNFdmvISa8/9zW3EnJAD4vCLUvmVZhcZB06BFy1IX8yz
dP6b2KnM+2XgrScbSbqbCgmwi2Pk8tz7vw7ilgSQZff5K+QGC2Vm7ATtS+de82A+35+OkMWUBYS1
em6HCLNr3Fsd+Ttu/P9xxVx8d3Seid77UHjnlDfq/Bb28CkLAZkDJVZT9yZILmDx5HPQiwPFpE5S
vLH+FHdkRUbHxe9XGWSdfK4IOiHeH/cq3b2kj7I4r4JHxBr5j6VV5L6PUHKt0q3mH+vZCXBhiwUs
BF2N0g5KVqI82HqQoaFrY8De76485+Z+BPC63rKLBAWR586qqXQG4RR9dM0FrD2aBzT614JcuIkT
q1MASrFAe93bdzrgRa+/hEnD2lvtOx7WzRthika52TmR11PzAXiUVFyFkFUUWF/mXOJdz9RIG3Az
c+qMwk1DjO2C/5UJA9NCXBbn1FKhpBZa1yZjoijuQ9jHlR6J07JjX5xgKu7vv5GzlzhfLU685Vd4
dI/bG2jccf+vW5NtB9I9kFeu3ZEkdjqFtuyb0MF0+34k/Hfx2njAGF+lbyJcbRrl3K3qSIJc9dFE
E7xaGtAx9etDriB7Y5UrwLQTTIY3Uh9ZxBsI1zfJy7yLFRfWupUGyljdDAMZ9N2UGfz1QTBsayZd
NUGFchQ1zhMDY0JCuH/lSuu0x5j6jOXEyEmf9+WXDbYGpTObJ7pRjXw7r56IVJU3KNae0uVjFn4s
pYx0JNoabVtlDrS1MnsSwTV2nRGF+OlkcQdOCV8XZHPYAXbf3eQ8M1mIcFfSRYjapFl+Vnf44xrf
fbP14zebXkRJUuGC6DcBCCHQuAoDrdicm6sGuBtY6UXw5FlD8JR3UuAAS4EvAgvi6iec4UcZNNhF
61A+OAZ9CSwapIWcRICOXPng/AHd4tmkDCSC/N1lcxi2IF8bdQo7SQRg55AidpmLzSxVUd9zHa5q
3xftoGjmKsX2ksehif1LyuJIxN1MgRs6ypDJ94Bt8o2ejbtGulLVoI8HYTlNfMXVpvyFVigo1lK5
FJcedsP3ireNKNmYCW6MRuEqpO5YdUIMiqMQi2oY7bHIEWbFAjSuRyuAdnkkwr8Zh5peIA/dRQTz
fA0zHkyx7yd/aElyi5yraYc9NVGhAgSEduwW73HufqIJ5M0RuKPhkV8DHQUYN/0RglfdoUAaH5BV
Vy+8HuWY6Ghy1ZRxWIDJzEN+e4Z4pSDicQHkMyi7n+KQ82Yq9zRg1Z8l0FMq8tq61Klbk883gtW7
10Mrx0mu0nNGjCyN22s4X6pLofPjyKa650CGQiQTx1DNi4FD5dDoOhL6Jo8OUaaICZR1T4XSMwQA
NwLmeD+vSOzbLfqWkmQCy78PmToOQs0+NywPn2LDphJNPW/W9JnwEP1/R1aQZZMjsgk1BKscguLv
Gi1aC9uygXWl3t21P0SWm30VWlNdHB7QowphmFxN0rnn1ZIMMt7t+uhVoJS7ygokIA8qihvwAWa1
ZjsKG0AuzADYW7+2UDZyotm5kg6KZMLewb7Yw1kzoKDgDb6A6BJI53PPIW69Pqjouwr97dzdMbTt
X+oukIbp4r+sbkHuKYoprPgarm2W2lLs+rep3h1U+FVc4rub0VxUznrnELLaQHM96UqziVqi6kMn
AvsMjQeAM6tCjTbWkOmyQaxp6EfglNfdx56iesbe7GChllCUe/qo6nyHCOfqC2V5WW4oZZxx+qwQ
lW7ghBkx9WdZdmqNokOvTVPNWvSSf11DKhVth085AufS548TYBeV0n0vMuzrR+Hi3LtujoWGy0ks
HVfZIuqKRc+fKy6u1CzSKBp8HiT7OTm7nV9f43ApTnJO4oMQU4YrUzUp2FZGkN8Hhf1UHQtZ1kzD
gx0zrLqGJUUVdUwcVl3dMks1Dp/EdeaRMzzw54WHQxVtah8aGprJn/HRNXPzyVYyLDPRg5xsvfI/
7RtpfFReFCb/8RsOuY0QPIj5nUw18TNYcIXJfgFhqSrnalQobN5t7Q8N9c9IV6GWsPPpvAA6MfnQ
OrigzP0hV5EscIpRV3vGIFIcl5xQuRXKIhPwc6lYbTH8/uIjLCofDkLw+O9Gd7/4oZFrEvCUj0wc
gvdFhJb5h4CY9VyMLpNJ2gHvjtOKXzBCO1duBo2IBTYfzGnyaHTU1Qg7H75dK+59W+51UgnUbXXQ
fq/FJj4TFEQA3uReuB4pc6LUN/CqC74fWmbBVNqDgWmmD5jJ31LcyD1eoP+4e6KPRQwX2auEFeLX
FZaetL5ANh50fLp2lXPqnzy1jk8lOxm0NvIzNLsRp9qkDAk5oR5fyBAJAxvBZWaDSoA3lz3dRowk
11ERtbk7nIUzHeo6i8EjXNg9LW0baM9uGuYBdED9ed2bYy/jZ7SrxXGHfM4ZDQ1PlVVCnI00vy06
a9DMo5Y+0du65+ZvczS7ajQHgcPrpW2mB0uZXa5hd99F7EmvCDBjSjx6ygskDQLV9BuAOZ8T/UnT
DXPHHJhBNyARTN92gL8TDpOxXJUuflOpqkwR4g3+ZQSWIR6I0jylhDmkgUuJghlTvx6nAUKS2nUc
WP7Vk3P2iBstDglRWsCOi9fFqQLsYZ7NjzvN+QsoSHe2RrEft54EyJF4oPsq3k5gRpOeiPe0biiH
PxMqr/E06dYEaHtFY+WLlLtnWvOSbLGE9XjbQvBQlpcrfRBXDB1LZUKntAYhCXuo0jVXXI5mX4kS
7dHk1MmU4K93TobV5MK8DcwbjtO2F0bvtwYRZDfh8X3yQ7nP4qfwmtC5n8S/EVT8nokGxJZwSgIV
His5LMUmCBBslODijiVqjIKSC7cGYaoeqX8+FZXcnpObNt4IIWyAPQdCg9qRucfdxvGR/IZaMO84
UfMm49jWJtH/y/TOp/6RAvxKzYQfSUpQ00dJH0zfhAjMoIoVHTiva6ylEr3JnbuJvzP2ssblUk96
qjTHBL5KcgG4P40RO1ccqKqkne1CbAOWvpOW+VqTdOs2bjv8HT3+7xRhJlgLKf6mU8VOdefyWS6K
sGYiiKhJaSun1vDRnpSfkGgpsoT4dWqtr7TF+XmfFbpmlxovKL4+zLu8APf7nnbcu1zU5qRSxAYB
fUJWbE8643Kg9XqaQlFN1+y4NgEiQ0Ja5ucnEhdiTJbPlHoGlWRVn5MWebhcyslht4FFehoohUOL
5nx9RzCdYfUXnhyvflCRhwVzb7U0LpaYmqrEtKMKVfVZ8c7XtQ599xh7bvFYmyWg96xu3L8iQxGn
Nrn6TyCvXOwRES46cMmJd1rEF6J+NO8T/svPetuH1t5rKruWLCxkU1ql06eAA3keGqyG6BiHlkdG
28CsuWnDS5PiRlz7MSk9mZUXK6CpyBxF/kbdB77D/v8GKd9NnLPlfXxdvvAns/kkjzL8zvKYi1XG
c1Ck+TDcCoIWGrFFbG8aJbAEnTiC1ZXXFwoCNDUmq/bsPBlLoyJNLRLFBbQNg7Ya4+nA1sDuf9ti
BwHGdtTefHfm4e/90BWDJoecBYBSXDrjPo+f3DDYIIr/EfViaAV6OPkfKjcYATM+doYW0Y1T1L0p
xklvB904W6GFS5kJcDXHl5fBiJ2W14d2us8xbq9Ds0VFobvmcv1WQs9963fh1mcSNEdBiNQr56zh
S7EbdkezSoaefQB1pngBT5h6rTNr6AQydUQ8jN6MLfz/QRh64j0t1X+eWs7R3ApKnOSRQmUvC6tF
yaqMzRWyYpWXgmOtin/TCwzAy2PYc7B2Q9GgZxXwh+81iGo62ahweY4Ws32dDik5FmIPLvvtHqfX
p6Fhz/npYi301NBgKho21NHsZnw8b9peNlVTTcYm+XVXODhaozoW6zxmgotHQhDP0b/unGX1r1ph
lk54feu9oyXpskmzN1bp7zvUAwRiz6yDkF7wdKyfZuPSKSeqOo/EqBxKTH9Qg6200nJ/TKI2RTGN
51UF2y9H8DhrlxLseYXij+M+w7INRzBuT5I7LDmI8OcGEVyXa5/x7yDK44hSIjxeqhuy8trm5HXR
sAoZTogxqoMVT2QLp1a6drVX9JOPd1RMBYIgrpHxAX5rpkk/XNMvosNRSnUf7cIw4813Gd5bPTWC
qMIYWZ4faNgeMaEI980s0j4Nm3fqbOqAcnjrTCfObWQloKwsj2a3D5YddoolOqk1+buWw1/NH68O
7nkoXs+m0sIYeWWIl5V59X+P5hmZ3lmva+SYYVadMIkODefCCERfrYKywpZk+ZabmSQ2591XO8aW
yYgtU+N3OOjzVYDEDMjuwkW1EAB/TEEWjYmsDUnzDSj+J/XZtpA78r/ZbcwZMWEe+1zbaROEx33z
xltaXkhD30HvS9OFWNeeeX60ImT1/D5qpMdJykM4/j2jRjnF/yA/kKo7g6Cx55F2InZ8xAaZA4ey
nFVu2Y4hpQ/AuiXJIa/EoGtFXNQc0XBu2DSdKSZBW/o7SXveO88fkff2jyWRrlumboPUM+FZFaPq
TPTra26MYg2Yxsjwi7CeY6afEf9AVWsn/UhmgH42qcWqNqNwuaOopT/Iy7gTAXyAZpoVo+btMM4/
XQm61mAfKwEAwF7ibnyzslOT/QbacYrmOAKMCclDTaJQyYO+EqSg0iDqvI9PylFNydhfzSM2KfwU
4Vx9W6tY/gcGgV9si5qG+WJE22+VHDOlzm2PoScRpoWo1aSbUFDwaRAobZOYiQc8CnPuJkighzrl
JhGHXyRrkjV/6G91Ebc00l43UmJzBLSVme/OCFTTPZWI5+2YA03Ai28ka9mHyeM+L1uiWY84Lfpc
hQA8r2lX+dQwO/xIwttNnRI8EDVFH5H70lWRUn3DbSVLQBGZw4sMMWuXMqqD2zzR/x2KR7/LjUqv
cGzpwDl8HQPUucfyvdO4aATRMMFGsLFZY4eNThpx+aOsJiViYi6weeUWk2eYQpZU/qGV0DScFBHc
0Cb8cbqPLef5Ur+0UOJmoFdvDbuZiPihiJDpmuxWYXhCCw0Gkhrm+rmhK9fMys071KG00nFVmKFJ
fxhiPYCTM+ViLn2TgC8YVhD3HFnzrKgLwYhyvJEXoVcPiwu8PLTkdbxVg9pnYH7un+V2OplEizYU
8nWYlCgKfXe1JyIZyrrJVOhL+j2KguSK4Ea1ckSmjpS4dIHoIUb/KdMVeoFYSUX+5dsvPTK1GjUb
f8+FbRAFFRXPDUVmW9IOgTOFIAz8kjt7NQI9cjy10i9vfBfjpnHsxPnBss7154qXEFrbEYQ1WAS3
+3q72RspsZudNEFNbBBWKM0LNyEGnUorPqv4ZmuDmpXfwUKvjwIatUAR8NKtuVtVBUFZLgqoal1A
6bflb+BDPkQqaCHkxkvgnbnKxRzviB1/IUqMdTS4qRl4N/PAfNBhwQFFduPSrqxnmiV5KVLx9t0x
m+ajUS3hFibV17TYMQenkhY36sp1t5Ddwsh5GoAZH52huUrJ1RlTJfY3OwdRPcjzALuz//CvASO3
x+zA5D/J661/lYVD4U6kvc5Q6kx7FSWQDp0qXOlB3RthfxdmlHPaP50QcRLuDoJNqMt8l3zWK00m
FFMA1Zsbyf1/ywdz2bain2H3s1s/kI1tFRR7N60jd9cl4zsPENh1Ler7c5k1Fedv0mFtDt4bf387
WknHaQBp78qY1CNmnn8ETwJK2LEvfEEtWZ/ejLewR0kZq6pCfDmCl5oBhSiNH8pYtgogMB7g68Bx
1uiG7AaMrcu2FzgoAW7le/gTfnZgUv3ybOUu9/dbknk+RS5J/gd169i1qrOnbq9d0foYUJh403//
2V3JVM/bx3VlMGr8MLmU8npxsm8kj6TJUyclWla8O75041rQ4/Cu6ZBebL3EKUkTw18oAKLGk/Ky
XtThIgmwkwCXD9arxvCA4uqVccrijVc2YHrg+CKvZVjohofUhKs+IEBAxrBG81av3JTpvkLyMWDB
4TpGVL3x51TzzEpnI+6FsAEyCMwqluO7nuw1u3BQg/mCTFwLDyoq281BghgO3Qz/cczkjDl2UxMN
7TuxXQhjp1eR2ONDAsc5HzHRNVdWAQgyORBia5cUava5W9Teo+ck+Coej6wM9hn9HdZuLvl5/vfo
9G+eMXBC5oXcYtt0IoWsGs4tTIcLoZUPOJgrFNkCogl6uPmtoiWrLCqzto9+0H+pbK+9hQXhoA9C
YWYiwTHwaxyD/A8pbYPAt9xLhHR4+YZdHVwlj+zhbH7TpGvXaM9bKXlt4krLhEm1HVihQgxGRoeJ
a5K/02uCM9pudARvPS6UC6vpp27sZ/qlX1nW7q+/ti8u5LDz73tRV7I4DkkYF8ozuAAc+4+Cz6YC
Xr2xWX8tTPcRSKlbpD5RzdtWEXMTw+m+qhGPzIa5DnKSdLs3fdGAGDHU5I4DQ2svpo3j/DEocrTG
ARLaML1FMqbk47EOEUMjasDUZlr7K1xl6SXStEnj6RoWlJaZ3JxqPZj0E9qPXaMl+MJMsb1G22F0
CRtzF/xrIhg5CBG+gVu71xt4EVcqKuUwiCay9zgwCDP3LtzBC41TkvJPeqk3u11g182eUKRCISNa
gOvwLCJWDeZYcT+PnP109/hEvaRp99NA/fmmKL34vRykOGGeY5mWvG7TXIaU4XLCZgoRtQoSm5gN
T7lI9BeEVOWK8CcUKZ/7OSjIE8lOIMeT+s1qrbeWdb8LukzUSYbBjcGyREFn3UM9vpvFMYjGHS6X
suh1Ly9VkAIyWHas5P1y3hXjfq1+/a84b2DtHwOJgbgdfR7YaeoYprHvr1ONLoL7MPsCmsHWk2im
TAhaK3FgPucIwwk+9PtGm2GPDHk+28hfVSXws+HjUuZez4clz3xUt/Svn0Mq5FW3Uii/6ZEDQukQ
zp8veVAw19/x6Tn6IqQ5aL5Om2nGyp/c8TD/2g0zA2dZdT3vZW6vUpG1ya9qy8AoFWjCDPAI02lF
Tb1bJQ98RoLr/ruA0iDiZsKyFIMaUUkf4G9BnvoMCvRzv6SWTigxwfirHiyO7mQyoSby/CLtKF1q
vAJn45OnoKunp1RsbgDlRQDb62hyAoptooSmvdv8nMcXqUR3DR6iTiMOmDetp5BerqcSA2hwGvU2
CZYMfZIDJTIbVveEtqOzPPA0J91/xobhZUG5yH1BoHoQLNQA/K4fLesvPCOB6WiKe8yDcKb8kP/p
Urdl6uTKVA9GWy0EQfk/5D/fvF07YY0JecSkV9oXnv0U42sGDVD8LokzjkUaYaZ4xxnjaDQujX0M
4avu+Gb0rMamO9nNf+QUgzRRCOFhL9d4QF18iPSyTy6uRvuf8iG0H9zhKz5bibnLbjIjmPsKekzM
Syz4oIfgePRbxM1JLpBFHvtwULmRrN2Vbordc4oPgJWvR9q5J5gpAU4tESrWBKj0nTTe96wTSwUE
SdMaFl0hMsV1HxdbjBzFlOGlhMBORihQRW4ddvPB8hzo5NT2tc13BUq2JRMfDAvdQ8w0eqBlCRTc
4cWkWfjiVC8RM3PYw+2jxjP/mYs6IhmIgH0kARv5OAFLxCt6Cb0IalIkOI4bTVvhLLjefPhNRLdq
+//iyvWUQ6EyiNjO5hoIFuz3Z++e0OMg62018tdhCO3beDliWhOM9lvqdveCIVICd62LecDtIQvx
fBJr6j0EaetvvrntoLkcaxR43fZIPJaLZpSI25MKfdqFqDHcm+LIHsFc4duHY2hy7SgLN5x6MfXu
h5fTru87gZMu+0pOZsagSP+q4VDoiroxAIb8xNNJXm8IE+lKswvGBj+sO4aErvu7LY+ZvDgTic05
Y4Y4nQAPOeueRL7VPi3uUMNnE61rh8DoWMtcTs0v8XmFbVnwhSjvShf/HLSB8Vvc8djnJQDPih8C
7TdP34Hqj9n/dFKY0wOx9TsriIkhTdDWVOUSQRaF+C4gb4dbgEK9gA6m0q0TgkxICk2JTQEbJqpW
RqrFIqh/Sx5Dc+4bDATpZV3sHQjEf50Yetzqm4GG4nZOouLnfYTYg65KxrZ16f2zPF0cema2Z2EE
95TBIdpMHybANOtTTPl+PO+j+UnJUEczFCErJh5K3XpQoaWH5zAY2cqpaZ5r6gARJk9hcnWiiVqP
3h0uLG1Xm1I8YyXw0zWf9j257poGMR4E03G2O3Ozpy0xTN/shLKRwdAqFSrUgCOHe/LYmpXhLVv6
s8J9Tq0rp4XSzy+of36b5nQxYm7RrfDrppGRQMFUZC75Ws6T4naX3e+gOMoqClYm3eI5agBn62XF
UguSBI6yptkZr1EUp1LN/4ZPDX6MG7HkglVz2xYcwVYclBJEN6SbnQgx7iN1JE7k3j/y3buoMgEB
AaR8g4S6tEdy17II2ynbWGOdscc9CBEhGi8WLj3CwpuVNEgTDpIN6dBxW5B+MVo0LdLwDRPRn6Nw
3Z6hl9fObpxSWLphkhrhn+vFLZYqOv8ZeU1hSLh8VMMUhkXaP1aiRwzLiYcNAHASy/rDSzUQvdkG
nKq0LAyXEOi7CPV2/pQW93fCdXD22DgLAubYLd/IlPN82qZFALd/b/rd9uF7okx7CrspaNF8oOln
m5kGZ0N6EyyJ54cO5u4nfmFrQYMVOhNOXwaqhBCce/GTKPJXF+ZG1ENsi5tirKTqH5nvmMEGEiR5
2DlxF2NIpvE7X3IjGhxTPGdW6m8sZo4JZpnuDQQ7hSlb+RcA5URwmabGETgJocURqHa8J5Rfyrh2
FX72I9BakE0PwPEdbpKRJnHnEm9a5xtsr7AXaTenx9n/YcWJof+JyYjv/f00dje3/2NAW7RJr/2C
6LI7/1eaBZb6fhs0mLX01HWOaHLIIxaUlK2xF8f3ABILDvx/L4SZLCxz8FtltBeyW4ubTwIgs48w
XRXQ/ntjm9VGsI4ZE7QZ7Of/ePKRdaWikZDB4O70EMh7R6ygnTo9jI/5eh8jBVUnteEjtZpqwCuC
bLHlOQnE/kOP4g7tuPGpfYsnMyY4zRRqSJNXGx+QnvR3jS9y0k80Rvp/aN4Giw8E2TeQ9NzDu4x2
C9OmsGu3JdQ3XhZH1vZLloCIVFKIlrJzZErxk5N/nHb5xE+/3Yd+c4WwAWdu7norvERCg0Wx+5vu
RsErACMvHkUdtqqWWV70rEzqDMqC7RWdQI8NF2UU0UyNmDCDmCrSAAKgz2cRKr+OaKypugZucSIn
y+aCjKvkE9ouus+eRGoh7rLgW36eJMJrI0IyoFnkEFEDchs9CpSVnaTIzO2FcoNdlO98zhoj/W7X
S1e0RRJ1vVq9di2LkOI1P+HEP74eYyTbJb1DXN2HVrBjYn7er29tk7vmH0QPMObnjmeBTiERwvVX
EfsWjZO7qEjiD0bLdtAnnBIVcy8R12kQCv6F4GHktvEgW07/cKqFdS0X+aYimBhN7z271TMhSGwW
Rcs3Xz649FKZKqUXWpsQL2iSm+SyIWko0mPpfGEoF4A37xItaruRvhOYujz7co9xCHWpxpICr2Et
f9uRRzl/vpsoQW778z4loV1WN/z/q/jec9TR9W4F1w1arKbA30R8S8h9TY/Ipg9//p2lvSckXwpV
llx/kT+Tun4aKfVuijDsbRfzS7N8fUt4WO5u/UI7Hhzm/USXCTlU4StsETaUcy3EJclZnJY7xAKI
976Zz1Xhrc+WTqhNFzUFErVrSdZRUbkGczZYKZZIZ3mmGjUPKySYhV4KtjMMC0uZsf/AtU6nHz9X
mMb1GDDjJC9judIJkvmQa6mXEfBjUjqELhZ7/AmfVzuKTtIl0tvSXN5NSI8vc1GVga7vFiVJCwP0
HI/F07DFIZDsTEnIYN06LowrRbTbbehjjG3drPyXcpOiRjEJ57ee7I/mpztZRRv+F0rz7Pa5GdTR
Qqs9VTgeeEEKkCX6KRw84Pn/V/yLrH3tdbwKl5+pktCtDyXDdFjvohGose1a1497d6CzcVzVv7Y/
/DRrDmO8WQRf1k1mwPpqM0kul8P9tUqAI99+f18XijKor/vEaIVI27pTqKb07jOAXhLnEpZOr1Zq
Y2qV15GuvqPudnbrXGzSJQx6ZXiiDr0SNBHEPyNlMFWmQnJyKZ7F5xy5dicVF0zzJfP1cK3N/Ody
9Rve4i6Eo33xcT5srKMAJgqgz0C/vg0wZWfN3aOhGoHg/PNHxAlX3Na8PZ/boLmasEhHCZC+Zkhl
mKbYe0hDgl5waZnbv6v6T06xRSGMWTGtFtfta4Nwi9JLBmicXAvHcKHiG9Y9Cn8UPIJwzduBrGM0
BsVSueEHy+ZFnG7JHYgyC2KkZ58+RZ+f3TiXSn75ZRiy/jDX4lZ+Rsr03pVGv5Ud1urYk+j9AYX4
ccF7Su54jy6F2Q9CUKW/kyCeaDRBqF6nO1hq+K16rbjIBWTvJo5N3JWa9/7/UnreNZsknX5x46NN
E+6Uh74i2U9deEMfEZ3FUDeiRLmTeRgYp3yk2GJm2+dMTq/AibfH9TE9TzeBjLc60Wnfvw4dDS9X
djULT4V/kFwV4PZgqMjOouWJkSAqimsUeGGRsmaclhPLKAVio7eGF2t9v6tn/BOOqXsZPW0Z8Qsw
dA3Mkz6nKsC0JLgTVi9ok2G4X2cTURBkixuqK7iBuwR6sL3A5qtlMgsyBQWp3qhGx7CUDudVo9rE
GGT4KFpEeK8w0FM3vUw+sSH79YV9+ncvw3pm2cWN49Z6cus4VzjpvBcrNgfJfH7d9Vou0cAw9V7x
r9Va7PKwUeKkqGkAIuRVCmoWwpC5omc9myNt6a5w1fyBMNWK9ALNLirtCdy/DNcqj0J3DIEPPGsP
9ovqIee2ZecfjuwsqJ55nIzJtAKffck2M1XepinrV/gqlQYSd06OfK1U3RO2Y0KV8TlIvh6uWsnh
RLjyT51xY4YPnOKORevWGZadddv5nJxxndbDg+czXtScpF1RB3p6EzZFUQ4lOr35vS9q8GlVhUg1
SyezOlIBK5Pb22FraYuSHdvSLJSP1m2eGaIpqHDSk336rdjbD4hH7SEavYiqFTvF52M39R3pkVME
kk9fL65MM/MjTQo3dl8mXHaJcE8ThOWYwCAbPcOpwsflKQKHDVFgPhEpEXsSVLx9CrAlmATfSbkl
9HIea4UOVjb/9ykWrDJzTErgMq+uGWH/kOXm3JYnUKUdLNdyJCR343kLGL3Oql6CYz+VjkzTUV9R
gqAb57RgeJ2Y4JKytT32+zEoU/N77kUMIhg1+Mh8TF08CxYfvHXynp8ueuTvHs6/7UjH/0U7Vmsw
3p8m0Zdti2zInNQbdNZWBsFVXRIRltgymbjDnCDtO+IciRDm6T4DstOhW3kdR7tH5Cj4KIJJuuKr
z2sSMTed6MBul4V2fUUuaRHn2KzHHh89EHIhnTgOcQEBxfTrZD0GGtQK5hD1mBkTgf5dC5KzMm61
VD+7CJz0T8yVKnLwpSejmftyeCffCwxUUyyXZlmU4XgDli9Zgpyxq7KjuMJptefj4ABLZunNXDzD
fcTSJmSLV4kqvg+uelG8FxSduuQcjXRt9ePV15ByvKOTED5tj14hkJZe4FEQyWh2vx8C4NwBdf9E
MsOAjXwUMBvFVSR5ofzQbKFJQxSnldwFKTeTtmLUEgY2D5B4OE1A7vz8dgTIahwmZGQiRM7DQJXf
YyrDdqZN0NdLgQatXDmJL0BCpALqj0r44Kb3LK7nMYTV8zsMf9tJH54krgYFvCSP6t2LgVbS7R3w
SDKDmL4GsW4l6arJgzuR7P+qenXcADiQJEQO21+wpPI1MypPJtGcUsPsKfm8tGgBZyGpWmecWt7b
/OJhOYSLs1OTX684HkFxA05UzpnBdAvmRyL0N8mrHmB0//VVqc8ERHNChLy63/ubZI83UaSaz2y9
TuU+tR+blGM44Gt2tjXILT92W2ADlheXAs/+4+xNqFaIhCidYW60LF6uY41Xat+7cQ/t+RcSYzYG
frk+EUpB8AWZaah20cgBiRmIWKBXLh8ZnGX1aH0WairrXkWo+rVAsUfmH2RyiQR39v3aCulxX93v
/maZBNALtbisHvyqetZZOzdoCkzy5Pwe8Jx4FzTT1mTHn/6ikwHvjVv64f0HV60cjm46kaub/wkS
QoPUZqtavvrpSQuWH8orDfJsQ+WqH9Wvx6Yg7BqbmfXDByHR+SX8gbTwXCNNMjiUNre82jlaqksZ
uMoGMMExXGzhkOL6nx05Q7uytU26gW8PBxZFMchJFFuOjqqnNybyIvRx7gRCscRo1t2+0KIe4/tu
8YVNnSHLMIIx+9VFaBNGfuBNxoMVpk9YQxsxEXyid/kdJh3N5+hL3EwILcVHvQhFGb7QItxF6sr5
I1NSlUEmGsxoiebnxRg6KCQGfy/C8D1Nftx1PH15qv7jPyXpxGbECMqJwyKGxJJo9rp84iczLLNZ
nK1zy7+qgZ9klfXgtu1mZmeNGDOLSZ02QDjrtsE9B5zvRte0weDgh6scnIrZYKDD46cx8Wik2tRf
+igaFMWyr45PJyYeXPSRPEcofrt4rXvXmzrPWOnFs0DkBzCWF/4S13t78HAHzY2w3jDxfjF6h9CE
nzt9kKlhj+y1jNl7Bpj84eKC1fh1t3739lBCsjshuT7xvpuOE4euuF9jcXboauJOo/P65Iq0gWT+
F2U9yfNO5posJc0JBMcl9iHY5T1ftj9e0SLG5xnpin0rDe2puatojeEjQBazBRO27LHQDUyufN9s
xrG0aXEmJvC+J8yOQd8UOg30uHBWKIxkdGBC0lLtCxoGSzJ7KOFDtOvHRMLPX1eMpT3/icg9Soge
H0Yu1rF8DSD0B+07SdGdZFqE1i+5zlj/b9eCFb5JXYdWCZggo4jVIrbwwkgIe07TQPUJyENN9H2L
EHzdWYwXEUf5enzq6EMm2NXvBIBGNksVsUK9TX++451+YZrGRJG1EiTxiZCX8mWGuHD/tcpKUN7h
rpqW3tsFHgRWKC38b6UtPMJ3GAq4P98LS+0TyZrp3Yv8jRaF18QRsVkmLru6tcoiKCIf/vj0xz/b
7xSKRmxU6Q5N+yT+K2TPglU4HZ7NdiSx6Wxn4EDRJmAOoO4qTnrVtiDUQpWfIecR26BMYoSQP6j/
AJGCJs8d1+ffjZZe0RQQsRPBberI1PHg7lYKOOX0RbL1yPeHPe9Z7mynsA2fDMzhDo0emX+3bq72
uDT+bP/x+EQ2TPO4yPIL4BM1SB67O5NBqSfBWLapJhZr+2Z0tNimocm0S47CUp/V7jBlMWpy+3P8
isH3RR4ZrW8UHWp6omFz2ML+vePwrNenNE0OMh14LrF5RLZOeBUSdQfsNHly8zBurCtmVDPrSH0o
3DEHyj4QxZOGCIFT6/hXOnLVRr5wdmuziZWY3kvt2agnatgoMQvh5LBN7m8k2yXDdtMIV/D/FB9g
DJWthbjVh3bzylK9IbZdQf9CRDkhPwv5q+Rq8fyKcV1v6x7s6fAkMdsV6OYD1EpZdNtkQr6/CfRU
gXfNnuN/gkOxyiw8bKsAYRSAaun0yB8Ywyjstct2JqdrqQxi9A+paZIyWEg4pjedVX4ONXc6bXJR
S8NpAZM8gu7lICu1ZVxguOTKpm3ga8iqrSNZLx/8jVzv7/sAuSuHHA25CHEu+cvpxoo6HgG5dd8C
zScAiuiNrBfdXlk5bCyJU+UeckGpqjZAfrYlZblw9VdNaAZKIO0RvrIIyPKXcC6U6kglGo7Qr+2N
xSDQ06V2NJFKAW8kjo6irJE/EF9dw88qcpc2WPtKjv5vbe1gLhlL01VMafV/jbWx4wLrUdD8vlOn
jIsxP4DvTWn8YndRvTggBBavB1suWevy7kIFjlgjC4g4baa3yPqu6PjFqfLjcrMxdCsgsHW3IBc9
nXWwaHsqJAUONkwetkVY8xpyyFK3YkPvi9sCgReJEbCk92r0BNS37Kr9Qz2nt66DKiqWYWrlKWUF
vPSOn2qpxREz1NJHg2UUr20+XVzxVHZeO5q4WrpB/anxUtCfNWVejpq7vPkxZo87NtH6y0vrYO+u
hLYg6lY9mCaIA3gixSih77zxntQMB+MH9bKIMFRBFR+ziI5lSQtRctJBU0wGFGTJK4TpALvGx/Mr
K0gMDuomsD+SSYnpskNzc58RqXbwvllFlq9N8MU5G0/Mg+d72TzYGZxbYkYY/7z/fAL7/ptPAmRB
pqwuodmwPP+o60eu2Hs4ylGuzDPlhzOjXfYFmd+TfHs3+VAzrdYX484IeSSj1piJJsr3Ax55hT6C
FmFoY90H18j3T0r4n+Jra1Mq7n1Wldwvi56YWrcE8hop4ijH7u2t/B1y5GBIfYDY+qijTdBHghPW
xvgdO9R4hRQSCfEmQgxEAb9VzFIzCLEAVjW1h4zrykbh29WkSzH21jlBSHxV5ZZqurcbp+25XLV8
UOw12tVLLrIXl7pJVQlxHTfAz6JtCB39iRBWfoTsNHej2opsAbx2p0oBm4JJ/42FAUJ1sW6I+goo
jx5Wiip5Z5MJfZ7EgKEoZK/yrm7EvMU9y0XIO1b3d0CqzGJzRkjcfzpYcUuVwcI6B8rz7VlH99GF
9D5F6eSB9Yc6g3+LcHIjpX1GBcwftjTl5s163jTAKg9AeBN615Y6UZAWcrXc2T8LbD4fmS9nNMYs
n06//eolho1rIZ2ogk4PDEkCluQ4AE1reKPcqdEJJexV2L0m2vagpF1E+oeZDh4Houh2P9G23LzR
RNB6Yi4+dVp0eYW0Dnmz0sEX8o41HlQdHSJ1bgyHX6p/Pgl/HpsGbLQ7UvdudVt+8NzibR+oiueU
Nw6JtqeWE2b885r2VHmjYcBiOTdpRxCVUvTas5VGJpzzl5fk7Ls7jyhOakGhHgJ9pqfU4ANrEEMU
6kgE6e2Bw7IhcATroK0kV9paq6N1tLoarvX9LEy+rsLpByOSZHYQcPzOk+sC0ha7KuMUdOZfBit8
oQeVJOaJmimrplrMmddpp+3Fh1pSFaB/cJ4AfNF90rwDbdEU4GRhMzVLl3Z4n0+z4e3HY3HRsZX0
cq3v3OcpXFeO6ITmp/cTWeuy/7zLdKkZPjZcqsLEgLuUH3lLmKjpQ9BjtUvK0N9n64gfJtrXwJi+
CGm01U+oFlffETEpEockPHprPwSEnDnw+WTR2qHrz03jCHsOMNZavNmCnw8o/LCR+jtES9o4jLS6
ThcYZtfs1q+B32AwihEfNQ3ibQqhufvEILn5Lo95FlmY22jt2ejplYQEPiNpK/drQbGbcBUq+Gu6
7Mk5BxX5Wajgjgq9DaWa9ZG2pAtw0rxwKnHFhctL81QGMbQRX7AvTANU+0lhaRd4NrgHAQgFh+6F
5YzW/RfctUmnfwCM8ViOXOvtHgT15iujCks5RHvCBEo18pRizqnCapxkkaOiYhUWmxwYqzd0smQe
axc2hZT3IgC1RHRQbZEaklOE8DTLHGXWGYp7V+SmJBdYJ5iZ+DbiJBMGsDag9/3e3xlYhl7Shrzt
9oAmb9KCGq44QYIeQ0jah/Hqr89vL7PO47eUODu9xUq6jQ08EXTx9EFeAEN+lE4+DCHAApnOgAqe
Ic4e7tkWOE/hrOvtRq6MlqQoPWylbw/Frd/2dkHFwGSI91u1BUG/YU2nuIIOf5EwCaT3yuXV8HXm
ReGfaea1b1/b7wZmL8cmqyGGY9MBkgtOF3l3NJ7mvSVLMeKQX5oU2ULEJNrHBSyK99sDCxzqsnSk
rD/d9kqV0JY8NX7e9L/GK4o5RBUuOU4mKHgnkT+Bybi6Ivk1S1JNtnwIK+gLlnSB/9zoiXrSKbyr
FH7YEhh4kElQLyujukZ6f/eSSpfnT2jie4K4O1UN+AOYKQ5vUe/+2kZvlyrMLCm+UPOypGz0Lbnz
/OjV8/TckWuM7e/oW3tVV1cW2U1tZe0VC2CsVxZCrKK8CA5XWwZE7IZDKXAnulTthCy8XdVkbZG1
jx3zt7pApbEgc7LzEgURMewYxAA0t7Bhrkq7mUcJ5pEvHMeokp8fD+QxUEsGbJNOmjLYdxBJWhEj
zEFT8ldRCkmGa6s7cq8xrTBR2ZF06UqmBYbkxD+p0CPxit0RkT8P6XiFD5ZjhR3NDFXlhoaavJMd
9YLbqR8rBBtXN148RhfmtuEVjXcqqKuqfw30jLVo9DAhnVcN45W72Rp3IgtiN0z4bh0YSF5OobU3
2xJOIKcRkejmetUcUpZV8/Qf3HAxkAUoAtmdMwXJr47GRc+qyZ0wBdraZQjPlAQLkQ8gCEO6xOpu
f5qj5Mcnb70rq5kiIZrZWfgb7bVLGdx9R9WIFAe8YsdEgWqkA9uK/r9kia/XTnsjYSHYYrYG55mw
3VOIH1oRvgWO5mo0aYyZ/B72Xi/o7k6+0uP0JPxuPT/hynBLRRBVqo/dPDttIFngvhTx7O42BKIs
NTUdU/wOIge+DN1xs/W+8sh16gY8Y+lXy8i3orNuvVzq4epk8O1TG26rSTUcwUB7E+XNTcAIgYEx
E7z9H73BDIhC2Vapqw7C7GBphKAi3iFMykQrydHyNLJvWme1Olw+BpVQtrBgz/jm6c5fzvp2iVq6
r1+bgJsg5BxO7bmmxZiCdu/E9GikokgBiVwWovshWO3RBYLyk/7/an6viLHROup7uktau1rGsp7I
yT0XNMc/T0Vgrb8+BmW4vxgrq5xJpPmmebhM9VBX3TQY1frATJMkaBZ15lHReVJevCu5HfnGBbIX
qMNL4Lo5gHUs5F7448JG8Z2B1jS+dUWJ1yuGNla+xPylg9d9z5zXsUA0/e+RC77TRtlFRJfztVYo
1u6WtUYkhbSKs9r3Bq/QLHfSfNm5PgwEz/p+ksEGSXyhZWPmpbkBO3U4WRrXwaS1/rYIzOwoIdEf
RqzYqR5gqZMVltQIISUMrp3xpIYgO0BSTLOSV6SVS5QbQIRU8Pyi5wrW5OdQ0kCAooBnDtiEv97k
RGg5hxS6QCdYjJZx+WusaYWYF5+bcF1wkrzJWr2f4NwshupZWzHpAh8/WWgkk2MsI3l5u2tj4zXa
OnAUtfIAFXFjA+ancvR1xNF4GKq/911FfekriUwMTKhtjwfbaALYk56Xo2DKSrO9iEk8fpiwCna1
hlyE7asLBK3fumto+lOUFvQcMfvYkI4+x6ZZdHLFaoXqlMl0Qnz5QqZOGAysn740AQLeL3PAArCR
feFL5A+Z3dsnNpNHEp43z2DjekjlaZ0TDSNFVpWR0nRfybmQXwfygaJYAIWtJLNAmVJODADcYAgW
ouq14AdWhCvkrRIfrJo/UscTOiGW5KVUZz3sPd3xDsC+RB+3Yx1s3cseDk3WScNxSbSCKeT1hh6E
mv6H9/4IwGHn18CshvYDuofGY81opDUMFUCHp6JIMoEGvrx6N5VWomuHw/JtHUyB4dG6mLLCYMmo
zSvbGjqDBlFHKAeqc8zeSujp5aGaDwC3L3UB9lM0NMgeUI1+9yYEoSHOR82ZsQ10NMnZx1heeZ10
nJrnVKlLTtLpEjPreza8xTmTWpwMLiIQnxCxX+DXc0XcQ0jxae2myIw78/+nDpRF/ELUijGcsmRf
h4zC7MrNBtif/wbSVlEzvwzZMcxkYQZGEe1EhvQsLunhqT8iZOv79sp7VKiXFFelBT6KMgH9tNrN
oqPxRP8v4RXnQghnDzz5meYRkQelJ7F3aqnoMtMMUFhD/11KbfQmqMoJ6qm3FEYWJARsWGnyU1H4
4hmmPF0vfmZ89RCX9PriUxXqspkvOLRuU94miU6KxL61wO3JnrDJ3gsCC5Ei3FIT1BmH23u2ODgF
5ZNBevcUQ6Y6pTrOHLhGYbkE4gzGO/T5yTUMW27FFvc+wYrEnZveQST0w6IUTsKKnVlGuW2/gml8
1jPyilA9OOt9BBj9Xax1wPQj+AiHfTU437BHrPyVvkobbmeGIZ3dvn3csn8B0HKZCXaY25s/0pgF
gQ5JKP4IiM+jVHjGIJDXbnPi8oLD0sSP+gdkKoUwUQfM4d0avZZst4g61Q3Omdh/2h0AGqwRpQiL
pl0GGTN4GRrcpBg8Wx9YkVD072TtkrUALQDmaDavtBk3uTaOwRed/N9VvNbUz+yvxS8Er6JxZHE0
bF7mpbCHwNMErC5tiieUJxQLq8ibd9tHDWFGKliudWI8omZpT83C1vjUhbzZD0eGLyH3kan5Qqw4
xNeEkqwl5HqfoVq+NLIe7NmaFrhGltvirJYmNl9nXjVg32398MVt2dqVaMNWZznYLZgXchhFsXvS
OUdqmS3DbZK+NQorEC7kt3bBmoTyB5Dptgjf2HeTHaCCIWvj9c7+sm4mugG2No0TFA41lfOXEcTE
m6OTEHQhD47u/Wbo49jgJh5kuWtCrXslNPMQn/xEgkJfVaUBHgK5SkVzv7d5x4CclV9qCcfN6vWI
PtHm9Wq38u8q1acqJgQJc6Mpa1W0+yVPGzyowzAHzQxf9bagetCx1H/IYjdl24GBv7yh4ZPCKIJ6
JddKkQr3oSGxOps2AZnlPnWPj48U20Nj9MKqqW9wvDUOw/fXhzMiPkm03coCbdIeTsFCkHLjaxkA
/jV3MkQC62YSCX6IPpxi8XiffB3AoSPnNl1lKzYN3BUpEif2PxjupItPu38J6d0l+u6JoXoEVhJV
N37OEjI8X78tQxYvWv5WCaNn2+G5onjqwCfYtLfYO7ErtB2fFZGI92svNvbf5hAe21+XrooITFJI
AgaZ23I+xQ+L71kxpzMUlTAsUPwmSRar9D+uFmL+EMwwHRNL0aep3bNQfTkPL4YP+MwB488ABSLi
u1TABfQZy+erNfFvPniD1WIbR3NUi0gkyu1qre1Et6ljC7duZ7GeA0zt+9glb4CO8h3AgOJIDa1D
6GoTK/pxT/eGZdSGGe7JnAVezvnfXE/rz4/nr6f0a1jvU6iwzHiFrpNwPmkqfvix5YqrwU7k0Qns
icd1svYRxbYkokosvXo0XdRdEMhBfZhi3+SHWAmevARWt6G3RCVt8WP0GzthGWFG2CEYskVOBzGo
7zq5BKI5jtPorm6/Pz0YMj9GETMd2903uK9J70FPYuvdSGgkTl9uNp4BcL3FwXoiBCfrsiM6CiWp
ciefkjGxbDbRuGIu+6P/dWDa1qQMp9i5Mz/lIFGVf+REmmN7ohzOkdOCF7oFYBqg5r1QAtOPPjbF
zz7l8hOJpVrJmntOwl6W/ZP1OvBEliGP+CIOyxVnBXb0aZWOj57LTv3dgk+52+Y4gwEiYKmTLQZi
ubCU3HMHKKxMswQBLuRDwUlKcsAv5ujarhKWWaUt9bgMaHXRh8JtPT9Iu8zH1sv4Bm0EQArNk85I
3Q2+IrcYyA6RVHmOMHMsAPc0zTLq3wdb/HELYn7CBq2yVJCPKCOI1xO3mfMoZdoZxr0+4yZDKcsJ
UbLZig+c+nK/8ktvbt4EmhA9q/ag91T3V1dAUikAwlpJFlX7IIU7Apo5JlXDaZoaW/4GMM/q8UE4
IPP37e8sMcODSiBPc5t3FLeOmF1Gce0sYECLjb5r+eOrqioBn/0h8fg+LIODz7gPa2/4p+t38GBi
Y667eu/y0dx3jLadhuZnRmX97NlqSpjrgvrdQw/DLeFcbyVwJAJgEGj3xaGyOyIaxI/rtlQAdKx9
mjqRRPeaP2POPZAIS02g3E4wEmTCtf+xEXh+jMWThUJFcY56sYIuls39Cikxw4PVHMdhWhbYMLIO
v2sCXFMmyWKmpqefwXIWIxkA58KLN5+l9K/yVtbVkVTGuGJe6n3c5SZRrx2qNpFwAER1RWS8N94x
K8QTv/KraXunc2qBRmPkAIS217NrDQjPhxusrqRj407ngMSVht/ubbB1kuEJ+gb9d0NT37YjQGeG
lnoiQpzjPjLANSjy4jkT4jQNvbfQA7BC6D+dKnMwONVuN34cdFiJiWiRw3cIdl8gRMEo17F3QKbs
1jPbE0P2HGFSwemCR3LMoiwvHQRsVJU3dueWxsF20hr3B+be4Gv9thS2UBPxn30wXhFqYp3xSuxP
9aeIREpsRpmL8eIeduO3As2Qb0FXrrfcZRlEe/M6HKXOOXmog6KwU6cPQVgbVj5ld8Ij4sqgs1y9
a5JkRlJgaZGsYizObP9C+rkwltofKJq1yiYNlKmrSm7Ji32rZZOq7tTAmDtqwIj383BHPbPop8J1
u1/AFlcVj01Dfg5JXLlF6srd4p14NdF7FVchgmbPA0L0QMeW0lcyMkY+usWUSuAd7b+dljvKgERi
uN53CKz7XaQQPvDw3ZJY5VpTadRwGOTijdByMA5D7AFZTJgpZzPS8+7n+kLp96xn3DiWpe8A6slv
SfhW9jkP8LAV8brlG/aNgxlem9oH2r3Ryw9HXMPCmnhsC29BKWxybkfKYCqmPfyTHlNAy35G275R
XNMuDDA3yGuAE4Qt+JsO1zX3ZeaWVNnhGS3eiKI4G4zlUnwdlUbeS48CGdASO8+5zCOnDtzi0+nD
cgMWPv5ATTLcQWdv8fwqLmFUg+6lEbMClGI8r4xTgodS0VY4ETEU+hkev2oCyyNpqPqR7Os5MDWg
IhIhPnuP5ZnA3GK/YiJXYm7iUritOvRvRaBLP+HrI2f6qsltP6XE9pHftThNoL9U0Xpo6tQjNSYh
tIYmo+q8nWLqPHOFkuq9KkXkI2BeLr2tg7KfEsW7H+eoN28D+AcFL2NnVADdPwpWsZJahsUZm86G
rIDDyJ+vlqR1AQuekFHuMV9kpB4pFgMt1ElF4ZwDiU3M41YsH93VjMD/qMTSOMReQsAIAT1fhWfH
QuUP7Lj9WOy966PLA9jBqsc98pA/XypxtECvftcxCydrCA42I9UbT+4W0rrG63XZC7EPQSNroawK
kFfNhFxiRu7vVXdY9n8e3ZqiGYAy3LEd7kB0oWRmxjolXDGnmmmHhdOL607sFLo9vqdCeRy6zi6s
I+SLjbg9IMSvSTdDYWTAwnMU7tGSwnRXu9AVN8keA9vpM7Z+IPQIWwx7DVtrrwHbjzyvk4+oZL/B
iXFx+z2guSUQ/jYXTrX2VBotndWTejSiTh+U0y55qOe2eMPsxctpI/x8fkPkBdHiv5ZuV+eEdMI7
rXRC+jHvbiBZ5r4aro0DF5gGILTGeQ1nPT9o0+9t2TNu3hhQ1c+TbT9uXeR4/qfi0A0b1eCS5fBz
tIY4V5134Phc1kftJcv4J7C60m+IH7meeiacRgOwlZD7wgvUBaPfdssIiA/WbuL/UxpuMo5PTrcm
lYafZUAI+cekpB8gffKUayBa6fHb2UjIMKb2ux3+vC8K6ve2X4R4jgZtBVp64oJHN4dhRvg5JDwQ
4aWbyrGVZ0tpFITzGEmZBi4aodMHV5Da4zX9efHi0cadoK24aQPY7urg3gEHosfUhQjcNZ3JTMDh
V02EEED6/v6j2tX3Ov4TBkRiO8rJ0x7kaoPSPSa+2tlodh7Lx2unq5VzwtPFbLWDFd0g1J2zlAOk
Hm74F1mutURAkM6NLq7pni1YFXzNNtS6xgnzOaIgbTmmHL4WGL8KZiWO+R6LE0CQqwla2EC0wxfU
8AIAFkvmz6+knTyvnMu/uBmFSbVYmGj0aWGtpTnzjF20Y9m3481JxuOQaENl9t8JsjywzcEbWlev
0ITSG7cXHhUVrC7t1VGgCJs73WskaOOqci4pykHpvYBKENNvQgw9sBZ0I5iwgWr6ye5+4+5epco8
jZj5tzFi9fPKQc0E3H2C4tu/MOqrwO1yfLjdwkytytQjm0HCPmifF/usdDeeTUmha7tGZI5ixVzb
jnshi3IHr0EJtmaKEbOwlaYoB8cqkm5ZBAvb/nEmOx51lKi+w8w4kYQoVWT/5I1E9dSQBCRtAfd8
OAYefidR+nQO/cVmm6HuV/KPCDBh7Eb/KZL0bCRQ+uZwGcp8zfEvSd5iEMkRfOSNCv49dBVV9Xo2
egfz4qe8KhWkgFk+DdNvuQzkkrRnIdaXFwnIyl7Da23MCHls0Mfr+MCIcWXEqA2Np4U6L53nLVdf
g+U55ecRSrhOAgpOskwR3KrqLE9orBuEJ8kugxlx3Xn/4qBQKANIgbBGzuINbq88iVZnhAZpluyg
LhkZ8gsg7rXlFDRELq4+92ltXjvZLCDWHjvBW2mID/0GgFzVTDAQ3QzjPVdopaDUhmX4zo5c8en1
gIVUQhALegcwg/B20hlncM8vYtEcAfrHQBzbFmpNFTKe09LQMCGUsEuabSAtePWqNE0si2VLWsSS
7q6wYiUbLDkan8PhYa81Wjb8GZ657aWn/YYGLDKymY3ey6Gh7TVWFkbnMUC6MeKbbhDiGftW/wz5
kw8rnFAeRTR7+EhP17CUSti7JSauajPWDc1agRJ7y/nPNoa437+wbvCKwx5Rz/HV16d919EvcbYc
H/2TzGoSGMueO55/sotC5m1jvyDGSDL9eVpPQ3wC1te4XtNXIOiAnh2jF6MODyeAmJTDu4CTaw1N
QjaiGom0CjSBctvmDHkm1HwgmfRVXya/O+xRTQxEes+DhSqR4HS+Kp7hfO+nTZy4JYWzdFOzLpR+
phM3r7aZ/ekkWIA7QSKEy7Ed9GC3gDI+HJgzxcBnWK5D+EihqFHzfr4bxsZ1YdcN5gVmf0Obfxpn
jCyUKLmC8SWCe5K0X3YJdj5KIdyd5mD1OBrMiQLBpmBxr0vlxnFWiRwyQ0LQhxYJJ1gwVHzC/9RN
j3xg0L11ZkXKFOgdLJRN6w7nYZnChRnr6qATg0Ng5RYnRsTQU9bEhqufOLCTBUkVieXqAdUWvkCL
dIAVws280j7Z+3pbCtPs/bWcVqVcNHZeDnU8rqJIfWLjtVvHoRw3+4K5Vr7yMOHzKHal4QOC5oA0
88L5J50Gu+gLXGvAcLNAx3MD543XXBcW+zMU8jnB2WgG1ip/zKQZ5mKNHLvAppVezsGK9mydtHC8
P2+T4ALOisB0QrxRAg/DaOMuoslkYKqR1Rod76P8zMLB6eK1HHrg+AD9Z+DoIl7r61+hedsZShm9
inAiS/f+FbDtK7SJFMRx7xqrgCR0TIfNFW9NRGtgR0WWq8bCypA7tew024T7xP3H7f08h5rzTDvv
AywBxQohfQWyKIiWdhZYO/qmYGy9kCEDbcqadjbtd1Q7gINYtTPQrWqjVbvz13G3SjVBBgDRz+lK
MVSq9DyJzAm9tIc+H9EcGtcv6VH92URzz+CFEAF6PUpqDvOb7HErmHRKLwQJSMY9SDQKVw+QIO8r
FB6Opb9ve2DxK4GXcgSnNKTJkgTs9KIUaGoPh1aBNDazujs4IruL5KVzezdclqVqf/eOy3rge2NG
gx/aBLalnDyrW6b2eMfmAiWI92zy4Eri+xCbRH6EFAD0JuYFzdiqdndPxxI7i532r5IHnSpeknbp
hWQ/TjwTjuR9VbE9kVEm8y1OmuLPHWgQ8O9ga3cvVGWgrhr5d57uecqSyY/QYkkmU5INVgiH1IZp
9zBE6uTeM4AlbidVfcfQ1e48O1m4CUlPtFhBO9s1Kw6Uj62IXF91YN+Cpa1YpV4tqE0fZTg6++IB
gknn47pl0q30rhQv7UB3z3HdY1dnAa5BQE+9sPbCWL1IkwtKJuAV3pmAyL3gQlSCKqHHzmuxgNsk
SqAzeSfMuXUC+HqktyFsBBN3atYLGwwCO1ES3Zjsz7fGRacJ3Ms6ek6aolavBckP7AAHGAcEashg
7yHReXwHJUtQHPT/Jv1C510PXFr7gltc4VEsqoCS86NrlTB2B5sLB/odSVODQ+ZyBS+rwEaOtsxB
Pegz+ZnhfZaOhuF0e5u6xCkhXotR6x23RPYZz7fgRu3IUhnzNyV3FZBd4v6NLgRkkJgukEENImUb
5r41NPm6lKzG0ib/IY9DoQ5s8E6YfEfQvhKiqBnSEb65ccvyo6ebabPGTdIw2H9UB1Hd78iTAGWi
umX2+UlsHROzkV606K4r1JmpNS5sphTHF/F14S8BfLAPIrSrElNAD3GfIN5ejfRASnkx/YA4L2k5
JHXRP0savl5duGr/+te1oQLjoDYe+dlXqycpM5IFOhc1XpQyexCw+K+s8B0E7ir9jkqkFYUFn158
YJIG9YcV7dlPrl7AijsNTiEqCPoc0N/3MRDBmnjXZ90dpeEYomIftUt2zxj8H9u5jqWMrkBkDwMN
lFZ3LkvA01KFhyohA6XKIlnKEghQ9hJ8O2TnSudTPyAAaIrE14h7JiNHhxH/NWtBeYrA1dTdxhsZ
QZELR91EXkc4sGjTe6jdzxKSPJaYcRHMUY4KBI0jpXJ4wpEB8PMWx0cpIFHBjirV6nO22Nc3mSV+
Fis+gHLykrdhyB2NYuedEmK/a/6kUBomuhlMOPduQRQyOEL5pqJ03EacqC+CUF0d3QjORrjMyqoa
cXTuHjPQ5jO+vN0CpV5CsD/AC/9M9SPT0auIIJg7O0MvDxBD5iHCtiXJcV6Z+IxX/lzNqmzOdGM5
Nxd1h4CuF3b22xCG7wDm5Ozl9QMZ5zmyFTiCOIMFm4mIH96EmipVnF+bGqc8jjPvgErJWjkUKNX5
d13lte1np25pZk8Yn/vE87+lN/o7KVdhY5ejomfbqWeGlCr2r7drgRL7KrEsQUkLWoZ+BoSi2Mu2
SiC2yTxHRZZdFmhHn/ROS+8z4q/lysRU7tkQezP0+O9hkGF73M56RaSLtzJahkgSA8koF72Q3Fqq
uvxXQLcDKZKbDkAWT6yBqdmHhKR6CsdwZGkvzq0WC3Wg/cUSef69G8EyoqwxdzzYIBCJ1qPZEvfe
0gOTo8IHDo/DsUssdE2bwAwC52PAErzS5aa1kHR943blIU0wvdZRHVBrHLrLVdqxdy46V1LkLujI
g9IxcEeDVgN4tmQhVkgOpDbwJWC5CEShATZPatUDHrp18fO/PuWdSQs6BeN0A2ugxeSY7r6PQjoS
i88Q8EBo3Z7U4dNaT2ro+49FGPzPRwIdvS7Wcgwce9Dnc98x2OywtaZgdPxvx3ZqvHGt2wbqsCK2
56mvBiDu2Mu/RmAwv1OL38NCRAVLDwfAvTDbMKlReqeSHNSMDmWGV1CHJmunGrSLXC9+TZ1YP01W
9Pc9+Ip8D3mUiOyELbBHlF8Pr+kT9GKTsZHTqzNXg0Nek4GLCTB6hsPSmFXrsFVt/k27FiXtaGIy
WqeujM1AOMG5CZaXT+2xR/4g5yW/tnUL8Nr/onIDfTVHbwr/rCpS/mQvvt9RF8qO7Mns0CdX5sVS
dRmR8dWACx9TyDttnTFqRM3iVPxrNe5v0LSvJtMjL+fiilUEG6SrB2v2Uv0zZHzj+kJ066vq3Qib
bCmVkSSSas97xow54IUEGzQm1riaISc1WbOK508BEkcUp2hblMiIyPm2OEG3LabPKgexPc0HlhmZ
lvmszMWN1vDEDhWIHqAB4cob8Mwj0m+sQ60oxpbNMqLXvRgmrFKKuVuaXthnetDRljGRg9GUIXhq
tdJm2rYH7p78tDxtGfQmV4zZ6HUGniwEduLbn783DZIQk5pRxMWO0Zif7UzYxvBtofhGvin59fpl
9N3Jw6/wI1NIQCu6L1CA/6iUGRGllLcTCfhLz2pP+ucL1WzULDqySYjurMezOZSTIUDgEn7yGpCM
rHB2vfKRZ8SZ2TnHTYfZZOmpXUtdpa8pYUKERAhuGWzpzOrlOcHPG5yOdga34IAlgXUSZXdhJklk
jK6n6g2uZxgQEnfM43GgiPWzCos3qYuWKBiN5CZGtXKlg28bAOdfBw2zTtKgpeuKwKglr1FOHfP1
CjytuTl/eNHqbpt4HlWjipj7c8Rf6PyCDuvA4lwL/8XliGXF5Sp87F5orsFOzbHHCXAlHFaEr2jk
AKceL5h7usEUEfnfFRBOVM2NgUdWiDTPlEDjnctgQB+CswRUHuRp7vgsD46eLwI044Kr47/4sEoI
S8c0GyGH/Awso3ImfTOMGjeEKWVIOh6MNvWxXwepxhWb+tGpCzcvA7Fl8RBYDCukeWG37AWPHzJV
JWZpCXkKK7cHI4DfoDcLwNYLCNHcXBPIOdL3qklSB1KEl0Z9h9SY7HadWweLuO4G2+/kqQ9UKNhv
KeVSiENNqw+2MEcViSiL8BfQNOc9M+j75h+yLyQ3AyjCcWv8pYXueNetsGPgfLMbhIJH0YKB7jKv
/6gC2b7lEbk5miCCC3wa0yHx7yT7dZh1N41buvmMJPvoojvoZNnZz6DzmJW+o59Xb2bvdms3hVmx
B+zAYy7SbwMe+kKhXJs0yCTOPDSTlfTb6zLxZ+1anJVY+T3U3GoztKu71MalTYYFVmSZyByQOOqE
C88G7sGcrK8yJD1uopjO+J49PFBEqfUAINqqvenk2B6nEVG1ioWy8rqK+rjT+YO7pIXWXnC0baQQ
jw9nc+4rwWJ+8xYVZDBouzV4/KT17R7dUNfzE4zNPWlSOCF1DaEqExo4iM/h6SbJOZrToC0SFU0W
HlOGaprR9JufR0g4XV9Ys0BPuLbFWEn5aBvtauYM7K455teky7r0CWCwSWVxrvavyJZkzhesY9fH
F3A6+CZY/DTPJSCOf9zvwpm2DBDBtr0P0Zcq1pD5iXM1paN1pmQV7fy3BeayQVJNt3fhGwexa7cV
pBj02bs80H6sK6QzQF1NXQArkcPvcOxpG7Hb5q6XYfKkGlrvLjGIQFjLU17Wtb81fXaTnivuHShP
XuoU/bxaXi7a9cZDdv+XBgmty/Y9g4d4DazFhrYOtJ3ndaaQA5GL5Jtlqui09aONzZus9hDotXM4
TCulszduvAU3H1pGI5RmmbfDN3Pm8CeIxBoChYnZNwEsuuB0DLOxdee+rfsJfwYCw17ypWGVFHvk
8/B0MPCLTVGDjnOg4qY/LGf7Cvy+VZKLDaHsgOcZcNdPWOsEHVWGZ0SIa4myNtq18eYSwSgwX/Vi
rv+A4H/jsaAbzCMyIhVHrvIm1aJfl490dwrwtlvKDmIpY9VlFRsstsUDvkHLfPFBxZkN9k8HT+rb
mjMY1rMQ5dxggpglVvhCqL89KqIE5r22Ty0CaXWcPc68ppYzTUuiWY7PT66KFhEHyvGBoCSAN5Bl
YioN8O+bXCQSPSvGGLtZAfzfNoWrbInsUYHzCYXC5WNHgM/UPRLhMCnEJwKz71VhHS0OremkdZUL
9bTcM0689GQdokJ5TKzemE6e38dNhuBkqe6JHHs0TymcE2UsH0h4cwJB87U/fQSu4nw0kT5toFxZ
53U4U6mfcKkvb1v8Xg2ZZQkAPJJzKpB1Bdze1j4p1/1XIqMgH4oCAvfKPrbOuLkFt7+Byz3a10C6
25ISlTgmzx7LOzzgWE9q8pcM/109aeFvvSh+G/0QlnR37gX3oPdWvTB9XaELXUkkh8fb+giVt0QU
dnETxdt6r9cztxn1VT/6oLB4fctawH0ViN9AAlqCajOIgBRDEIAmXsItj4wqHXxNSd6uxu8thAuX
C4qCP+JpGSTs+2EPLBd2hrGRsJx5jX82QXC1daCzX2hVYAOt6l91UyBvBNB2xfSpyPzOs2MUQ5Sp
w50a1c3/BXDi7ZavUD8tUfrtazp/zHy+aCKrPjjy/DOsDxWIMM9HaJ2u0RqNavXZRSBc/UJJTP+T
a2RCzarY5XwQu35FUMwudbJ+brNtAfQWb2i2V7JHQ10pTIpIwBt+YdRVoDtIevuonXv2/5dd67Wc
nYd4c3nLGOSlJw+vvNxoXlhdED4BuyX/EKclnZVSirksPt2a82rGDhA3ZAlxr+mY+hzRcfKKeRnh
+KxINV43Yi2seusumDtb/CsuPiIzcHBzoPsiaUSj7sGwitOHwjAUDsoB25bnYQO+/+IMMs8CkN2l
5+ULEaPCv8TNOlaV1yCy7QKSQhYXCIAz3CMsi3U+rWX3NYHp1YLATM/W8FEFehtTtUsgYaIHip/4
5KV5EeyIApiGZ5HB75860XOqDvhcHWIAdBs9XPG/F8MOxwSwKTarWzEWHA2U/DUbgXE7jsbWLKIC
v0j/0pZ9b0zRjNO6fFNj6RSwq9rsclURAkOIMQ4wuVJeh/uXpsjkTrmefUIbQAJMZ7dwcNBw4EkF
F8jmgGIPMBX2d+NpcrkG/MoYgbzBb0d0jvlQ942UsKfey0GqB+43pGf1EV2kKl/yFhCZxixZm07R
wYbf92nitaSSEfA3pb6Wo6CG4CHsuVaz9yVGHurXuFiHlr2rp4NMtswfqKWxBFhc3BKuD+Kh0YF7
x3x58W3HVz8CKUjeZ+m7lRoVFqQaQ2tWHZ93lFe3XqfBOW6H9pG+ISHQd4AD05mUQLn8WZbpzLp0
CMC7+DLnIZsnsseQKpD8IGwpC1mvZzNalPR2ntDiQSaXCg63xa8GiExNXyEA9alChtfryzzUowEO
oOMb1jGuYfjF+Wjqyh2QqUveCoqhFJvkf+AuAZ4DGfTTS2PeZWx3o8WCoxeCOTK17Ha85EDp3NHq
yYYaOSghTT7LZicq/zQm6rD0H6C1uNeUmWitPj65de8QTF7w29GqIRX/+eDysAqLVnv/f/m4xKu7
O3tZKkq/c1b64Vs//ETm/47J2DXOSKq4++R7MKj298WG2c0Ds9lchtlvxuGXA6iaG/lAbAo7IjkO
WVY2O5JYI4b2bLoK39gjQ/5nYe1APYzpWioHPhyLwL9MTw7mjFYaZzObAnGW0vhYBjoAudUmufkg
sxSoCYd4AHi92j/QKl6PhkXB2cDYxeRu5atQj/e1WIX0UQO5xx8cbj2yoZQK582bnO5aUfADw7FF
K0FjHd7g/+jlLdQU8wnyDQCBACn8qely0SogrFjDMLfx/GwlUwLrQvabOozfzbijuukmVwlfXE+r
VaVGm1gee73waMM4AOcpJkA4LPsWZ1vyfxoxd1Iw0/jS0ONS3fmElvlpOTLkQJFr5aEMQQKWnWKG
GdOOxXAcFhusrFTCy6N9ZqOeOvJW5k29UpXQri7EUvU16JV07cEMgDcxr7jbeokojBK75Kfyl4/M
qTf+b5cEZEBJ8wyVGYKY+9XZqsFLgwqbltHA7ZxfZLBa1QTDI9mPS5otjZaYEe9DtJYunFkiBGiU
vEC9t5scn45NyQ82VnI0XT+T5lqewTTbGUsPMyMUy5H87pPPnwPnEfHnTOsAgm8tL/M3Td1WhcAE
svL4eo6WoIgBsnyp1CtMhoopvvcOMmsnPgPm78+wc4N0+lZQamsbBNQWPhBQMlTK7TUjafuz2grC
H2dy+RHTSAn835m15PuOqtm2f621htsifCfDugadns9GrNeKKIn0IUXFOQZC3pbECz4rgq0l2sna
qgB59ZXLlb9hvk+TUJH3C331cwu9sGExZyv+kxdOMzmnsfOLjJPnzILPdswEl8LJzw88SrfVPciI
CoN42ADM5caUxmI4e93td9hxZrcINvJpZLsTnv69wv4gpahtaJv+0SMRF4F54BjBDvxMQs6f7Seb
Gkkus8DITaeOvTTy4I5Tk5EUkQec76rdXuASMrvDm7kxPTyba0uzDxGaR9aNfLm2e7fp+9wp8shg
DiDS5kqiSnb8f4/DcBTL5XGZGMwQpQ+MWtoDhZjemUnQ72dPX+92+9NosmGmeeJXkBSekzUszfK5
K8PTh+mGGP6AYUn5IYgpBQljtkogmVZTWWfFrfirAE6jippAsCamM07CUcEvXQ2Crh4XRlSbJ/tF
I/YXyonx/O7t1l4DzUjb+4AWYGR47wtZy82uSg4LgZDvJ+Ns0py22kxKMjt9OlbU6jl1coCuv/Co
tVcm+COINN062kWzlCZ4X3fdSXjsARSDBeVQ36/3HgIx6PRdlHNrCW433rIfKi8ji4sF+xNKoQlP
zRulSRQpRmd0QbvyP8dYLBxLBPqKFDgVwbWp4yFLFL22uiNnKt4Ju7e5+tCakUEJyM+cdkISB7AB
U2CDardFzQqINsC0j8sohx2z5nb4+L79IGhD6kCLQ2OZ4Weu+EyJmObJUGyHBo+8Cthe37seRjpj
3MsiG4+AifPXo75jar++jFpqOBs0kIA7uUun09qZABqq3IGcTsaYqDDb9NOTPI+Icp+P/QBfD8yi
fSMCiD7LAepIxIDpEUTdVUmZXmhEAZ4CJaHWZOMojamR7OFqV5jW2DANTMIl/UBlqNL9zNV29aFD
myxtx+qdFbvrdQPSx4cGHzjFlymFCFaLcTYGcoN2/SU4vitA73nm/qYGdut8cvqcd/mJWn5vaI/h
bZxGrsPOw1x95eRfulStDwWLzcgz1Bz71V74gW9BQNkMayzJ/ZSB7GbmgDVJ11ZQ8P4gUdBkaiLy
qIYpNUOykeSKKwWffbzCZtFV3QGm9oY/nwGBshOfYmv5Y9rsHsiSal0MJK7mwuC2we0jB5Eddzjf
WHvWzdPh7/I5hu7RUWE0dNm3nlHcTFFHEXAD3D3c5dorP5rnk0rHugaAOD2DRrbk1v6E7uEjnMRg
7ye2OZKwvdYiTIsZU49GWm5vx87oGRYukez/CqFjqaqh7CdFtGam8YRfT7SKxbhDOTV7ehTyAr8y
k5PL2D74xiAP7WVH1lL4yJq8lCkQGpZNtBGTmp2e5SWazMrH7XLvh5Wh18N38yVmnDkOJKo14qV+
rG2/FG9KT1Y53It1yLXcnrGoHtHg2TFX+6KsVS1KM7XUJGVmDREaaJYDPgKy2KVvERy3T4qiOpTe
hrLqAjZVoRP21qj8OXel+klhDhV78afGuLjCKWSdw+Xh3XLO/zwMw4oqUxI55ilAFb4TJVe6J4lX
v/eok8Oos97yf5cIlwG6IxlRS7uhlG7YaJ962G8dOJ7tyPqOUepQILnSh492JvIWOPp+cnveBaAz
USEIT/POM3qBHtWjlPx17SmxE44g0bk7yfPAbMPiogY2AK1e7/ccVRnZO3DNVHVu6MGfjkvA43Fc
wsetLaHeikzMNghI6jiY+YLmSji8iZx7D9YzZ1VwMFXgPDMDbvWcWBCr7ux0cLmPrOhiSLMjB83C
qsNc3QtvQrHFSkJNBUe7kx2BTsmvYohnTzvbMMlo0MWPI6X12pkNRX96WYo2Zadfl4dnK9IDFw+O
teTMspU1cbliGj0bhayvv/FMjBDxwSMHy572vL7kwWfyIpb8rOWy5iGvOJkadZjFsFKQQ3Ztb9Ej
P3yFALKo7tjinKeM2TYMqJvVu5Skcntddc/PU4Xjvtfp4ns7PbMy9Rq2CWFUhF7URCA6aOk5sy6S
CU4f0lkREhElnDFO2gT0TU9inKWt0qSAidj9RMJWrgvq8g988KYwLxROBzbSESOSSd2WdX6XGA2T
ADz2/WILVvbSh29d11BzZLmtZB7Ey3KTX6mmWP99aGNBPeN0x7bxv5b9V9W5pZ1fHQBljxsiifa/
FSsOpI7etnWk9kxMkr7in0GIpbNo9QhXieLFo8EyxRxAfjI374bY6CjCfHXqsMzYW0XzYW8+CsTB
aCC5MDT0kGULH4VHgSKxyTveUC7R8oelJXvehxQO0fyynJC6iyz2a9UlL5E0HftH/6q3tkd0GE37
pQ4c5cVS6Uxqvmp9udn4Yezgzstkmg5Tq7Qq27Pe7jQZtsDbDvhTIuugECvZ5B6GIGWT3DbCo7vh
5SiKFAH8/GSgrwDA+iey50iVpyMf8ZEwRhJPDYiDJr1n0PSARFViMBc398WEHE527aqqwyc46enT
Iacv1rsFgb1wMnDudIqCvDOcTa4xspYQf0rnLIXec1PRuzVbNVWz20FD5pYadhIXhwA24Jr0s0SY
kf+DphPVZQPcgMN6N7CHwSOSEi495KxkItUbACrJ5Tg3UNNYeNNcMCgXGSXe911fqEIKitR/4w0c
sMrebGTbSQbJsbCRzvwwoytu+WcjghCEfpotfvZ6bWIfi/jqVrxJu+XcMJt2kvJhforefZVGlSzA
3LahB9XtJdvmU8GnxLp+KYtoeFqeNpA0nRMbHBD1id1G5X5WDih+m9qM4vK6HFaNQMN/zR3YEFsS
LhdEL4/8eqVFYWew4N0Ux5jmc6+jClocJWc7ZiAwvSUkFrNY0u3kHxgYfQ+P/W+J8Vgzo2LKx/e1
veOr5kLWHxwBfueuxZRtSddNY4vJSaxgr6tBIO582ibzh8uz0GdCmH+A1Z/k3uRpd2j3LYYeobsl
jWFVD62VjcsllpQUtf9TDtoEW/HIk36pyjYskMOOYnh5TocLUyJ0EBSKMwRrWBdld5T85lAihYsy
sB+vXoXbX95iGANisnL1DSvHYD9Hh00bf2E3fHrnTEPKk6NVH/zd7MuzU8+l0BrDz/Iq5bW931/Y
FQp/Guu74i08/i5dBqx57CRmEBsWZ0/BIPQ6RKs2qpItfVSQ6Vk5WOHtCL//sMxTnbzUfe7sXukk
qYGL6m77zOR6gSGUrjufLE02K9WaBiybCp3yQ8hCIehciCldrIYRjEUqKplh3QF0Eh1YGSIo2nrA
E+YsopPoWmwgR5B5yw+el/48w0lOFyaRKShQbuTMCqOADNHFIC6cbxydqAMucOULIbY0SmvJl2Ti
noyd2aVZ/E4jwusnP6FZp6Z2mdirhF7ub8LQa3jWC4LPR7a4Rnh0euJD8UQkDRnQyEpTN7wxDW5Y
VsAQKuw5A4c64GvtjVvAz/+/v9gRv+qLu0FC3Qw6X1wGxHXoUuUfnLisLOeX/db0fUqTS2YuGQtk
6gAKO0qGoCxRZ6d1eZL0ZntW7AmzK1rG1t58bJt+XxXsOXSIwi0c0bWeorGLgrkA6mbR4WjGsiJt
KimjnIdohlpOS7JYMtRkICYHfhATLkf1Bv0pe5H1yNdONK7AjiV9BvoJYMZcEqw00fHqzTMfXLor
Q8YPl9pKYMCk/Ab7QR/0K64/Ik79kb+rCjfa9yOixiPjR12WmDzKJKOEIyHjzEBrkxg0XnvhlFkO
Uzp26UiC1yCuhI/Bb+o+q4IIqcPKowvloIbyMzA9eEzWpxBj5kExpf7BNbWtCy3KGPfiyEEVGWhy
pOfUvLLHW8aWU0LUr8N1DrxHUWSxAQ83jwBDW0qaocUOUTBAFz/FYOTJftNDlfyr+DuWxOWACz6r
dwNKEexayfl+vSxNz5eth/mvI5VnjJAYTxCqd0HzDJQz9CDLh3fKEAxPGkQqJ46otaqNleBA8WZW
zGTsgEVoJqmCXbYlO+9h3A1GrI+kymlzFqLV9IBFMzvyYBrksWur2qYHTtMcL/rt4j7UDJ7U79aW
eHDYvP50XTWcKs13chFQYtrVuyvyFUDyiEQy8woVZAQ3HTNUph4BbO1UocDDv8p+RaSygSQ5A2I8
8LjTIT88QFkp33F9JmdAaJJBVkuwftzja8LmIAtnTdXmHVrQFJ8+SVL6lxzfpzs4CMBPK0RmV4N1
w4kCFNcIm+mEWTZnpKwbuZ1W0RTWaNwZ+FkFUI+koHq9Tc+M+qkcZxL0vx4d8AT/WhQUVL1il+Mi
GGURji7GFmnQ1qzWHOy/LG0vQVSYqV3Op5AofyuLslFPWyLcTD5lVfyc0IH6xNhTZvW15em3MDgo
4+ucNT4ff/3hv/Oc+I1SiaD5FVM2eOnizzf/RNAPG9WgmrBVLN+LaOzacVpnHKikzMlzXbJy8sOZ
GYFGdWS/sfKWqhaWiVsEoLRbV2s7fLfC0xg0p2SnrYylB+C60WK9B8ZE7eY0r+ayJmFSOGcIGgnT
1WjhnhYJKRuo39q4M7v1HQzebYUASYR7+uEisbd/lgcYHw3OvLNeScR+jKdNis9cHLntPcb3gc0M
HnVb0NiYCltI/TdLHFsPxoxdRTTYoPHIvjX1L2cYK+lmvZu9aFPzXNGqJ+88O8GpfL3o6h7wvwHV
XcowFWGMZzO+Fy2OQCCPjiSTbM0BeIHBqqIToGr7fxOYoeOtpb1EI8l1HVIkcZmmj6SQyBh1LHc+
g7o67A3qTcNuNdljbEKAqRMMho2vB25YftKqqz91SWSMlDt06r6HRlcObrd3RTWt2KFw3eZbmHX9
WjzYG9NbA7wMfpFkF9o+MXwO/aM2ZmctoWCMBn4QQidTjtYRl19yYl2PdQ2YjYwB93IuRQkmhx5H
I8WznvfDK/lNotsWSR6KmCnRnceX2VHhnAt7fqhvz8PmOimLg7TbdeO8CTbxOfPqK+OFuCoCiIzn
CpkcXRtxycv39z9+UkqjXGq2Xf5z0WtUcRTE2W2gfNvpDSsi9K41TtXuIZxfR//CfsKJzflH1M/C
iptE8m1c3647qsTwBMI1XeJwNGBtI1na0m81LJ6Ia6HY3r7JxtgHkVQLGGJZ1EHIEHp3P1OH+foN
FWyWX03UMpH9Riaig+NBnO5K1MVT3fMnayYDLYxpmO87vpbU1SRKLoKfoGaRm0V2/+7j0Tg7vvCM
isVMqIXTzDiY0XplJPBHdJNnk8LE/lKrPqn456JR96P6doHFcOxKwZAQTDGqODrNmxWxNR5uQmX2
cKgpB82kMCNCPZ3fmi/2+LA6FT/B4naEWF2V64RuD0Q+yijJ7Nqby87f/a5O5BxWg/Upq7BnqerD
bPA0qSgugFu8j/0tjRqW4zAMj3Uabwx1s2F+bsnRAZ9kTEvafb9lObpZw36nG5qDTuubY08REo1+
e4FNCqbmYtVtqZiuftuOun6D28Z9YviA11uWjNe0+CzpQCR9NCfonpfxYcyJDNFfpyVmgGFp7iY5
YCF/aV6oSkPucju7nuJYGrgLy2gp9OHtJc8slryIJsWYq7Qn2uRhQ/xXN+joFnqUCkXdSrJHNxZ1
pWWpPInreipUg085qpuZbIKcFAfoyo0gly4e9aflmjemRPSVVPsCeZSu07l/mC9W8jyzRgY0UjlJ
yUtArxk0Nv4JTXbKnBX9heLZZhwF/VV2+NCd9+1UllLNWczPbVP4RzlfQjNpDXnp0PPpxFrl5rCg
gSX//Mu7iyIYm1Jkdq1HFk8aFzcuaueGpcQemOicApHYxM/2ktB3biWDtqmQLWQojxKufek86qp3
O6GtxW3B4huCHpHWET2UP8e4uw9C8PRLHnf5mCjAmrdEVDFXbc7NhHci+90n647XRw0x5GtttRNe
SmhqF/LALqAB4ZFRWxqUVi/mePhazniZKp11up4g7Jy8Oh0H7gwfUMK5Usms4R1+WqGldIcK4u+X
zJpyQlA7QOgBM4VhO/1QE9bpnDCr4Fr/xgjXVtEiKe1SpoQ4M3hWKD0ly+EERShNSr3EShuHIoly
WiM/HcJHFtLk/2lFNrfKLR7f72idEVwptcaT5IJRFkRzfXvDbYqvyciEKuz8Q6MKp+7XrmgtQ3I+
23w9gtmib80S9qFhabFvKUjbrA0dNkvzkfV7RGbin20/rLImBSFR1lb+R4nDhZyc/I4DUchXXOWR
rW/384ITPmoDLhB4K4A3tTakZb4FHuW9EQNaKa6DSgr1IJeEzqvhpS8tBn+ObIJCAT0dC3ORRl66
BAD2CiWAhG/rs2vJKUdh+jGdQvl0Nf0V+4xvBMWi91ti9x+o8TQpQWfLQ3IGDd2+GtZtJo+04n7l
89bWYJ5XkGF2Zx44Aqo1vvV8BvjpHnZdyXDPvCBCKgigKHY08Zu0jgVMyIv2n4k6C6jBPAIhy5YF
uf4UlcmFTpDtI3Sv3Y5uuxIcIGwckUwxGfKOvA5NyckUy2WH0/7tc5pOjE5EMMDfX7jncwoPHmuq
IhK0ws8nZCTwg95MJPqBb5exrkSL/u0bSa01cBmWVIXlgH/THagW8BkVzcS1HouT8NkboCOs4mQL
Tf7XRRvqGcxFxeknZqe0Hf5mG34d1KokyaAjMluO+w1dLSn3iDb4WyZLZWhjBZm2VCBhdkhRsuE9
wTg/i+advRGtcLI4fvia+6wnxt29x+cc3Mp2pl2dUwMIz0Bk/mf4I7BN/+xPu89h+pTKFGW1eYPX
xr4w3ZA7X2wCKOd2qNRAA6keYWi2wGFzhgpgAVES2dcriIM6KMKjTSMk3GqFBiRiXgCrEBUPkvR1
VD0vNxx9YljDIswJqCzblknCPD5qrD8p17seyzW9ZlOKC7Gx2wBWyYHXjigTDTmyU1Qzh6sWrbwl
M2HQBNJAqp8AKNDRfYaBT8XAMJ1CT5vQmhb1oavTAxxFnBKNVcyqit38YCCQ+hrT3ywVnEichV+n
wANqHI997eUsYkKzRIpxrzxdC+Jr7+zk9kCCjT89ctloDGjap1K3g4PAtc1m3d5jykUvl4UEk9nE
Z0FNnSD0Tq5DdXUfB7MXVsPBQyEmiOiI7AzS/0+mfI7ij0n4gAwpKxYJEYWZnW5FhrN/Kq9tCoHL
huHdjkO01YJJeqqkEJa9LXlr/DehS2ehsQ0zXkudsf6A9iflEpK67dL0BqEsVPQi7L8f1/twvbf6
A3tBnxED6Uywd5Ur0u98dVIbEhi8VFYqKbQft3Io9YxyLFj3kXKdE3PjJaTFiXyDEWCxTAbnI95w
67C6OhzJIMu60BGs4VCl3tmUP/R89iQ7ux66O8NY+FxzvJltCa3ELidGEZSvzdw4r7rON5gr9/fd
2ZrZgJyjJJcmZIOZAyusWrPF7u9IRHXreldR+xNvikxDUOyxueQSZ3NtSb9ntA8Z2tFX9+0XrK+J
hoAmw4L6HP7i07Ai49iE6Ud001g+cKNBA/hcLUxSgpJdhkZptW2LMZqEsoi9cNKwPqnjFJXr3SN3
eMHo/h3vPJrdrcdxp1RirjUHvXmO+pEmWZ55hsJptO9O/cqZK51Bl5xPd8nOxnvYSDA9ZWwU7Iku
Jp0YktAbQiA9JnBxdYVxCkcAJBMY11rIEar74j9XSe/wzt/WreGcVfIrU5n+eKz69LGnbGnSi1x5
sUHfkEuX5Dz2ZojmcvxrNYjRp4nKr4f8fothCEE4PRUzW8uVnm+tn1a6RnyHwDeTDqLGM2wvVnBJ
ux0oA2tTg85qt9a65/PIoM36mKXge36xOinlsaZTUuBbsKx9+nGoSLhrEa+7TWiv2OFf5GIYVVy8
yLCD0CKGnWdrhP/KDUG03tyFi1ljEKybhLjkJTXG8lZeZMp1dCqkycn+lpdinUk8aQRTrAqlu2+F
0XgUoaplC6hCR3fXaoZB3EjtLV3MiPTfFokYSTFo050VKYC63qaAyPCLb0O5acFvy4A7FAPhccZ0
EZHnAZ9pCpwEmPzpN/fv+QHLt+mSwNCcNL1RMh/JZkmH32METpnEkHQIkBFotDaAIvfRVMw5BnzD
Pz8maqdUVXXcxh4gwRw4/gPhISD+59UoL7SrCiE9vqhQaxlFPt2gj6xWojU5y/3UCiWwO+cRXIrJ
YnIT4B435ru134hAI69adrHqJNWeufRIxArGGU2qVqrs1vaRZkbjzbthGWL7HA2JDvWEv62YJdhu
hpRqxzKJ9/l3IKe4Iexl5kyhFAIzay+ioP6e3mwSReGLwwF7WH6ItrnU7B3nsxvf2/LbmGpn+5u8
VOYwk+AX3dTe6/6cClAXjiZv1l/7PDR4rehy8DeBkPY6JsDmaVCaJFf0AR5cn3lDyXFgGUZwLVob
I42lhiN316zFZlfyltqGbKKv4TM/1Ht08GqE3Jdl2YASyH0ZuXLt086A5D1VQch5PH7L/SfXtYt0
4eFjnjQEUzzJ79UJeNU3ZFkQQX9glj5c+hFkYC3Rmp4hXmZJaWESSFkivepBUoJ8XyCi2j5HreED
70/fiJHQDepsKkWpRNtAB5rBr2p5H4qNGNrdWP911ARzzvlGnSF9K3tGCY/XwAY78vSJpT2J7qUT
4wiarX67MEOhi3UCEAb+DHt54cvm9qo1IUmODUcXK4O2S8rHddbjhnaRMUrnA9CedBXZSw6LLKYC
cWr6yO/nQP/GClrYX+v9dlJ+9KPEfRFGM87ymt0JCa0n1SyNiu32SztwhUYVgpYnn2PUQU5Tlpgy
J+6wHiy1AOIpfAzm0eIHQBmQwNBAzsVdlmAOch0A6LomCr/HxgwDjopNrCJAo8MdAkRKFcwCwLgi
fh4IMI627qvf4zOjKVYZeX+C7VxlNtJir56ZYvHcLp7ma040OCijwW+RkCxLXw6kf8y/SjAGsWqE
5H/CvvlSFqrk/07E0fWcMx9Sw/Lf78aEwmtgXn6xppxTAcM7pG6cB/QLyIx9ws13osY1CsMFWzwb
vMIpanmI/9eJLUmpfXYcTJm0rc51xftHMGAJ+GegTk2Tbd/+gZTPatOS7gTP23SyAfVko6nxjoPY
vk51i7H8ZlfQT33Nkl5XFbM/Lfp2Vjn9oOjL6bU3fi+JDpm0NYbgmjGAPyMnOjpqBLDdattJsYV6
6gWKdWRRrTMV5tA9uLqmvLMoTiCzMUrxFBfSihiAXjSJ13LvilkGSgC41kzqx/tSwX/mmv19TABF
LMi7ObdNfDSGx5CZkk3nz1Rh8wtN939KabilmmCgXmYq4kbcNzpgiUV1YzQoA4+6axhe4ETt0lHP
CjE1WHLo1NBYNA+a+ncn2PSo+mAeHPS/18Mkh0+ZteJ1Ubvr4SN+uUpMD89s9p3KKK3xenxH96//
FQwjhXHa7hYFZSNmVhTHKpB1gsyFr4wgdOl1tr2t5ojXJsuBXZTiQd6vvcyOYYyyKVZf7/AYpur5
Yn03z7rG0EGjnixCZnuDBytohmOu8GTxanBRywaK/+cGeFywle/ZzrGVGpwPAGh/aGoPlglwf1hp
SsD6wteo258sCdHYJUAIzg9TtLpuxmhfsgwclLsI3mVXVq01UxYxSQ+9elg0HTrTWwaFx9jJFrZF
NjZ0K0b+E2+eraCo8iaXZ6QT1GNh9f3Vb+PrG7kVqmTYUTMM1LwEGBfsY+lBdLaudYb/nrmVAA5b
HzStSmSHZ+vpsBlzuMIjRHQuRw5neujGUJOwt8M6umLoI0Hl2pX67/2d6Tphg+dWwXGHAm88k7w1
ByzcPpzxnvSNLiQxXeqvbvU50ehkBNDYYN5pR5yKECoEQnrN6lvoi4ORtpKGmBAFwImlx6RrfIxq
SSeTvuTRq1VPcjUFOcpO1fO/5FiebblrPDfSVxVRNd32OkTcHLLTLLwCcWA+CQ3sUpFsFCqDlTC1
CPabREf4+ME7xEqNi8nD0kCwyNpg66Oqu1W/Nhc0NMN1w+Yki86lNaRwhcc+PT2y598Q98GRCR3o
2XOdDoWDWBvADjYFphSAYd6jL5KvikS6rHpH9LxWESfcGT4JTPAchSINGfFNnKJ7Qy5s4AJcSYdZ
aWAJLO4gXWCXP34S+AcPLeIzOOBbjzTxP6ZwAVjvexBFOU629HXQ0Uic4OblYsiiLZQ6Ixn1LYhF
vna8/4eNUaeWzhnxNFwtz9v6PJZtM+yhUZA6sZ5/586JsXylEDb2ZxfQyaCjCBOYFALznGSa9Hus
rULezDw4rc+QepxFPaymhK046r92uSC1QGT8fGMy4Z89H7lPd36l7zWSl75QKKSNb3nyTXUB+BWf
caaz89ZhpSL6DEvxBbHTD30zK/M9RpQX89kJAJIJEGKrEzQAvlY1e/g/lphsNclFf8xZWNfGvp1x
8vXJgeFOdv4DXL9S1IRcPnGAR3sI/9eNqWceZ4O8ukMbT+QG55ZtRfJt3ftqD+YbUvbMvTrvglHJ
Hrc2PUT46+EqLlVWFInNjhfdCDYeR4Lv+1CjWmk4NcnpPwUTqGaIG32EIfzlNZxdaxK18hLFaiz6
0Nmligca6V6id5JALApjlcgkg7+F1aC3rp9jrGcAH8iuE6nrT4gSLkEKIzudFkNPSvDBLeA/wzZG
r12hyctAm0QK2Xgrl2RTpJZBQxgHHgqq4BQG01tH8JM8q9mBZG44RNPGVBSynB0X6GYLkv/xMucu
cybEjDnVUUY83KhfIhHkJlCmNARldM+c9W0qmrV44me+On+LjBKUAS6y5bI4YkH0VG6KKcQvaaZL
3wn4Q7eEz3eCMF1rB1zakmXTNLYGkhMSHSnBlNnB+mchXKFL279qJiQcqv/tFAHuw7Zv5UWXKpdA
V7IQQHyIklrUzf0zW0AiljR/FWnT3TKATsAwReMnzOUYqvcQYN71ULQK44yGSFc7kI0SjWnJO1qZ
viq5k/c8NDSL7aqFPbJrxwQwgDNh/F2wB16UnPL2zUjlSc2Yt7l0JA6r6cWq/6/d7Qw4p2Ccim8D
KK29o5o8/il4FAScEOv9EDU78v2H87cRn2aljt9Fe/rN80D8wlwjaiDJx9ZdOPB8Je534eXQBTwb
Ok8Q7Y0mmyBwQKGu14fthA+baktQAV0yFRjqq9KDp0O9W037PddebDiyxWcWEZ52fkf7sC7FP+fE
mSJVm8D4yZoohNCl0tf/9RSprCk+7zt0USSsDNaAejBLIA0AVT0t0YqzbL3fCKVHmHKqrnF7f8Hp
+OwK7RbrpD5UI0YVs1kZmlA7I+vgumfKNvHi5eVxWOL/Vg9JoBTBge/21L/rJlSRWHAijDHkYIW7
aSGzBuiaj1IQuwhfqM9CEP5VZ19GKFzWGa2DXnj2lPyOtsMhT9LJ8tSR5uqSKiphzXJqu+CSKrem
i0AB9z21B294pdxzr7xKMNWzrzWTn2HzjnpGAZM/hImR9wokx+QLdR5sRX6d3s7/amL+5V/S8V36
gKBhLh0FOXL0N+6+74k3eOmlgVxI/XLKq81X6KfA1pZkPbzz/zbz5OTkTKNFaJxGeJGC1GJR39FP
MYDDMsRTMf42H6kUlZbhYQrTwgFIo9xpODubxcZFlTv8VfpYWEnAcMC11JWFq7Y/d2BfG23PNZ0w
ibEQgO0BiTWXlVnj24Isjlav2QJbX2l8hmZwLlqgakKuk57vQ4WrwNmCQkko1IVXaSfls2nnVyDO
NdEimJQOnq5dbScjYf+GyWHdiNtokjKGzQ2CU7QSZDw2PopjMLR4+VoIiWNeCWBaflh1Ubc5HRkE
xYPWJPib4uuy3a1CyY7dv9qZHL83SDdu/y2Y67Jr9gFNYjgVJs9pnt7UNDXFn0fLj2X+vxmwDUHD
SFkMX/fI74ZITqqlMfzvvSbEnsRUD8wLzzULmkljuWMmRl3GRBKmWfvTGjXwVXzt7GUNEtz5Aubu
jEAaxYM5EqRwDmScguwx4f80MLCuJfDBohKntPgZVkLoTFjgFTiA9Oe674qvgbmYZjiuXEWAnNan
OMf4U4VSWVrsNr0ssvWpTj1yxwsfFjGPD+denFYgIYJHh4N/q1iB1wCTatzyduqZed5O0pnXq9BA
jpOlxyTYe6kQ/JJgXLbrTzZMqWkqKQJO+VnDb7aQjI+nv6ZE1r3NHwwIeDGcQNmlkz93R+c2/1fX
sK56ekQ6+hwJ8K6aHAGWFH+Ct7AL0vAFGFM6/8yINZhg4lnf/Ol/+yGB68pOSVce0Qf7yekPevSW
CJqHAUGk42IkQ7NAzNmfun8xoirA2+E31ZwnMJYKwZTI9qgXjk7wMu2kcMIuf/u9jjfpYgnRtxNT
pBeXRxHomf5ihGyttuvJSzGX3JwF2LTXmpu35ihGSD4jfUoG/vgxQiKy7YK7d297XKeKJJrP2/2P
E5oy0YigQdLU57d1VWy8GzsROltSkLw+eXsVUaZjZU4g6ZOvnW0eEUoEDXD6mLPWqwqag6LD9g2x
XTLQlpv4+zUczLAa5opfvqxgTScdE0qRzQIm7aCmpGMMrCnF5UhIKXf4GuXhM7AaAizieT5teOul
vqpnbw7ddHnzBff+/LAPIAOEHTfAtr/r0Ci4RnltGZx6cBXoTRHCddnh0gYyi20QfcV3yqTrzbXs
oyp7OLIQrdqQqlMiXNHBqp2s/YZDidpUozoYb9JUx+BMLtXycco/8LYFaPQuu8nx83lf1y4lz/ho
S3cc/nzwCkPrYyk+TraFtAL1BnLKvkS/feOQL8KcNkCWmM3AcotlZn69DCSPqappn0g8tnRvdgxT
2aaSSUW6UhNIU4PMGjbZREL3VYrB+8iJ17X1r1C6bYBSM1x4J2KqbGRCT3YdteCEVFnwZcVbJlWP
T4pg6C9xT2ejtaZzt2PGeG33WQNTUkU82fT6iqMHFY2icfeEjB0YT3gseQuGyJXKmoa3mqWWr6jx
95ep8yVosOZQk9XYabKKpho0UaTauHdC24xBrEw2sGvxXg6gOLWudmx6nYrvIOztcrPi+8R+dnii
D7fOFt4+W0756JcNMpeuxLnEnzv9kHEsxfcOEqkQOfU0YnR6JvMd/eo4dKP9r0qvzy3vsl352X3A
KPxFRMJDZc2HUaqtOlNjIembyOWhKjpgaQhpzEklWB6L9CP8pkPZUW+Ojdk15g78eztulNb2slOH
ucBarc8gbKr8F2Iy/QvVUaZDDC8ttgUUtRqJNziLaUgi2LAuu2LlIosNwesi0p2DdZnfUUnovsBY
JZU45eAyXW1P5H3umRtALojHia4FeOlEmeuDCmDnmoTPrc8GqfEUNfkrSfGFxtz+OXUs9ylVf7NE
CCi+/MdBiLAA9w6Hvb1HhHAv9cpJAKAXtb2dEomDOlH340GYmW+7oZ45vnbn4UZtttL97E76Q52r
nGL7plR12zfAu2dWxq09WlF5K03COS4UCLGONbDRNx+4OmILTjAk/+6Z2HXPd+oMPSS7rv6OSNEL
aubapcNAa4qYdnKNUXlymEh4k9TMKj35YyN4cZkesvd26vUjKBKYYpHaHwjoTbiExv8vJQ1OoReY
a/ITMIApG1IOGvNlZ0CNay+WNxyy75w3clsrWfYLDVeUej29o5gkZxq8MA8Eyj9hFfJRWAwSam5E
7AXzBHvYlyACBmdtNEwPwqMiki1MY4bcAFNfm3Atru+s931D2LUsM8APfZoj3eDui/85mqzF5YUK
8nF5oQkLPAQRDXfQygIAxgxzLzWrzp/kgCAWtGLKMf9V74Yeh7A81xvcE1RfYrIECl0Sdoeu+3Uy
WnWjVjyIEJJZLjza8+M0OgvPf4lvWBRrz/0W1OR1sFB3d9WzV/cq8Xq5jyd3YNABpVFeVtCRdvOS
FWBShF6TSJtOFJFwDJ4SbmnhdhjjrpfMz8+Gn8519I0PUNg3/HAcRMRIuHlhVpQRWfPfHVwLfJda
tIZr6IyEknt6tqvzTYfUK9bH2nT1rEXz0owJQBmzto0rdf/j4LV0NBpMq8tDxOspazLathG7kUfZ
6692W3o64E2+W4sm0u5fHwT7idrqDJni7qJwD95L/VD1ckyaaOqXt6uwWKzW8FRMwqijwHyxICwM
on9j7GqMrr7bTj0d2gzaAQzjnH4aFlF9vPebvXvL9v898Iyb7QiUP1kj5+WqNWNrW0IrRASqBSJj
tFTiPoISH+HtQHUmqpwJ4SEnIWoj2sABCe+HXlQJos2G3z6u3F7SJUhS4ET/LPLmPxKjk8jDdFtP
tEeuSlhC1L92bF3oIMHzCwne0iKJdgCk/ePZFDT2egPtn6w3gZh2jMhgfz6VBymUH5g2YDdkKBaN
0O7OC9VY2VIktD8+ceNQZU2idy7GlRzb4ZcaPw3ZT2vGDecT/YqaLSN9e2QbZ6iluhvv6nURWTLH
4nib709l9aONH3Q3YZ9/pO6q/18bf0LlYcETp2YcmBfeUPNLnAr7WNdhuakfy/HV7oZ1l5F6Jb9j
LPto6hfgCiXUlp9Z9FYUzXqqgbdXzBGyhvbKx5iTSrMjBhi+7VvHLB6s3eOeXTgg0JEAJmAB9Po4
aqtdiY4cnAmBmpeKBLzUut7BIWh7BXNNj+f9+62PAcuyKyWMfd2GBr8EfbLz0Y1nGAB0XmXldZBH
+lbd5drj8OX/afQFr34m3bC4gtqLqNomfmKrbyqjOj0yaqsfiqlptPHATWs6fEEc0KZgVbzoLASU
nPsxCI0yv39WaQtwxQv/E56cx7XEDbHvWr2QV2GAUke4gwPgf2YJGPxcx0BzBFD6t8S7+ZFyxymc
bELuUjEXhHcX3WaqEP+c69LGMJlNK2kaFHpj5/17XtykTGn3dMpbdHBRTyzQYm8qJ5qaggZtJVJ/
vxUszIQtE58eySvoAlu+iXfG8nJrj3tM3eyfmm0xGlaq9yQNHE06CSewJYPw/tg3uF5HWXTSKW59
yi9cEuw8fU4+Fpj+xblrC6KyNXxyMXUc5VdsYhIfw74mFUmYbCxeWV1mujT3Iz8E40OZ6uOqS0tS
RTGkuHJU1CkZhjfBAfAtDgoII7oj+LSADIinIXSza24klgGGciLfDz5H33hJtsWmLLGaVADAmbtW
cA2hcB4zqfdu6Uw8QwBxRh/ErO9hKypFo7tQnyjAPiwtrvPd0roP2pnSgIFw1Dh5/RTuwbSmC4rB
q6pwD5e/6a8K2/sjch9IVmy3rxyIDdF7VNcRalZhe6CcrbFqpSBDum5u7kRGZepufnZmFZsfpg2r
YwLZ5SR2oam1i/B5cZT39YLxbELhZU2c3CnZMwpXIHisRvWtfgNwhuESRClG9WY5t36B2dm6Q7/K
HjQArO2tQIqyTMTzcswCeGXSAaEcF+GJ1kKi8vyyrRbOhGS04l9s2zOXx6K0eSuNYRRGbhuZykUQ
0+M99HIy8Tgbl1j8SNPDxeQ/xcuDHbHZMxfBosr0yIG7hczg0PnzzPJTMNSD7xK8kIR+MrHJEjSN
8QDXg23IbJ/nUkXazN/cuOz8u9isiDNFoExZ0d95DEViOfnUbwWzsaaW+M2xy72eMw5qoVTSmmsK
MZ4oTr1wKRtk/UW6nLJuQRvSKFByvndwKemvyb8taRGjxtUat4U4LokhxliV+5fpFbPTiG+3YuPg
MDmlkwMYd/psNvFjEN5fOnZkRNpum/k2XT7yrD/lH3hmy4VetDpqx+xjhkmCHruokGDHL2O+IwVm
8WJSpWQvY4IuGj5ah+2O1u8Ron3lOaX5Nm/a9U/SqwcRbNEgPzv+GNQKToWzT8oyxaHnAV8TY0Ga
ShZC9g6Q6e6nXhAEpjJKEdxb6H6jPZSBCQDosE7dw1fJ3l4kfgpA5J110lWHtcgqq4S240k/jWeU
SCXpWtD8j8+vMZ1Z6bYhKDps4XTLTiFZe5t3LsEb5hlJB3k/V9ishZqZx2g6GLIUlORVmJyYfRBO
QQcwk59WnvY227YOxCm2YkkncpIozo1xTbSRa1NJ1bHehYeW17jxtcQ6R5Yf2qG6yS31pBrD1cwE
LKfNuKDcJAtXIAjBBzferFszYjAKk1ZuZJ5vqMMTO2i9f9cC+uAepk8AYZ+yobSIQxP4u14nM/Qx
wJnz0indHVgtOTBCCrqpbVME83dobjKzZ2NBst2ADTPqSEuqCxzhrgm7F3vx4fizIOITqtLzBYr/
xkdiceaLqXkC7tnadU4+vfh1tYamsW6Q5MeW4HLtGI/z0K9fsTF98HqRlh0FDFpRc/7LrxOOoXbs
/NmGOyS0IQKinfuGiSvdyTqGyJexnHnjyS5Lef0qmjdX+OhdRTqiM+Ln0Y8Gelem16++ga1nYzjM
vnX0CsDHJTUXkeXdIB/CbUfqefrWnENE5R1S4eqvh2lZYYcOXmaQsHs4Hy64B1WiMtT7rmDGi9Sy
5rVDzB+1Ak++fDAQm6JPhw/6S5bYQ4qOLHH3qY0uT/LKX8xh0oqUzy+PxO8Wmjx1U7lN6WgPtsvL
ebC9+kqD+NQZhyTRFEZYvIdwldNXpCCU4/llaP+eJGn+x5TH2EXNIm4TiSGAfcMLELqO85vHk/OL
MCwg6/f1MhpVSPBZ+CYqrQ/A7lgwW43hZuFrxZHUuKPREQfUJUSvuKBbhPi1aOuG04MWmp3jrsLQ
mJpgL7BoyE1lJoEP6lYtGRW+Vwbh23Ni33/ls439dZCl+e0ghGq4+KTGUmT70+u/tNMsYpPWrt+C
NriST6uOthKzyQxANAmQLEZ/zJEM5oFwg2E1iqptI+v8zodsXB9+pCvO0YAemwn9dg/eIR7+reNB
jJ7t5zSjbAr5ESp4WOJj0Q0YK08KFaer/8B25r8mynStiSr1h2OitPcDuCCMFNmEYNUbf01D7o3Y
cJvda6uZAfHh177hPPc04MumSWb9dyHIiBF+/4komk6NvuDcpBj9gKk/QK+8OwhWvUiC4lNvhF12
98zqdziYJOHwwZYpCgg7oqLbkPxGzOlqfcn7JFujifXHemhNSDtm+N58VtdneW2C09HNEdBrTgIJ
0pqlw04Jhwp6ymAZlo7RhPBjeQd6T4BjV0ELxRgljGc+q4q/gBqIxO2Y+dmCqtbkmc2u3Jvz7T1C
mtkD8ACA4XP+vsTJ/iNznmVrChkZULMZ22HW0YkrAyjCwGt+yT5l6fjGnR/VRilmwa9ldWHkog1E
R5EdTbf4ILGeoCF7SClpRYkOnHTfZJ+YuXA4v4RfIEHlnImz7BEUGha+tZWC37QanNMsEl1X2p+Y
pDe9yPj6IY7tg401KARDChYzALgHnEAG1ErGvZZut+uHKGa6c99rB/amcgXsWFzKF7CddnoCthE7
bVbsHs35r2mJgzPljdI0xTWVzOAKdV+tPjn+fxarAxlCxzTjuNNkyYuJAdjA87UbhT/IfyAwT0mS
SY3AFUhh7D0/uSNa6o3CK+unS1Z0Ms22Oh3zVY6wAh/JHBS1QbIrpYOxu++ZOzCtXWJT6FwVmFdJ
5X9TnU3Pdt2imVDckE77LpYAlgVxMdJGHB1HmoGr5letwE+kBDC/UzOJR0Wxu6a4OupgxFRfAk6X
4efqyqI8ON/BkO8rINrwUY9qbwqrGOTSUzHsojdp4Z7Bmp/fBVvR7uJDH73gaNh+2qan/2k+m2bs
zmavwV9q+rtOE99whDE3Gqx/Q98JgHNDc8VyEeQZv7aq1LreUXbep5xmEYY0NZ7crFoBuRJq2IHd
6X196gIOMIvrQc+WXKW5MkVaabz1SiGNmemsiebDs7EcEduo6/EYTpHKLujsW3dc6XwOoeeL65I8
uEd/1cwszteSwBWJixwJNb2fnrwqfH99UfklBzc6PX2nvKPPcGPhVTnN3kEft2Y4YZQOYwY37ML5
YDe+rrB96aT+DI5YF27WybcAbN5P5rtmMCEFc0o/p3JkPfvckuSUTfBztlRZvPoZxREQBKS8EveN
kO5wNJ/Go50h9HJio6Wqke5h6yKO0u5vP+nB429fA9RPwpY6c8GIuziYal4Ceb1834NlSitPaB6q
wGQ4qZ+npR34R/Ut0Ruh6i4++gMjaNqS1l2YuM6azfrQPfbfbObp61w7oGRYsmXKgfv15peHeS2E
6LKQHK+7ytjeVyTUgPe9qh6+BDzuJ58q1PgKcofbD8Ie8ewjVMg14siu1ALGeai/+nd/uqCiqD3N
J13gVYA0r69fyk2Gk4bEZE9bfD+zbA+cPGHIBGWscjZl12v42nafVBPop8hOMGY0Qadlm5ijjN56
lAppzmOtjGNHh3MmGmGDPdsBAbz4mflXSDCAY2Q5MFIwTeqgQr55k4aWQ0BfXB1M3QPr2W6eR1Rl
EQOl30ygJdzGZQIJCvLakuBrsWm7hmgmfFpb4UcjtUs/MpmZQIaoT3wxSnwgMUZPeO5q4qioKeul
k5g/9Z71ywBvqaO6U/6NjjLYFj5X58caKHmyfRNiy3hblXo5zZcJ/3ivNDDgxQ/5Ghd2m86t4LSa
Dzr2J7ScCcM9FgFq/Y4AgLmJ41g7oI4icBzh/vphlTpmBNzloVgCzAruh19leQCWijhW4PZdybXY
o+VKySnnCAzClgDApa9lAvNaa9/mYd8X1/xUX355+V2nqdtR1oamyVufZSjl4Zsz6Ujnv26qaEPE
+zIgJLM9dcy67mhOgD3npEsN79KQECL3V4whhcIX3Fuhy7AVEi466B1ZQqYFX+JGfl+v+PIeCM7W
3+ATXJJVDhl9nEQzh0J1CKqZTHjXwITHpAngGIDK4kwKhkluvwWEsW1NCMbmXv/bEqgO/Ix7msaG
BX4Mm6qiKBaqdBvCj7VG4uOHax6KhVIOwxNnLE0Rd6UmHyVqqRXJ40R6DspKpDw0TkKASaT1YQAq
l1NFycggB+xzvz+F79EqhbsgEssWbpiu2Oiy9AMCHX3nTqpk9JY9iqOa0c8Wy2GlwnU5hRM3j6zb
Tax5H7RZ7dzLvFgy0wSm3gGoRVksHXAz5bsWUhTDb53YSuCZhcH2UD/aF+SSThSQgiLcuH5cAssr
CuY0QPYuSNayr6Z57kCb/KxO9dk6FyBG8LDcjnTj1CczDEmzutHsRNmBs1gfdxjZYEJTfX/yCn7O
4RH6gv5KH9H90+q+4S/kL8/s+RPqmSQSwJUU3abBwuGaHRxC5vD3pfI0kcwn7ltISbGEAahVlrgc
JTxv9X5cMXe3gQOcOVtfZvoGw5SZe419L6+Vc1AT53KGUhY0UlM3OKHKlz8sot48D0oW0pvEVknd
fCvbtsno3+BQlrJ+WGDBRStjwz/M56tyq79KhG/bPRrkUO6sgoDl1zX2IhdYTwt55m7iK+CaIRcU
59pNCd4X0q3lnWNyoZ/XjfY1VuYeL5wjHKqh5nBjFXerPF8FF1PsH6v7pKYokIlMEPmCMRHbpGpt
FeBmVDgkThi9nDNE5RcsA7NB60OLmscEiGUQ9bnnUsXtDE5+ra6D2A5kizK98ai8g6pMr75eJQSd
qUAXMY6xaq6U2vsxKr5PyNErLYam4rd5g5Bc4gfmMhrMkSpn9vKTXKP2Kj2NMKj7jRrfT6fe19WM
3vPf4EFcsQW2d6ng0nBmR6dDH2qFLli8NeocPtde5S+bND/piwRjNjxy52+UseqynU7z0LD2DTeH
1TLQwn0j9pgqRYjnGX2pwACvPWWgIjnPjrUqCjtRnJe7lClEHV2BtxQQRU6Nd8/1uyTlHp8G3nwc
ugDfJZCH2MI8JP+c8C1qHmgN7gqUrkv66fgVGHFwZvDQSXYYnrneqvcHNh2K6alJKptZaMfOo/Ez
t7+rlbvUd9zI8+msfIxLdDwxQQu535sueRkll+s6zstBWfdfGO8wEVYjAAmd/0t/jDCdem37MCd2
g4Jr437Xgz0McEQOr0oWpQJf84ybPmzSNm8IgXQZNuckviIr2GHXMEhAXS9uegeMgQ4uVA/qbg11
hyfb1rncgOfoSSc+DMtc7ZWH//0eBRHAuOBkv+S9xdszfSk5hqpzLSCUOdp2TF6GmPAe7hmiC/qJ
P/d/dqm/CLjCbnZzUZQLnKs7dikBmzs14UkChT8jNX8C/1YiWCnD3GWQbN8TnAy4neo+TrmXt+IG
V696XzYCukcQC+6Viog95sMrXh00cKKPJtkdbUghygRQlspRrCp17zQXvj+J+D81w39hj0mQm6YB
GHd4Js5Qj9+yFxCRosJgiikZ1BHY7MzJNexGuYLwR24jRGrjGG0W6n253CJFY8BMd3RUmOG4uMA4
Q0yg1h2srYR3+Mx9KXaVFGM8xAVwbTXqivp4aPOWZ2xxug3nhmiDkWE4zO2V3K88LJpeB2DOF5+t
hP+hyt9rf9TYxMrQpokO11M/mt6IUCtX2hN7FHnj5umg7NMjs+LOiSfAipeN+H7PB5ARpejw6Vv/
+kTECi9CtiUTDTubHEH4NOyC/17SeKoXkt8YS27pCM+gfKg2qOYRdyQGAtgrC+nep0hYhwiNFXqR
t773VG/v49CLJ3dYvJ1nE80gEwclWAfGLxhd84NnberB17ZbWu4rv0U1l+Kjij5lt+f7yNZ5XPx1
NZZH+mP49+F5XuUBo9O/tuVYWo42pPsLBN7hbbFlZ0TjlSRQx6PspCBM+u2OO2DzquId5EFFDzW1
EcDAGBBkGrynAyF0Sg25jQZOGnkRj89/INsS/lvlidkFmfUsn6CyEXyGQgvJhIQri5hgE0GGmQSG
J+XMei/qHUtqGRe5meaHDWS3XzbG+9NSI3l0EnNdY/C7BSUDK5xpvNPGsOxhX/WaZHl5Ia2zhPcA
vYB2Iuts3NsRAa1iNUbH1iOqigcx5VV5/L7aPZc1O2AkZotKxijp1Bxo7pEiUxej2nsjfPOIwsYg
PNBKyh7oOz4Kn+o7njR6N2sCKBZy1cDNsHps//57bjtLeFXHjHMEKy8oityHGzgWfBbrs8lksxnp
TffYakqtNBkib3DOuM8omE6fjXx1LYvpSdCR01Qt6Tw9dIMmsDT8O4qzsV3PqCe3rCkwz5Ia0EKj
JP4SbJTeoz3ebQeaYWf8rGeLDNcbOH6MMksy8QuniHCm0Pa8DF1pcCSo0DY7HB+D0LR5qp9FjRJ+
aR+AJbiPWsCX6l22jX8dYkBgf24+Mxqr9NZP8oqjPtqc0iFJE17RBhH+Gs3A7Bjk6TsOESIHr606
aE08GdSMAfhDPLO9kisQUYNc7jaltbWy6i6LRlNAEijliyyGYh/MFeqRiNZbt3DBwe3tPgcu3Bjo
gLF3EPM4OFp+Ns7Pf5SyXK3pF9YFMhqiXHqXcAwwvkm2W5KysRdDpFntmWqpaI9u4AJ6/ZoNiWxx
yDmoyuDJ1KP1h85gM8JsCf6FJB/1sdpLerLwgQQX2IP4y6jFmP79vpjJGUrYOTB1Ldsh82e7Suj1
ty/WS0c94VPrVykhWH1CnRblx8dEdYHvCa7zD6S5GoXpSXZkVPXKmtITWR/xJhCKFGTJGsSL7Of2
9QoUuv61JNKRS4O1Js3dW+dWQM3skJ8baalOLUjNNV2Lrbvj2k07IqIkZUN/ptk55BJqbCPuRPmF
ihcAl929tcdf5F7k/a1I9FeUR0hdQe5CzJjXBfbp4cpjc49aZEWPfdV0OBqKCOp74HJ7gVj2MnHt
iRNJ/48t0jvd7TlPcuFA8xFmaKT+HVEIFNEQx75u8HLQsDhBDJ1W+wNCNoNyJbzNeb7mc//uSMEz
FoYazoqQItyaYX2bdOUmXtQdBgvKYgjWDHCTOKnHfwgN4Qma36+t+cx3Ik4C3o3pbXzdKbu8fcId
h+/b+xWGFAUoEBIhZOtjWTgnb0MZpxe625XGMokcDRYSwaC2v2FIC1f8nYJBYji4IGnfZB26V4XZ
q7mVg8z4+ueB2/e1VGmsHcWFhHST3l6ZE9woNXdj2JlNEcOpR4ePf7nbKEJ0xa1hSY+YvXwoQLPM
0yZSAx8GoVhzlzkV1wbBDu3tUHb/gVCJcgGUciTMLaizWAwhsEHm2Sf21KwnaSXLJ9NX/S9ruk5j
dTReKEE988n/8V8AGGXvTjL5OYGlwlpfcvA525o/o4Yn+sw4nW5nD9jKRj3u7kGACvRHZXn8A7/1
ozImRT/TGpEuki5tK4kLDlo1LNqICGzOiwpSc2WJU+XurJwmxeVjODVOZomvpYEQjcQahLoMhXEk
hGJWjFVQXkkEg3XeMd+KJtxmmItcPTrMk/4tgf18cIlTqkETXFf64VWtGOlM9pD9lbkAx978nHwr
uHqvzKGKLgNUzaPKN+fSkETzIMgeIAQqHHSL20QGWDEa3aLkBZvq9PoYvvpdqOtPvZTLLuflvB2q
5Xf8o7sqVteLfYknEMlLZWtPliYPz70YLPi4yLO1oSgUGzPPAn6jeFBoKnZ/TfSvi7yVduxhtPBH
wloXwKS8Unf9Iym3gDoN1wcLWMerA2/za7ydhpHw8ALHowbc0ZBI6OQaiCVJV18xBqU4ncUaRW8U
PY4vrpQgstOdUybnLBR2ZWzdL2JdhWJuat2QR5wA0vweB0SkPSyS1Q8Sugh1dvyH+lh8XVHFIlMu
E/OhyswitX7sG76i39H3X38JD3iAZ+6c3XQVIP6Yxd0sNDsToaYytsR/iShEE/0tkAccRY1IRDwV
lMlnOjp002MqoGV0IYD0hSVI9sxaQ8/RgZB/eYmdv9Pq3rH2DKVUe2XM3Wbhqyg+DV8OnRdoSRAa
XphtFA3yCaEwOLFnCDBslVoE/5fxdB7lWMAre5auHVqKzADi4t00DkxdJ0EEf/iUvIL4pf+lLKi+
bpdjLWr6eUfFQ4f5p3bqIXFRSyElMOuSlE0fcs2nFKUCDkVcpAhraEjoUtAHanxPIi13oiyXwdTa
tXz0+fTe9lgrWHAKltLHro6mN3jQpLxPf1REFtAXLdWEOZpi4AhpFJXM1UP3NGXqOEEHCZB0AGty
l9TpEKiKl/vPfdiuXgcaeKoPVqk2ZGwdfHMR+zCPpcNs5yPch4mF9bXwZITZuKCdQ08QnVJUeOUT
m8XQDRzemvXhtJp6wP3KMcyVkr4aK95XCIwqusQnPky6pQFpJr/ti2XFbdEKEXYbaog11WB/2/BP
8R1Z+DHEVnhmX51Ql75k6127RdNq+INcsjwtu0dxO83E5aXPhYPXS81aRT2o8x488JV0vNMd0nk7
jGDlpPI3Zc7JKZeScu62bvLSQvt0GhJVrDZqAeXn7Lq+1GmS7umvo5ZrXXlUSM/isLbJbwWr7nxe
Vu18x3KwVZN2QpgJOMEQpDhIyLE8GaMFOEBQTH9Fyvel9Ihs1w9Orojz15OLCJem9qyXpVCSMdsO
Y9FZVkc4ixcUE0KVk1FgSYuekHHlPAU0PLtxFJKI2khnaOGuJgc+ezgpWJ4oPPMRb6nJH82orPsy
XbReexfQsXLbXlxYa6gbO8IpV0pALwHvvAmOBSKlbrkAntC5QjLYxWX95b9wP5eYDRskKm0IULAM
HthgpmowgExKN1xgE35RNec83ObDlJPgkvWvEcBLza/bXZjq891BzItx43qBE5hQsIQ0/Msnz7Lt
NVqs3ycZNNbAhYFsoFY5qgrA+fDC0i4q+3Niry8F23uTEPd35oU1Yx97dq9mPsuXUihVV/WxD1SA
rFUVmC2uD1trGprN3bdNuqAD428Wzs8aqQzX+1G//ORnMo54/2g12+daIuTkt4Ed3OIlvjyV/CsX
o40qcVdny7JAQh15pT7bOtO1yk/mKUCPIQhr0efg+Y1+dXfq4ke+XJiVJk4GkAlx45rZvZDN0u1r
ML7UbTkSPtDpbH6fWUHF6Dm4sQf2symbRSaJ/RGys4fpiivJRexJXuDziePM4osyufiob7QoEdZR
CmNvPcy8Ni3arm86PwctAD7pEofhv/fC8F+lU3sFtMNvc6OJWJYUUs9OMm1GClE7F8PE/1MU+ta2
fN8YgarsZTCCPnGwmPrgkQcF4Y013kJmkd2D52DMMohARjttqyXStT++L3efy6mKIHb0JA+bDsbR
IMkcXwCPvqweLdpzWe33YXF+kP2xoJv9CJ9OYwpPKW55xXGa8D3aEVV7G9GAq118iv2Vytk6nBjL
g/DZEW2JnMVpUjwnwI+JH8GM5PnExmgvRV2DsVnUXTj6jcd/JeI5UVHLko1rCdm9H7nmD5QqGj96
FIzOt19LJpOijRzXPnPZ5ocwu9DTslUopdyawKg3v07nhYJowWkBkIrQNEYh+f/XDJR+rY3gFIim
qf/z0KpQVsWJxkKssfiDsLlAXS4IxA7TCBII78RD+cFgPQHpqxGVhjHjhGRpEcOQ5wu6V3q6jfm2
4auMVJN1p3DmyZ2JVCckDvBFq2XkR7WPlKcByfMbOUViJQo23vnVhMwiqVwXQVHsB+nWnlf/PXdZ
1YYDfJVoKGDu/rIkuaxKPBdDsUaq/F+t60+cZ3mQ+dQswESlsVkNkg9OW+8cActBq7PqOfuXBkxi
RYTe2oB0xkEcfn/uz7XMq0vIzD4WxGOZU+wJBq1ppbYj0/yPZJ5C8hpt1szRn/UFL8NPqbBrZYhn
v0ZqIhgAh6iyLPX87Gjnz/mmVuOGSXzuPHZ9GUXGDF8WvQrVgQNRHd/ZPZ4s3uLWPtJs7oJfDoDh
5YxpB+eA3gWwDS+tYG/SSj4zIeb4k/yAtjI1aoNL2sFBLOvVl2BvzYD1xd1yI5DcuAcSIyyVIwvC
A+9+0ZSu692S+rq6Wk/ZesAZgV2NYwQZjMOkxoUH1bh8LzTldut6ibplMHkRQIUwwGLfKjCfwyo6
0TG4H/0590NhOzJZC+3pgn02qa6l10DhymUbazvs+XA/iK7mssL6ZGYIjBrlfJj7ofN/CQqSjlYn
Fgw5eLuZrOM8pjJQ+zEjE06n0Wy6Uv8OKy49BBbU6SN2PYF+4hx1JjvG+urgRcHb+Xv9TrXAS/IP
ygp5dsz9E2lNf7kw59BAVAcrfzSfo3U6SjzrWNvuWpZCzp6f59CEvaxJJn3BeAGarylBE1g8O3ra
lSN7UPPwKHqUN0dC5v+zaI+ltrjiizByOIdbHA9rx9YWOvyrJU3Vm/AzEVJZNlosYrCbp9jwglX6
GQPsJERA76XTP1UGbITBmum6XbLq+jjQVl9lwa4ECNMfczdk07ScwNb50VhC1Ao0o0OGjDn/hz/P
0vub3nUpz0JOngc0HImXJo3z2L5X6UBUkjkbw+d7lB4T4zjXbYWiXCirSL4R0sKZ/er1ykPd69/2
JgtBYukpPRxqFC19tKSa7+ASwsLt8vj7DoH6Pbl0uM0Y1M3YEt6Iok0nOjjXx+99KkIYvhvapnh6
fhtE45GwJ0DAl4vGPQDy+fLdO21nzxIJjoeU3IRw+1U2LRF3kt3u7ejy7PFM1zOL28wlgPGgCWNk
ISuDhfHyOz0C8PO92lD94TjvG3EtR37RPJlbf1j/m+k3P+783692n2d/ziLWaeTgxM8a7QpcfiYg
2CNvhPEbPhcNXxzYlZGJEyrgEMyRB4PbIVwwD3GMrPyKFki8b26Ukzdz74ON5IIvH5M7A9mlBhXS
+WxokpWyVU57jJHbbsvOrZs2PP+KXhn4yNmtCve+RGn9F62Ip0mRLrRJ1RiRo4kyEG64+V12NJsp
tIRu/YLMr0bdfHAkE/0QS8Q6nM5ehrbm1sg3WJtDmX++gyDOYJBq5R7rYVolfeHU0vtlV1dnwcwa
A6sFcUv3NcD2VtA6ltRbfkDqHjCw8MxGbrSgbQSZTQqiDVvmboRuTrQlrF4WrwwOyzwFP94Dq4d9
seBvLD6atpNcWYtjmVIG2aRFYjeRHFaM/Wy8v/Nb6qJGY3cDtwJAhBEI9SXwldLmbVFXuY8sZdL0
kpmgeUQtoztA08tQ7GbQbLNzpUbkR339ii+KNaGwPR+tltBPX4JZMXQtdp7jXqfhM0uTTiH4zEO3
RVJCmFV4i0SCJvMmStn0Mv/FyLmWUorZQvN0iEyPyX3Jq+VAn6JbmsVaGMPLUsC03Wk7pVVU1RwK
qj9X1MyWlGPYigREg8po6UvCqLsUh7TpWe6Gv+z5yUzBpSbwbkJO/LK+NlmVqwpzMU/mHAAln/Nh
DYaCJ7miX0ORHrAS8/UI6ZMxiLQnUJgzlQeQ7il7OeHAd6Kw7wxB38HqOJKHpTmfWlIx3JCAp7YW
KydQsk5KjvXGLb7+U0AKXjQDLrM2Eop/dJ6HBOyYeNNvmAsKEVCr0HVWRDtKtD72eTGQdSVysF8F
uBTxGUc/o+AwQfIzX+2edaX4hxl5j7Fl1zRWibW3advzET9HPt+pG46HVQx12PpoMhsVeJ4Qp+Km
ZA3U0+UDTKkp94NojewkXhp5mVCtbfWRT4i6tD5UHnGNZ/g5rE0LHwcl88lAl2lowrvJ9pO/2c/y
bkC9QJnXruwMjL64XeZhSXs6iZBuuQBpx5YdHsj2KXFz5OmywUkhyUPDaASAaW89DuI1/d1oZhwm
fwCiiGf1sEVZR640+EpFnF6CgzP0x77KLzrIpkItulED6zfvNWGVaFYte/PWzX40Fdl8angf62UO
isv5y9LuMgASmAMbrtOdwXvuvJJVI7n9WNcXdMc/+xr3SURMwA9HxE1kdzmDYE1Cw4PBW/sQKbWi
DxhYT7YGzUtMmZ0w3YND+qJV60XRv638w87RqBIqugVGLWTmTGGVwcSCrxQJEg9WLuXlKNhqd3sr
M+aioCDYpZLLPZavpfEaaHBJCt+U7Gw6zbW/lfNvp1bgyvbegoZ3yZufI4ct77t0f+cdgis6aFxR
THOLsb53MpJGMvz6+1eRZLB4dgezVmsI4xaCyVpK3R5qkYYVfffgsoQlXYe/Rae8wuEf6oaqtGia
ZtVIN97wAdGUy/9TE+GZ/Mk/9liVvijJTvVlH0Sb1iJXCCFlSB0LNcBwV7qqFks2EFg6ToyBjKZm
ZfCJyFlkizotYCNtnG2NOopzUE/43fSqin1Cad5WFztW5GkGas7YJYig/nbpExwEOm6H6KmoNqDr
l1urHnRtY40oeYfui92k5iREfWplDaPXD4UsLa/Fcb1YNWSMQ46llicqi+lWGIACeb7cQOuxK5if
OCMuwEmX+3smlJQK8TB9/sTxCt0+vG2ebHD4/lqhXXyWjr9iQ3fE+oUViW1C0L/X9ZwX9yZV9a2T
GxQA0bmUmIQkPWe5Kn2yg8BR34exWqWKzXrh854wMxGQwmUEoQHa8wfkYBSAbD1u+xgHpLHoNprO
BqFB2yiOMtTAGv/KDJ3YYQCkHK5jcfg0vDSe/w4vaHceumL8EDHAuUBpt5rvvPz7QteXeN8dhDNM
w98j8NEsYU+2cmSkVarFeV2KqJIi/yUAHHiWzWTzJJqk7pZi2vavuG9S0irw2pzCVFpXrQjCpr5y
1J92vdErUAyulsniMT9/fUyiG27PbBAZaaL8rxEPZThTR81AGtjTuLLAYvtylBSod4ANr2EkMsFJ
DzvtT45sU6lXAuSQE174K2OUBIXLAxZXVOOhG42tNybCLGhCROXAfh4krTYTR9rZ7wx+DAOxhbAi
cvtN8aSGZ/I0rwN3KIEtARLSh5gUhPXiSkAkp7qHfT7TyGPN7p+wCbgk30iy7Mlucyp7n0gePZgz
XOzHyRMjxDT9tBgrJwiM/M+HKDNVunNqLJOwFvRGiZWhDUVUuRajhmzfHoBJYOKEvb5/gWnEF76k
FBcOduUvku8avmlhD+arUf4mUG9712CIOCn+uLm6E6bMYBtcJyJuiafseAnse6ptGY83CoU0nLMB
2ydo3B4LyPUeE2H6wM7W5OaWIj4tvQcVYzVKDX2+bGsVCiEdvFuUrosvF+lusy56BUlLui8AEaL2
A5RlRCmt/afbyy/uwmuXGiLrsWD1v0LwV+UtZ59FA9xPIbx5pa9tHODFMENGD2CJufnSYSBtnl2Q
MCTgjXqemOodg9Kq0O81W8rshiv+7H3XuxUhRbaNLWUf4tLjuWxI0ntuKhB0PzOniAJdRAVIoLjK
bVxlo+xyKDbei8BAZ+NPndXAq2KIHk+HaqcjzX3EcAwHGn143j6cnID2ODrIWw6U2SHDvOyvpInA
1R8daA1/iszmWHMvZ2GL4yqNtLf70Vd6XPf3yG3yHCLClzx6sxC5NnsZGOPdk89OJ9oi+AREK4pN
VwbTpVwWpkJM2AXpXBKj5J8g+zTVRkGAaNK+b3fopnuH2d0/0C+6PHnBSNoUEgh1D2iwfgl13cpu
r7Mm3NDLewNmQ0FvJ9KDg69eIYfgLhV9U2Bl5xcCcXIMTQ/2pZ9F/xkpUWVuMta+n375ljJdclfn
zTaBfeQxCjCBkvrMwl+I6YIzVW917xNs5EV29rduyqnH8D6nNX+sRCaV9rrAVl4tVBD+HX23ALE9
R6Y+ZWpka/aR7QcIShs8x4Z+kIo2R30N6FCca6G1EPzw8+W6eqUxbTWcBDxTfGJ26hTDbdRnKxHi
Y8ACjuwu2jPaZ2d0tGSLLhUG7s1R8fab/vxKCrGzgys+cikrDpyE06CADUQZ8riCtdFsYfd3LWC3
MfF9aHD3x4n0LZNG+6AT5qZoibSGaFu45kA7BwHOJi1wF7/iRka81IHuBszCrSy656VonwJFTk/g
AsvJHVpE4gY56Igp5faCXdVYRMb6VIeLHl6gV1vdZkQvySgOYdo7DHDYxVyUCFD+5Z0oXC6DA2u4
qDuiqBdAwZZfnVUTQTEMz6eSYtVwSjZhR26L3mPSx5k1Dewh0MHP8LzRhOG5qczli+j/jYIXuzA7
aLMut4gA7rq+4q0/Rir2yG/KXiS2iAlMbLq1RRC7FnuWN2nj4svH92WF4Iija7bjgDj3fU6nD28/
xvFkgDiG26U90VmI0RVSL5sR/XiCgdf9L/Ln++2rTj2uJVhXuIfOXklm7g4UZ5cVZcbOOUh8qQBS
QWfI4LKyqNhdiqxHmc4+QJksHBsdjjFLk4OvYkYpSnLDR3uIApl40wzJgbjMmZRs7TLtRRjlhCHe
+N+hzLiBn9ftCujQ7uHclVR0OWF7lUlTVhFYatFiw17xFLI3xmktw0JxZkyADwHomUdcFo4yo4n2
KQAylHuEHcxk8YfCZJumr8Sr6+RrB2753agbj/gvGZXL7O97EVJukHJEdntNisSHiGV8pvPtnik9
/wuLb+6F6tCQjYh0PBe4wPbIaMrxGljTwT4AEZ/5wFPy9+my0ZGVlTQTd8+W5CHLx970WBXnmBs1
yNRiYmt+bj86OdZRcR1bKaDBuat9Qm75jV3XpK8+CpV8LiqQUz2AHDokBkQ5OUVNU/HogrTvMr2s
/LxSE1df3pF6HwmMfy2Qeg7nNUz1/fhcTlwI1SgOZubkhFnHk99wb9qqXLjqY02qbuVyXOdAZVhL
p8nOAl4cJJlyMoQ5f9+E+nnS5HgOj9/z6wWQdzScFFRNJd8w05TeKVrnO48PiPSEEytQC7hSNeBU
pw3UKQLwCqySP0SPHLny/8VcalUeg3knNTsbBnVWeqb0bOxlvZqoJi1JfQuDTaF+W5yYgGAb6ix+
polWh6uypkqT69Evp1w9m4X/YdBSC2HuFKEx+sA1F0Fc7kAqbwYsxC6+jbKLW+CblAT+r1MtV16e
Rk2FYAEjLswRtT1qODU1GlvLvT49Ssyl17JnUJ85Z9aTRCq4eoIW/QP89HhWxNpZynR9qiy26KWQ
9iiRlZA9N3LVN3jG4167IfviZ7Lpzf7P9foUuLHhmBqEtRVYf5lRT2MBW119U7IqPwdVNp4V5gDG
MNX133AUd/7AoZ5ktlJb16uHXvHuurU0RMlB4EnR0f5AEZq8I7YeiOPHj1X87GnwXa5T5LcDn0Rt
xkuGcTe1qYIFVdnuHiQEHP2xxleG3XE5PpSnXWk4BSgG/xusCQJOEK7EczgjND5SrJpEN+DivQJR
9/HKfqUffP2QLFfHmj/XucBCVkfhrXTv2u2bu9UjgcMrva7zoNPLBNOszjhL8MEsfPzN7QoYUxR6
jWbW9P1uHcmbX6SB/54FFQmvqdyFLt5tB/BAY8UFG6F0JPla+1vm4BL/zTqLQs8zA/0Gr84vHtXB
tjyDllfI1HmeZOCikcXlLspn1ve6OcTo9SkzwVadWLROsiVPl7v5CfFq/eo+LOux9dgKyLptgQ0W
nfBWkw7Ym++Hu5/OhlBMedNooZLVP8Bi5CYaaKL1p9PtUuqke9K/t5+cspcBOUtIYMotFKtufC6q
NITPDIF18BjNeQXvec9tXmQgBtYW2z9KGiIpz3zTX3OXgxtRRk/83BI5oUpUcH3mGVNKRAjhn0yj
ET0mXwTH4WWKIvfCAFDEX2fOmh8c1TtJBmpuilYrhd79fOi1C3J+Hqnat229UBHN6kTiHvJCsO+Z
J6c0/nLffVT5kSx4N74YgiHsKB8rAm0FVSAjLmUwMx9a9Upy6utKWdWgBLso5aeHATycAr/KoL5o
r9YxeioBx440S+Yf/Py3+canrdQ5jyVF0RYekHbbezUiCPVMnYzTbbW0eQttOzSLMcOIVxWtIEnp
RWt7/hvlDvMlEmTYi0xzGbEJWeHZTd6zLZRPd9/+AucbyEQ/bPrCW0l6Qof+1QGpOf8De1iUYXl1
DqqoV0MmVgiW+jQuPdgOQOOCWQ9nUEEF0LLXtDw+f3fYtxE55Sjx1JyR7P1TQZeTsggRCp8vzHNn
IgNg0otiCCWWuVweb61pfXnjbR9DsfJJllsQQXAf8s5rj/OIZLGgUmBJtFly33mgffv3EyS6OCrz
hvv/aog8bWjzylC9EBxQb4OD1lqs1UBS5eIuEs7S0bubmKPFZaaIwAXhujyHTRtFg+RJERYtkQhE
IdQM1WjabSJwBjdOdfA5lEkmAnQKoxSJI6e/2/4tKZAvkP8epWF4NciwgTLoHWM146GVDjX9Jxox
y7MdeSTJEviZy9m5cyr2beWVzgeH4/qqQ1l39izMElveghF/VHo3WcXi6hcoCTTPIckYocYw+gjT
qQvO10olSHzvizakqIjTNXmIMbyU6lQKtS6e0XlAPOOQL1yxhWqprRMMaxdf8yPEZ12Gp+FQg+sV
wii/9hN8QM59j/XrXxmys0Xus5cG6QaS7zC6KRL2bSsyj5RcZTRBhOIuqT9+bgEDRD+4OTERtCkh
nRb/Qbz9Y5+7Xf3u3H+Jl+9Q5u3pUDEmQhsczihj9KUC7X5P8lV5gcQGykAG7u1k5u4E0aLVr9sR
AdCjRMginRLOgnT1MRV/EBpmsNr782p4/K6f8LUNineohqQBob2+warJXia/uo7aOZvNNhbLjAHA
kMp7QRjLAHGNBJR+H4LLETLdk0VIwdIseKxXxPJew0uzYQuwW1KHCeeRQv9fvbY8/19LOmvrYAWD
5Jy9ySXIDBdejpqFi51jO198sNEk6sNLgJx1tm3DQqbD4nbsC8tclu2ptBRj+996cZ02vFUu5ay+
CEIFdZ7bPUb6asCwZOvWuzVtiGHTNnFRVp9cTw+lAHJ0KsfC+2RBqzPQmty1hqPNxIyrOgt3dN2B
aB2FpebW6V8F5G6WchntT5Sdl2XY8poW7zzZ7jYDI5lfeqUZzMxRCK2oDCaZMenaYF/SsznZxXK5
xk3/HQpZ+vrW+O2Bej7f2fyHAnzz/o64OPrRlMh8C6zUY8SaxpN3cjeIEqq3TQzWQgSTBE1D7sDr
reF8HwdFZm+mRINifFEwdiTh+BoajFL5DQTNgk2QnyxesfT264TKK3LTXKLB3Gybi2FFVm+8KU6w
wkfDtZKJ5nADERvbUP/SM6h1WVntV10909rG+jXG1VwUacL02NAtElVDRdGsER8VjN4PTPVQqTKu
Bx0VlJcS/SOgZKsEX8dd4QeZ8xg2J7MLzcDsguiWQoM9lCxcAEizKIjtxKbAj0GXKdqG8o46Qafl
LpIuHvgw/6fMILkGcGcrRVroLgMbjrFJUyO/dP/IHIyAVGE2X77QszxW6Brnj1nBpNHrxHtPzWy/
UJx7bu6DSq8asHrDAXHAkRpbKPlCpxorY3JyUkRmpTY/Ijlr1AOY9rqNgRSZnoJFQnwXpfxLYYFk
Gzc2EvKnYtGRfnVe/78LScabZjKb8Qsh5RE9uFW5s7kssMAp0guc68czu+MooEXrngCLa7j4CzkZ
9c1aSBbIuYUPJAugtSi1upL/2XqCweVgdKiu8avCScrYzPRyNXowDLvw7n2skQQ8ibMOuTW9zWLn
1fy0rI6wZm0RdiwaVr0W7ChntWeILJeCNe53kPTHWL23VlJH8G6cxQYBMYZKwEpMR3Pdos7AspLW
jy+1tWXVrWZZs1UhLldMZnwaoC6B7174rXuxiGhjA6A0ZC7LX//q20mW4wTQns43tXd0yn8N5Lnn
3YyeCanDfiR/dIMGxB0Guv2gl0cSsXbUGSCRlytDP532K9zXstVUxTqMUPaonmjf+c2IDumDttt3
w7tC35DzDbl5wEcQxNNqwHByqATU0vF74tFw5jqh2XnnuktrBK/7dbRhoMTKt5I/xM2Zg5xRype5
W3coZwh2DtI6O33uNOg7oRPeO3aR1MSOhddiZM+VohKWA9BVqvxx0SGKOkMmNtHOKDhatQtP3LB3
rJK5RkhqcbKQvbBQGurr2fqbaBnRyCZKzMzkdsYCnMltP7iAOH7KkhXDhLj1YpL+NVhVSLt3yaqf
ME7F9dab9ispuqLzw9+nJfnQPWAReZ8PXn2SlK7fuPtu/Zh0Vho7ybmWHBwVhktNnq3auJobl3k6
YU1HqLI6k5L/bz5VfQqKkkVGEb5DCQlDQcWY8G7TCM+1cEQ0f5BkWZPLZLfdJ+HJfNCEwsTjr8fp
Oa43aqYW8smexoud5QLI4cGNVKZT607q91NlcE2/ZknZpm7pycEkK+byyQjoDmKd3tR+TwsVLpTm
ZYZggbe/LeNMYcHg5dfyMJQ96EXhsYMk7+LO7wUjzvFRG6tjIfkeU9bDg/s0j4q8EXzYlVUboyOP
E8M/nYxG6he2iu3PV/O8qKhKwcq9PrawOZYCd/D54b4bRBx2nsGxLjYvvUrK4/BEJ44w81gnyJWh
rgKHWIMu5zQvH5vPuGm/HPaIrS7bWFC4ID/3IJFuBjmYrQ96MvqUuWN8s5m0qraGg7Ky9s3/y855
KQNnn7l21lY/6nnJhexlYXxMZhsKMDt2Hqn6lcRnR5wEEyu/EICgn20eJpA9qF67oufIFTsVJRmU
mDTQZkkBNblogUurmafbTodAMJ7aWeh+BIANkSYdJsqmC6QB+UN0fvXjYJmePa7b4WlS647q1ay+
V7rPsdvffOpFxOLzwvkxl50/HsaDX3bLvFA8W0nIIp9YVTk7jMBiCPXumns6Yh9LAtCkDE4OzfmH
L6JMszfqKZGUGEndMd5/EVY8j272kUuTtyzMux4ye/MCT7o+xXpoLCafABdLPdCkHEOE9F6YcYXK
fVrI8W3RLNgeZHTqU3wxBQqLZXSllUkpcd4GzJSA+G3/fdIv86Mz4LNDg22K5Ow2h6pyFXyMpkAQ
8XaKB8VDqVIfaI5xIFdZ0Fpo+MOqrBsb8pPFjWDoRu1plfXAbMiANQm3OZYMcMsL1ZIRM8hPoK7u
Wp3DSZVIySDWdeUggJfTMgao9pmlDzK+3CvZcR3gP2S6fTUDdRRJVDoKC6QTbGSQnniCXDIa4mOW
z04MGtoKVdA/d8/Bn1Zi+m0O95KAB62UB1QdltNexAzMsev4ObuOIIg6QE5u7KNpyOKS46kuty0n
4o6L/vbmJi/M4NHQG7qrpLvu5o+HmvjgCECjF6Ec1P7GHcBIvWCYeRbexiOhmDYZJVnnRmPEYHyB
Fo+J5s4791bW/vJKwxPAo581P6iA9oko9qz7HH65J3ykZCkQLgbLuI8k3ONIc4/4+c+GVTDK+F6k
+r7X0g6HJnq4Iou6FTpAj+NU+sbo4/fy7pdPiLvKZfkLaXN4TN1ZC/f9wPJgx0l1b3yQH2NmuYuE
qmcNkjoIQs3buslBc3ho3DKPRRl9hxhfo5j3evury0tVk/4ZKf7MqymkpmVjGKMC6ZA1geo5KVu4
0coWZyjMkuBLHANk1EPgUSV++fwPoPAIcSM+FdJw+i4/icZfCLIG7mQYHKB//ruo+hMEtYrp7xhW
bjGtj9DrixaTWKgUSZVVtAdNslE03J9Y8wNY6GBp5AtNg4Ji537GLIE2x2/mvLHeH8pXNwinJfRw
hymxptJredZSUtpgst3XdGuFM6a0TZx5uCvLPoZrskickWUEpl+Wadmo3Vu8IgMEM5TEhwwhNI3i
Jn1BTCf+LEQmoV1VsQXpQGsJntCt4yMb905N6JAaH/hFPKOS9QaXQ8aZf+Ys/MPfUcp+M6PE7SUq
pznjgxPxInhF4him2Orx3FpV7odHySVoVfrcYogytgY+PqIsTKId/gyI62ZIJJ/aIKW1WbWQKTvQ
iFx4Nb7O9N9AFqMZ53dBhCPgQ+G03QaCdzczlNHIylz4i08L/ZKXGPqx11LpFQYTtNkn0/8OUqxU
222GM5w8Uo+oFy75XlXRD5IbT9aMeksabQfwCFJZEnLKJVqDMjrTgGGct7AE0uMeGHhKcgP1WBWD
usPV/LianS6eEC0utohH6DYeVNoACpiLKj9Eu8FrQUc8K5K8ytkBkoyPEGTijVs7vGGqriecKYFE
UQoQ+cwEIVWpC3PJditDZOzj0wfWg+ik9tE/bA/1YiJDOOAA1ZSCZn0+Vg0iOgiBXw/SL4CxWjdB
iRA7JaYkoVoJ8FQwsXkStCnoyjruJNCSOFgC5d//jkxl3XSgm6LVkF3oYNFGKt/UGrfTs60Wmguq
OGkMIDGS/KVkT8o6A/UI9yGl5Rps0uh9zNudOh7nGkWsVS2d7S3IQR0/+SUdNs8x46s9pCf81JHL
vGcQLM3oB/0I4wrd0DF7N4fA6lc+e0aVYVnnhqUkCx0DlVck1HCIidTmeKzEjiAvylMLLlSJkOTT
Q55WGniAptrSwH4mLnK7QBDPD/NJ9oW3DUHj000DTdqXIJwEqqq8pnkBGs/nmfuj5ZRw9xIb0BDV
cgs1AxWKimPo/CoQ+V9+yZuLeIo6z+vauky/Xdb73V+Qvn8R8vCFDkkDYHFF2lxCONwnY7gOkG6/
rREZKUmLdACPM3bRiaIdkrNRusR+C8C7qu8/tcxf93FGNkDH5RQaaFL3Zi8sdESRx5PYpt5oouGm
AuOxoarAxiQQ7pcGiZNoMq19hLGaaThWGyDPbjQl5vShFY7VpQ1w3imuuzeSW7Z3GmPLb8508nvB
/4bYwqLYft7F0RK2n0VlBLStjCrwc2sHXI1Zwql5DIKXqf70MxlHB+nnMfhlUFeK3xa48N6KsbaO
8K1VC7IFxleymXlxBOHU/ivDqS6/xgGL6yqoFXbl/Wv98waH+ikE0E/YCmQ85AdjR0M0mRkMRSjr
3W4Vprv2+bXigQLzkeD0mIyZ/luTzscmoKu5izJiU9inKXvbLavuf4Vpt3GVz1/cYtS3EzqDOqXn
mUfwHaFOhKLHNouYWwH4dN7fVF1MG7CwYMBYt/K4Bxzxy3+hn7IWMnL77x8F0ynz39LCm0cWP77v
NGlWrE/+uGy5tOzepasVjB8aNEfJ0aQKrzM5fVrBdY0G6WrXfAx2qxwvPVAAjXdMa8+OLZuRnNKN
ZTHI67xhcDXXHfLYNXJKm9TU1E37UA7nusDwpwO/1b3ui4JpOwbUBiu2OnUbfXEl5ln3iIZY3W3t
pm/FoFbTVwutKvIgRjl36tK8AQuLMVKwXhdhuSPWZCwJ2LjSd6wZZb+FVpC7KcsS5gXhvW57KcXJ
NdVz+AcMl3Q/yFcXRnpmaTIhrYChixOaRw486+e4+MkZ1CxY5Q4ZkhaDfosVP8by7hRXdm9019NM
dkS4nallPJpBu2PziykONR2bF5ncb+4HTLFQCqIPmedECbFBL53c7TFUi6sn5JXK60S52CJuJenY
EzFvRGiAoSNoUCtGF/fGd8qD+Ww0OgQ+Gv+dH6M34i6eNxRDWVVVttwmuSSeVAGR46ZNymzcFCn2
aw1YQZB6clq0kkgk+T+h410tG1wSHvg2PTswJiov45RBYMkZ8OmiTOSUItoVhH7veOUSNZ4mFCkV
pcVygNXgV4TMMKhJHRUTR9xBpkSvwNhLD/gxbSKpIxsoQt12F3HxVbg0ljHTQaZvW8LwmI+l+CDm
xdMqH+UWG9sV7HLJXQJcYxS0qqH1tY7VbF8zrqwh7ozmmiu7jRnOuCPZKAorFXtO27AyxgK8KJeJ
oDbL93wQc456cWQc6WzcCD9uw9JNZqdrJbT/P/qISEkZFfvk/0tIMq2aw3tIvQ7LosOIJzPchF9a
qKDxOr+ZAm3cSJTsnJUVbe89qqGNJxAqL+cmKUOKJpiU9WoZsJUpZITNq0TW+AOK7r0A9fCOlaeR
B2pOqeaQkwK3OsTOwK6MpD+v3w4NdX0X+4SzQUjmNQOf8swncty4f1SnrCNKtGucWQEG9psk5EaR
uT7UB6RFEKdnXxRjqrEQJelucJQa/4hKbj3XDN6jhKojwJC1SE35f2p5ekpnlCWHkxD8Aw56+cra
U4ut5A7dSCHDYWCg6roGzgEefQKyq8zP26tgQ9VQhn9a0L5UIcvlhr84RuLv1Gs7t2vdzE66V5Rt
v7ewPh9ZtRCBt5tWEgkD4aWLSyGC6h7dOoQPJLsrWgrUna2bSc459Slhk2bj9Uv2ny6wVQQ0Jbz5
sp72/aYYyOJomPxk5o0GTGtwR5CG99U03r9c+uqkubXksLPtCY6hVQInRPi5Q3YvqZo4xs5gU54I
AcjfhUkSIrMMeCZVP6XD01IQDCiZn/zOfUyDy8jp3DPiSHPbA8r19C8taL3Eg3qUYQX73qKPlJHU
L2zEclmL/R4MoXOosMOx7SdXR9trRtVatrwBjm8InvPhvbG9mG0IZyqMGOr2Lm7mTZIC3iVZvjUl
0rQIAm6tP5OHmDmQTzrNdY5PFqFGXYwpHHF96qPhxruSHIQFALP/eeC2WNERd3oT1oei/fOmNjDS
UBJQha70ZFYsE/6PwicHNcKa5p2pc+HPFo+jKvflkKtyolUpQSJfZnUNLjSgL0yK3ea3x6k1/Gp4
BLDoVuKuXs8Q32wW6JQxGi1Hpj//UoTz1EYnVioHJIvHhWpZfj/JdCp5JsYRt2Jly9ch1KrWliJG
cffUeYvW7vgIPb3I4rPWFSKAdK51bRqccQuirnZzEV6jP3cvEkMgWUSP87Mz7MPmiIwxRKijuef7
6oItlDV0CGorD9mQKNApTslqBrbgZX/2Yma9//u0LVgzZkFbQRESOQbWqlKGXYlDj34jnjqPJTu0
pbIifWoQWjaWFlqnfBUTIP8pdd28iYNscDqu9qwvfPZhQaP3XaoSjK+AVNYG0yakgs+84R3r4twi
Ydir/Wy4+2lu+wURa1YRySKLa8BPuLZHvMF9XT9ILrJMF9rDLfMhuPxCaRiKLXMQ5Sz5Ceb6OFc7
jI0jz4RI+Axs5K/U0eIuOTLRfQEfVJll/zIanEwQVQqCRoV6e1AbqEqUVJ+I7XDZSsIae5Yyaa9z
Lr3cK4BB6cL/iV0FAyAIrxzVVarACPFMD7K9m6rwtpjaqB2M9VQ3TxPlbDyBRP/y5bb5NtpJE2Ei
zDY3fg6SNjHuGFG7bfXSiZ4Fkbrg6GcI50yibGEGn06IH5+rJVzNNKMCRfa920JA5/WLOnfXft1t
z/kmnscvhca8bxUkuUp75cPwLQTbsVdv8mxpPU199o3FukHoW9M4Mpmi+5fRtI4VLjMBawBkVFov
D5MdDS874prsHTuJwSA6aC22HgIKTKg0U8H5beI73F4rPAbDGs4PmfX80HLmraFYx0lLd3Vfh+Pq
Oc3uwj2N6mE6If0WxzwfDDAI5P50zLXBEucKVNf0NjAPspqhJYF7NEyJmkE3VTvvS2ooRhApM4t+
A/+iTf7nDQXO0PD0PXyTP50wmPOGmWG09bOLjjLDCi1Jvtl/Ls2tTv4R5KWia3VhKZvULcOYmZCR
Wt95P8GeslNHD/sXYO4Ayfc1c4pgC0FCq27nLdigjNfBFzofga/O+yL+pjsHQx/Ieo6QHrWWaJ0S
S55L5WAX7KM1jjqlAZI/zQrBqID3GiYh/yyBgyd5+t1yXlS0pCUhDCwWoA5jaaswI/q0fb+HxB9v
KFKlL0t05cgfbf3hTpTIyx5itT0EYz7bkXavCv0d4ZzR2TKDPMCV/oc+8PvV3qrHAGFRmB3Qsb8Q
FOZFKDHXBuLdhPlf6XC1S66f1JE9GBNvNOFr6poh910AKCjpJeym5KlyJ/JR9PZUSn67qU86HYgx
ViFDFYRyci/TSKC9fYIBNU7/OCKwAbuIA1d0RKctMl4QtwRPu1nJ1nQbjsLskxK33guqkKpnXD2g
IbNzbjBWtMI1sNJvDreYDi2PFH7ESEEDLHWjLZtUbE0Jo+2J5mGrBkyDN3Oor46QbTm1MRACAtTp
namBjWHMOhrjOcRxK4cK2NoroFwaq23fFqApyoKW02s0HHR9OMqD6GuF0R53n0AVgctARDy//OPy
Dq/yomyQG7L0yNkeI3bCdzgBO4kgY9BIpiDiuC9uC4tX3KDOCSTe1RjFy71TqeB68r33OjLEjcDy
Q/8quxdf+OD778/MsFHTGZwIYeXYUXPgURCLn6XgNE+QY2JF3XfcAW5M6mjXREIds98hsYjRdAf8
kg9iGGIAy8OvJWcPfxT9AwspIyu3An2QY54n2ZLGrnNJuXMB38ib6XUZjPJ4Wy29+olMAYmr1Z42
jSEmj4uMlfZ75MdW86JdxeiAWT4lmTV1JvFRbEeEW6HXVv7hppDYwzAD217vcxPcGUGzJ51AZIlr
CATbTrVTSCzKgrUFGLiwdU5KBbnLi1gcbNZgqpRzK79IQ1xsHQEB9MOUdktKAimZW3IA7teFEiTi
CZpoNBiOyjTV+xL24YgkokMh2j6Dd0xPUYzOCRJDVqQY4tNQ8gWJW9ztWTiW5X9x+9RGuCq/2Znf
SSZmfIIsgaqZHvpyKTZ66w7frfm9P7hAEPCRYjNG/77o3cyNhJgGZGsSfdsd3wh9EO2abfRAZ00a
U6SQYEoV3euMGF5p/cpIpZusO8DMdqTVgKvRX0BNt5ft801EX5fyA0lcQvn4tZEi3jBvQEl876Ac
+n6Ot9+lkhlQb0XONGN0j0h4hnC/UvBLE648y0UxVXNpIFyauOfnKocAOzRRda3hmVGSelqWjo3Q
iAffRed++2NCt08Azw+yP8t4RVS2tkHMSq4OTX2uHkxkN7B6now7X1TcbcDiGN/A9DPxko5ZMU2a
40WgKSAC4rBzPfyRL0FBepAKgD14aeb6T1WVLOrow3GhZBn2cm6Zao0xQQopmhpK51PakppWDYso
0VkmAVgJ1imGHp25+ALp3WIBg0EB9dVU/8yoyeQXQZwUC5cXUy+YQOktPsqePqWsgeMA1pWFQ79Z
L9BLhhA0hir7Eqmd7dilCq5CRuERgxSlCBDcpK66fZJgj2l1rMED6SBwG4zAI3z2jCuKZAn42+NL
9kxtUD6CPzuqKHxnVjhqAbOdcmquhReyPTnBmAz20zjJb9gVWVJsEFnJ7+JG3nH+9mEGWjlrndPQ
hSbAAYnoePqUy6B+n450bYmzJZSvpZsmpwMqhIERMcIgzhhzRjWCb2Mh63ZnQn1oEUUIKQ3SZKdU
rnBk7CAZkN0656VSmUh6+nTFOVdeBJsaGHRX8eBjmBZoVTJYfrCqganGKSfQMP+dj1guQ85+iw1t
QFEFOEQLwtXHZUy+MUNQEBNEEElbndPTejI8ImWwER9jCnLuwfePsu4gvcdgJK6/6IWt88ztdScU
ZFEJbugDI8EVqXcHtePmfAa6zRgn9Qo3PNR6tjdlymFU2LHP7mvPxZeyksV/IvJyhrbQxyvn0Q5i
a2ISzY7zpIJPdUOI/1FSexOrU+MsbIDMSmGcd1hDPpBsLHKjxTti2RYbU8VOETLYczMLPAqa/WcU
TdVEcuvoR+It+jgf4qO10gZz2xiWJ/t0R1QLQz8EteKuy/yVDxHUFlYNZzSIiFRo/VQzSNqHXSWV
CdUjicsYL17klM7+dyb1vJX4L6USlV6aUIXb68EyxC0cJRAxABAMTXtq20MSAXATDebKVCB+D9pD
FahKi94RkWgqaDnmLDaVFaVVbjSNxd6n0a/kn5U6K2zy6MpHH7/Zs92QtRHajMB3zVz+1vf8df26
1mjQDHTbVTRPvg5c5AEFU1GdEf4lSDp/2mm93RDHQsnikfAJI3V7VwF/+hW7CwS6gSHQHDC+dQjT
KQstTk0ewzC0YK2zvWc3kcqX6lLGEs+ND8rMOpZR+yhZ9/CxkJVjdpXLYh72/Lobra8id80POrZx
9ahEKdapjMBT99mx7qr7P00pZQqzJsSoN7AKDqxWNhRZ8JsLnJL+36pixDd9dd46VJnXd/45EsgA
oHRoVQBN1gslJdN6sZwe+yOWPbiXaJXMxkjsXg/vh7ibP3WUjBmWMPy1SG8rn/E9OdqfHpDEfmcL
lsa8AQC6Xst/DNRtrtHDvnV2znaYGYU1FBeEN6ILyvpz185jyCdhVg+DT50aOINIH+sNRjg2qgxg
END/KjY6IkVgKL7FT2pBDf3xe/kwLwqMVTJtawC5l8eyaV2dAKDqOpeOBgyspS8qo5TLHkvL9Muv
0hSA0kWlJLo/C/YWquNxCmL40ZcJssfKTzmKgkfY6tPhkgDxQAWTyJksoSz4LbIA+2awN2fwNRic
M+QtaJquqhvQ3d6/OhSBAASmspP6/2vwhdipKWGhPnZ8QrOZKsVvahE+ZAPcp8bJ1wonXyOa3b8y
2UkQwHDLk1w9b3SmUPU01XYZl7h6BK7vwbGFSjJe8Ng3CsCRODQCM8zjYg6ThO7Usb9cRP2mF0SH
rX0nCBuxgmi9uKa6eWoPc0Jon40YqHtQAo089Sf8NPvFd1e7jUqPHPUpOHJ1RVTejS+1QNUdgARQ
4FbVSXxG7Gu+ItAgig8IMfIHeu0szahYs2l9t+wgibhOdBXCttGBRMfpQJN/Xv0PoiNW722jrY5J
5nOBjnHI6UdWGjVBXC4Wu92EbU3lOp2yjSK5FFdLlDygeY5gXXxGFN4uvQmjUJJhS5msJcHWUYZe
XdFi+KkT8/2Ragv3VIJQPMdzf+DVOIOo5kwV5BlXlcOhNQ0RplfAp3KAEUX9NF96YWz8PIk5JSGW
HxA1ARjGCINGTuq/cUFGzBA0UIgUFNbmbiNyvPwu+dc1j5x5cDhrCPBCh2wPUSxNXC9YX35UqmlG
yv0i5MFraFU5fV6iH6TbSrrAe/8GHZDLvu5HfH/EvUILiy9aXdDoQtxueufk6mdX8oI687omVHq8
+bLDZx8JjMOHH5Xd68G/NV+zMPYQxnVhhf6ovGDEgqoj16onDetkO/VVDOPp7899MERyqbgaMFDE
2rt4KkgE6Ypl/Ky0n8IA19f3/IJ1VVdZObpTH6aNHcFODQdokc3MrBq7OHUAkE0L9Wii0+tJSttG
USj6ay7zYDYyf5ElQc+R2m7r93rk5OxlNQ7d5mxuPIbvulX5hsh/ik0Eky1J+6NzAfhNM5SHMIV5
Yl/0XoQpy8WwtL5Mwi19GV/WYPTY7cEPIkJgoLXTXn8gtDEt/6nJLUk18YQTHqT8WuvEfC+6vRnX
Iyd2ZQxtg2zq7Ykw+tYhlLktSNWb1YkoG3Or/0cVAOOl2mTCPaACz5xlZ15G4mQbcfTA8c6kZZlx
JKhzv98Pd5OPss925JNZTl0CGiUE3bgU+IjG7pNpNZsadouWTRCX6r4oeA3PD4N6iQ+DMQqMR1NP
zElOvBen9/G4jK5NNf/tPvkMqVkR/ZMskCp5gpZKS2p2FhQ818GOYGYLHyewEa3vYiKqHZ21ogbw
XVP5NFm+n87d+TC+bIScATJMad72UM8gZ6Pl8jYza12/E9KyWggotTpTh1VZHL8aZ7+X213+nd6C
DV58AkcJ2DMijElH1TjxiXA+wY2C7PUUOJ21wFHRMkkJlRhpidutgI1XjfNDxVSgo6m98JWJPyYY
x+tYzTClWeAPoi+i/xv04EDJr0AzGRxWNqKF9a2aKq0bPnHoac7BPXl2zO8vridzMrX1qGMWKUaR
qdygF8jzUGhY3JfUgaK3K0EiEx23TmsnOiyfme0zDyuRFQPnaUL7KYM/aDJgYTeODHLA+oSX5kMo
GN7nB/cWeuNUqkDsNiIUpHy8Y0k41f/X8ZGwrUrZ/L7l6y/hKfdg/zZnu+rBdEeLfNZxQC0T41dV
q+Q05oW/Rp9nmbvlL8ry2n3Lb5Rv1SoRK03e11wkjrzYjfq30WBE5I/DDo1D0mHFZrYjH4KfxwMo
Kg6m5giBmns98hlEbr+HyECCguMkL6Jq/s00Xe9ow6Qzy57PAt3Otgq6RhM41Ho0a27Q1OsBbgvr
7cPNHLETgkgtkMPjVAvyH3DAuqW+LF/LX/KZq97rTHBB0AnV3gf7bkFU0M8lVE22lU9+tPHjsUPl
M0/vHkNaggh9LvV7B25wqyhtySXU+A5Bmhoh06rF6R6v/sdKfKaaXis5te9WmDLihTNsKp8FF1FF
gkdpJ4Fzk8H9uWqLWOAGG39M8vWyvyKCUkectQmoW74WmEAIdBCa+oPHxri4yqQHfU/JDoQfdInA
zmvdvSgWL8Kneyqf0rkyODrYgoiKN9I97oE5AUPtJexSAVhHA/er8RKQAeWBEeX+HrNPFoQYW9Cp
LMmHtfN00CXrSzxXJ1pz+vdkuizTqHSKTzh4XQb38pAIDJmbwx+hMTxfQ55vI8TunII5MY7XnvIe
OEIo2QIu/HnchUCpMcrHSkLfp3wp/9rwnWMUSoWeG7snOVBzn821UATtICyIiZWRiNHfyHPC2c2y
e8GpKuP99NP3DhwgMzNIQ9IfdveimsaxgncPfxvV1RaeReLFEilPZPDBua7R/bTgXEl7NxXxDcNb
vrzNqt/pVJOpe5vWyWzt3s3e2hXsTh9v+rbwhuvgrGtFWfvtoiFpNDSpfL3KP/Pz3z5qCkzZ5QHD
fz3/UqTG98kAq7MmlmuYwIQGHNIHEaFBF+unAvWjlIqTQ2biMD2CT/HKCb4sENBCtdnZA0PvjsVw
xi1NuDGnSpXuubWIh24nd+QIw9xOOkeNZYfYmaxwMKC3MQXVDgW6j6uoc2hgmVFhANfZVRLfUVbr
82RoS4AWGLBz8gOlnHoKREoHL1iaA9srfcEpxYta/EnQk489jUFc2VgQqDTwI9SjO69JtfsmSyHI
llaaBmNQ/QsquBX8xhqLLqaCLzo8zA00g73Q/lbGNHL3jkSVFugkyzWfMcm8E85n+q01t0v9HSBW
xLSQt6mssZ2MBpgpePzpndcQuF61QzimkgRvfOZ74MOsvcQ+iG6cW+/WkzfaUGI5uAkWrzGkU4lt
b5s20hy7PO7r7kLxfEgzVCMfR4Pb/kaCObY7wwWOyXmRX9Lj9IfWl1klR1lCC/s+EN2UURBGAqKq
ZxRIj4+2pl5kF8TR/F1JjuRm9Fvt6U1wsezb+BpQ5MMdihAqOFwBfobKIBXnmSGK6DAVwWSsTI9q
u8u3vgQF5BZrGoGvWn3QXptvQrkmX4iC7RoRO393rvjUWZyPUqHIjaBApOWg1j53+h5jjOZyWL5R
uaYlyogn/fkCKGR+6I+/Rx8di1aCQfFrQzqb40RTqEkDzKOaUrleGLF82JvHEO3kgdjyBbBRkS2a
PAOrwjF0aYoGmRy+5LI2BhnaUskKGtYpaqkB8MvYTFk7uTAwkmJpTTI69jq2w4oNAtdvFe8zZzOh
Q2qXsVyHrdlB+p38Sf4HaHl++ZtmMB+7YwIlJ80iKcjaHhG4bhKRWv2/3fkGD3v0/z32w5RSw6Os
Kz8kBcvj+vutWFBNUzXQjwrMglLhPg328wQs3QVr/A1abGPwSRGSKUf9KEd+WIe8hIv48xKSRA2n
tZsSDQyNfDgMJ1hdnRNj6pxz3GWFV2ydjdNQqkS7TDCpSt2QC+BDq5/u0u97OnLY4iAxCompzOGy
shaP/F/7peNMgwwTwVSOzyr9S6Qboa2yWfiqCHp6xrU9n7WIqHKS0cw/NyUCBTDlKqWsRX3sPKcx
Qul+yu6sqfHAjW8Plw/ZyzKRp0+Wc9XDRzEBfHtJPsRBQuF66MI8l6QZtnN5ypLaXuBqKJ52mYN/
IfAfKlC+xqylHVab9Q8Cqm4rbcLZ3Q3pe/ZvedIgvaeQqeU8xqfKyFEx6k0mDSrfM39iqdPziO0+
qKBHXlN7w78q7/NxJOWYEiQZIyE9oq+CYQb09oXhvjhHfA1rdiLHGECUEFd+33nDpkUB1sGLq+p5
L076eFf1pafpNFhzrVyj5wpQOy5oycXvKqgrjWO+a/eWoMye2TJazSXvxEZ/Qq1A4Q39vHYzuPWp
N6PvSe9lG5LGY/fyF5d6gAp9XK8yElFnnPjLmlhsbLxG3NeddRgIcBosjlUFQyT66baJwyQN6LPi
17+lhij5wzxaQoYxH8urxvg7bkTnJLOqbtT4QvNZaWf7lxTtPem/4Dn9FQs1xSOlLfV13nJmtpQY
5lXkeut8A1xyj+iMhP/gov+BeQL4TZSe1tHarP0gN1S/iO6Ne97J/dYkrmB7A8zcYXSApEHbdT48
3MvkZnnqjmhGIskaWv1gokcb6HSNwuQKizS11vZHkDJf2WEOK3G+DwiTlVVp+sDQUEusdrJP2bTp
fGoQLiHCLAbsqBH5Wps7WUETbd+6qmhB2OWQnhxzTXiiXdccfVyteDn6Uo8j2lT/RlUUD5aCpLa9
1Th8ZRaFu/MR636uLGHkN39dE684vJw+0BJUdZoev2lbT0/Y7dMwIbyep3tIeENZAKogQ8FWZ6yu
h1lKfjzuF0+3mKE+RC6eR4TAgRITF8/9r0b3sYwoBNLpmKyA76YAUN41QBY7e8grK/wco+STtBLZ
Mm78+qyt7L4BNK9k/xw5ojhtfbpdyohuDLGNkm4+qhaYVlyP8eGqA16t9EAdmjczPzc3rA4pDxrr
vdALaBwaLOoAmyR3rLaJmuHuZI5Y2aGWahp1Gxwu2zCuBgIDWvnAPdVwEcPagyWTXA/Bo1iV4O3C
m/Au1iu6jnvMx7OHHS69D9Gip5vJMHNSx+Ge9Ps+qSDWLY7fdfIVOs64mG3pgFyS97LP3quxXkhX
GbPdmS1xoqa2tQlEQK6KofR1BiuZQnVBX1ItZ3cXERqskN+8DhSpPhZSheL4l+R1JKLU5OlFfP+L
lVScHH7/zWhahM2gL0h78TL8/KzAPn0RpFMvdwK847B3UAehKmgtFR5vqH//lKM6sciNVCKbRmqw
ToUJY+VgE+yBV+wu3KoZqEs8QxpsulGSGBUTW4V8AjstyvE52w3GpaIydBfae1opVUZl1shBvnIh
wnQY7ThAlmq4OyhiXT94Pwbzx3wow1pCE+0uh6ol5imC8/n3X1q6LoAtS6O0NkTzECcgOTvB9bV4
1Vxc4nlHkUS9S9nr1lZyF4wFxP/qTTYLEDRRWm9p/pQNuhHsMzWPR0t9TTKC5sTWTChhNz+Z8qQj
fCguGMTkGESw8ebQSNf19zZbonhiRntNN/kqM2fpBRcp6J/ppiRKsq06eFB5gHtystCC5uA7pCKh
4gHACG3uZru1QQz3hFu3mS53RCRjdiqLui+PbSjT9ZIhOfHeMyEnBShPyZflZ6SjmFzszEdg1B1p
zE5z5wycew5Y0QcTH81T/CLhXmNBYs25MUgoztNhX0p7hK4tRP8JRH+wWj6A7nJacLDKI5nSqce2
EIU/nd9uLMog74hayrjRK7FMtpavD9NpKqln6kEhAbZBwaCvYEgEXpEuIiJ921KFnofZpl0noujG
nD/vvzsAaMwaVue68fIK6jhWwwn6+/9CjGY6oZNkCPK8J389c11tCuHXjR1WhpnEHffmeNSvADcz
VUQAaCk6iVXbEjTqI2+0s/FP7S5tLcfofhaWUSCqwAbWDmN6G5EsLJjjnbNuKxsj596FVuNmlJWV
Q6bsjvHY1whsakR2fCf2IfTCSlRR0VgbaLk3H86dhv9ajrlsm1TB4X/9egAp7Cytp3EJ4KFMhn58
sdKr0d4VEeIGfGvEMUb0kJyNsTwQeWZpEVuZOj+ty98DWlD4Uyzr6jo2mcg55VXTtkA3c8gb6bFQ
0QU7ftbZCVUv9pNLupGVl+cYFdWYlkL6h1SDd7xDvgjmOmIV2inKDwv44lcFJ9YW++rAulSVk54D
d3l9kJX0Zv6GYKX9DfOg6oVYQWEZoRbje+a8hkPd76Nw0qLAI0J4Ln45IQ+faVJfH/38d4F5uzOV
gyyvd6NjVmxfz/klw7sVzKpx6LsYnvfazL6FbdJqLg7n1mkeakYUOLqA4C/aUAeCD96wxnkADlKH
uq0QfnugTJ7B/Dre99uQsV6ZRlac0RworwmzJmaB+xg2nUcKZnDbbGK9p7zYoaR/mQfx32MgHPNS
vyzRanPEEis6N8h0DC+WkZv6I1ojhpqe7q0cTO5qYkcNoy7So9TWSmUFEh5XI2h+9GskG1Xqittd
Rk7JhQ4iv4gee6QmCylf46XbxB1Z6IQ4fmVEWj+mnnbnYKpSD0gQdT3AA92QNOrZjnEneJpuONkx
6o6P6X0KBudrxmwi7VQjQZmrvg84xHkyedfn8l0CckQ+EqQMyixZ0T0gi2OMHGkhAjrFsZoO6TWH
/hJR4N8LZXGky/MH/2CMi/A8ra3Wu27l8fWqAjsOaGLt/jQugpjKmGVAHazvwBQlJ/CqrBrtmpTP
8GgTasbIWum7QoykVpiibMcM8zs72U8AoA4tZCLWQpN67BTZCKW3+lxckDsuXIHkxfHN2qv8qfks
3DUFvRBkJQ72utJlEDCsA3xfwYEcx5Ui02bwzG20FPmvqF0Q1E2G5fUdyWICK+GHqFo7pXjFp6fK
ctuR21T0f1VGKrefMlryVvVF9Q8If5jjuHDLoLdpzQRTToydOBZemy0DpHByvWcFlcF2XK9tM1++
6l8DHoZoA90+uJSTklgBtAMlPGrlhZWzNeApDdpyaCocyZqEYK/a51qOqgOK7HOgBK/w9A2aO8Pj
06TAk3BhpW2hLqql/oDCR//W5tNxTzZzzen7/Oe70gjtx2TruxmD4BsjhlJ0N1OAr83M4oPV4Pys
Hyq+iN5KdGUm2wSFDLujTsuuyurPEiDhxiIeLzgsZakEXXk2jJpgljPbhtlKiKOLTst8dU0EA0Ty
lqP+2qe7VdDFrmRSRZht15UHHxCJEFki2t3PDdUhSVq/f8/cS0CTWJk+WgLS3BvgRKX6WNBBX2fy
YBveNEgfmAskaPaH/1DF3py7A5XyCGhMcfQRlEWLIjA6w1uOLz/wriN5wnYBes/gNc96DJvW4eA+
RpKNug+QoBkDqm7jo/abEitA25jbFIegWdIkQUp09Vhr87DoIdEMhPt9JAi+WlyOUWSBZ3DbEFRY
GAJxhLGYCpz+Y+Lt3sni4UjKpD1uQ3sCg75RJ4nRORi7+i6V3o12oMnSiEP2kjvFkgt1sZaPaiIQ
y3i0KO80RF35QpE3rWrCuPST/4aZN3CnSUEtzz55+/cCJQIh7aANmxWgUnuLqUc5VxvuZ3cScxhV
jqxGjRRTMYyeid8cDE9rnp2Axq5h5tm+QNMvEhMJoP4E7KrZcbD9EbUcPs4+0Ubj+aS2fekzWTGz
XmILEiqm0VG9knUu6VI6hyI2QQbkifUicwd1BpsijtA6w9xwQHNJ5rNdDwHGJWl0p7FPeZyzpg8V
Nqn9CuDY/9b+MJo61q9orR1X02h+igSggOGrzOnAvweJ8kh1QuT8I1otZAfpwc+GWqrEoysbFNSQ
gdSuvhyc/uYu0TL0KtMCbeYstoqd16fRYdxdKfOP13/1Zo843osZq4PB+3wsXtbofWkyvxcnrvJ9
l2PoiMLuBg5G7csrg9AyNzNRlwSM7fqV5MJSHSQRlGyDFAtZodlDBtN2TlmtyA6/TazsZjDjHOFm
QAf8iMgJ9SHKGVJvewO4b0SaOw/M6GfiN8LPx6M9gxKNifJ6GSs9pbjA/0z3Ma3kbo2c8GPdp3V+
g1B5xbDEiRiRDHD2oyFaDQJbn8GFBPYTNC1Aa1yQqHKP4wg2BUzpW8V+2VJ5vSD/v3XOpSql/NMC
rwoXeEiC5CzFYb6BUIjk7hRUEqVQ/f5VNudIboT0SjCkm1FyUoJtRQehUFqfnNg0VDHrOIujv7Wv
vF2LyzYLU2LYveZXMomGGu0fVR2eUXoMjNoMNd3hHw7+oiMkUvfsV+OWsa6rBClEIEw/m2+MIlLG
wamTYuoqBaRhvblgGNTK7wtZ+484pZLqEvl+UEVHuRbuwjCJKIOJerufj3TyGQ4eKoi/NbakYo6b
HdBqexWwBOkPD0dcdWd0RyQxkzide7eRNi6s0d22FePBdooQQBa/gPITLPq6SPg/ywrO+EiOFMRI
ApJ+kUvLPpnMTpdibN+oYpTueGC7zKuz2Nvs6kIMMaDHSy1HcYvd/vYi/1hVKks2ztZBNLMOALxj
UOT6DA1voxSo+sKJ5B7fz3fFZR4db544prAmUnIyuHCynd1wnJ+Io8jwQcXfrdFxpumLQiFgRUyd
GNazCulR8tzuTUabZUVQRy7GMOcDAOWhfjD21cO8xcHEbc9iABNzx2UaDDLOuoF1kia7ehmEU3Jo
CdMTe7LVJE+CoHZY9XWJSZChvLuy0sqUBwCIx768BO+hvYzOzvbUJe5XYAbSP9tR0L9LlLUkwAQR
XJtl6ECPx7SnNOlLC1nVGEH+UkV06G0gbBCQI0/XwisgFtbLJA7MoxG7myEphwzSGKPgLiXlqbVp
E3BmTMSJ164A5aH12u/AWaV+mqur7NAATXs5NEx7no8BAkr7sEHDqZoxfbBzp2Eexg6CowOmW8p8
Bj2wJDEAVW6IDIasuN2BqajXWBuk9Rr2Sc1PT48Il0sHgnZ7m2hx7KXXNSv/gY/5C7QVekhyUf41
iE7d4+JT6uzK1SpGaV/1Pzh7rI8a591IrqZbgM+0NIt3cDnYSJyQAxC5tXZ9l+b/TSsk+cZ+gLej
5olfuCtURBjr3ekB7laF4OSSmXKg2/aenOjxxlxdRub4x+QTe78aBQCPnK11diGQpL3UpJ+3luYo
7DbQ/LTVXOxM+6WtSWTU9yekPKslJ/0wnHyezg49ZeEZkQf0naQdFk+9Worn5tAdkCQU+O25I94V
xa3TsHPaHy9G2YPO0OGW/ICNw3QbNZOG2vd5Y/nv9bA3BzejLLi1AO2x/poX4fBAiFgL9SaHEErs
TkvyL7JUExP4kBPecuAlTXEVClfoe4lrV5cp6Uowg7L6D13r9BIZoXf+gE/IYrqkXzwZw/uC6k7q
ksaR990PH/beFzIdkxwtdMVYuYcAC4Y+2DQC+LElLXHNFfPAVsW5S43YPSRQWaSMUIBd2mvNlPoV
ennB6PJk/My8rQPaQ6Kg/401v1Hjz7Z1hmxctpUa+ryEThpiTBol8nK32Lqvf2geBUyehN7DlnFX
pF/D8eo4Id+x6lEE1KqRpwdyehJUB2mJAmdMOdYbcrBsGBL9Nn5UshJPC3ckjueqDiqWVJoYj62j
yaqtiR8m2duJFnPr6XWASqoaZ4wMlL8l5GXO+H5aIsgBaBp2fa2GYXASIaiU3eZVT9A+mJ2RQeDd
uvc5IzNLC2ViCU2rfwteVnQ/eYlJ1Dwt6S5qhXEw01xSBHUp2dhZVe2BsECk3VFrMOnHkSbL2S8Q
TdhEW6/VAn80XAou6fh57rDe4WT0LXo7DT1PdMyf+1aojiCQAzIKIVOUh1jHbqh9je8AHmK4zBd1
r86YNbRdnwgIZ2W3YlGzHQSGI0ClxeL0yyANy4bMNpEEWmDI/e2adIA+zmKScyr/UrXzRMnI9+lK
Vk3UOrSbNZQsrnowvmLUwtBp+9tPKeYDIK7pg92oz+cGvcV/9iVPm8l8EIXbZyf8UWRysUnwAUl2
nuR8l1t+NhRlEKGh34PelYNmO1YMCdF22k/5MEU4EAlFUVdQbO+MX7MGtg19XRcyNqSA4CVu2G2u
uH+nwZ58spV04ZbD6+jOsSuErRY+jJK+n2TwOmmsubc23Qu/bWcrK+KY+IZSlHct8NmO559Cx4YV
Yr3yxg8ol98Y5Cb53ELHD6HjoQ4nB4rSZzIyVSNZBVOYBhCM1PyED4sbBkg5Z0huNmYdvNLiXWVp
fPp1Ws8+429WC3eLPF9uevsM0ftP4U0CtoYTZsYo2h+HyOcWOD5rQHm7fYZOrZAseMIX1Kj92k5o
ugvdIr8QEskSxmxAj6kEvMZDX6Igb+DQmXfajQ16xk6nkkhDBgciEeo2j/DvxqriM8QU+KAa0+wx
0SS/xZtEC0qtZAuMf+CJUddkgEYE4X58lAAy6xDt6O5YDUuzd61+Ck4LrUr+r1jd0hZy3iYi/5Tq
oQiDzUq8mOqTUV5I2bSvXmdW1Ew78sR4VpUT5Srv4DClf2yiEEPeL/LBsH+04Ro4sDy5zPIeMYIA
4Y6wBSUlriyktsQbQimFRq4flGSrbFOFquRB5S63WxKI4zqunyUgohdFqr8cHF2fMTrHq75LSm/z
t9GT2D+JiVnmRugxwr6nHkJtkyP+cV/tR1Hg8KLHL5+pJokxEe8fFytPyRRQtEojggv8YyMKuEHb
gQAt3n8B5kkSmchSuorxVjmLrdPWdWWkHNv3snFt0liY4uD0QE7kfsLmCfIMN86VmkxSUQgtlS51
ETMmzyjhZmDOMLh1cVWd4udzaMQMiOrbsWe4k9mqbHgf4K7lMUPLrWTIKIRDL9d+keD09NsBIh5t
5adoSETqgb5JRfzT6ZAYH3dVyH0RreowGMP3CZ9d/s/LOumznVtMY/SEf5jdU2WHwv8Hc7CVCJsO
3OgFoobtkt3pZKg6pd3tEa2fiJGhnu8E/dX18DwV2FF2XRSqiWcTJyEAUazAbU6+kH0uyT3iFfpN
4cXhZw7HQNfkQtxWohcAxUHbj9np0W4QymGO4V8VVZV8oA12J4Xp+CdxAkimHpdHVr8z++09POfB
yFWxNvWCjIYjc7Wpi3W4lpHH0R9Ce125/wn13QDtbN7rgs6Uln2otU4j3xVDkBLR3tQsAzSpHNSS
dxIuo2sM6WyGHm2xrv35bsIpvQLY/p/T8pWbhtMujoM4LtEb1Yhh1nc/GF6HhIKf5R3/vtLGHhm5
GHN1iaQJPvPukjL/Bcm5CKfd5X5V1QKxipBRyY1TAYINWbE0G8yItd2ZDk1nbBS1/LjY0SMtwwfp
6Sw4xWOtyE4SxtT1dhho3gVXcEHRiehXJorZm7Xrp8vIW6TjkPplWZJRNEQ4Kre3KuBvKUKUSy8W
m4oEv5aN24O+gk1YawKxpCkrHP20XsoXdS3EkkcHcnD6Q15N9ZeMqz6QolEFiJZnrJ8VV9TfKBRB
HZpgCjmy7XaoIHKS4zZBbyOl06rxGXVOvPnX261/wldR+4+tguByDkqySl+lqA4bNv3TwnTHXWRp
SEq13/qOCqejryXLRL2IyxyEr4qNKY0KwsaJGTzhdnbu8HCCWIYpeGogTeVI3O+7QciPvKK7vnE/
pbH0UCFklCEPSVSHWhIGMApwAvi3OBFuRAWBb/HhmVkth49mhEM4jnKYyeKQ2gfUU3iS0EKrxQkR
fUke+WBEbz8RF8G61ZRme6yDJu/sH0LqUb++LUjK4IdlXvHUjk34QqFpYiT/8yF6l4OsEFMJEEFL
iX4pAynJER/Ko/B3PDXItmPWkrWgkYBtnhMhsPmDVHXMZ5sZsQhfCe8vya+qaeDGKzjX1cIV4H0f
9T/Syb39CkTzq8c2rnx7mMUf+g0AHP22fcU2hVCz44UAEzjJelui8KpicE3SjGZAKVwD7UhnneCU
II9pwH4zHgfb41Z1y9155AhaQWqftO8OHBxcNs6ToF1Mht1kmooYwOqGlsNWUhU/Jk1zeSJwg0ct
xwWs2BDelPlwO8xT0RSurbHOuBw8eqcd1YFzVnR4ihi2BaIYigFfsQFSkbxAx/RW8vpCrKGuRNN1
Qx1eHlrwf0Sq0yb2/rZICxed+Va3yODMS28LbhSwJ8+zBwzDBMPiQX1wDhUMsw2waBS56j/CpOJn
USdL7LpV/wIvFnbDrOh9URA88PpXU7zD3vqKX0uSBNQsv9XOZSPis6/xDV5oKjlFak6cOefVnKIx
kKj4btnfcg3QYlPKMsVLT9YpF1a6xYdsnzWu+ZUjsLIFISnnxsoyAVW3bgMy3WbgbBbz+igo7iAd
8pn61rREjwomxMJS05Akoi/1Tq8AX2sBDyX+eBuGpsZuDIveKWKYtIrDJoO8r84x6hBuAFZ3euCl
e+az3FCozdWPUvLqEgD8EHG0IQ7Zx7sZ7gAf8KmILfwqYRQBXAt7YAnIjWgpT/Yvz3qKhRLaNGlY
LUhiIpaz2lvm55JmXrx9RYDIcpRaFad6bohjTvneqTgdUYRgpFGNaHXhTaG8Mu3VAzawhiP+IRox
pgr3klwxbf0EKp4n/dTZnP0aWd27H4EkAkIb8dbBgdUOXU5z23r9XQDGJPQnLGe6I/wOFiabXFuC
oXAXpcYWdu83ZPiIEZE0X6epQypAJCFHcrnf4verInMag75RUbiG5u5enKp4cXUNryWFhVPtJXyw
ltJCMCSFp2pNOm5TtYXwF3i7EP5T/PfN/gv7k8FDvC2LQwKkNpr67B8QB2PHD2ZbNrBW+gagl2/Z
wclHzovxo3QaeP7UCpIJQ4DCAP8F2K8hPT+o6oyxVnhGW5VHGkp2nK87XDfYytJS8gOlnFEIe+ln
9aUHqZ+mCc1irZyPNTE/sVMGtmyBgLR960I95knHtsxweEQ5B03BD15HzyyGmRVdKvNHU4qpvUsQ
08FGmNX82nV9lOADO6POlbf/rIzvReyaso4APqZUWLws7n8HUhOohqQsh5p1IZg9cFxPz8POS58O
9b2uB1DRRUpXxfGOymW4j0P8aYhEMEFLS2rO0RxvJ6vvfpN7SzRo8pyoOCxfaBfTa6vzcohnngzE
ExTOtLUqI6qPU6zFSW0I+Lx11LSRH6CHs6M1eOTfS5VDJAIL3LrwnEWdou8ErnzYeDzkqqWfh8Vp
WQRl9LqLnjnnFu8ONmpje/Gn58CqRrYlgvKYhIQk3T8Qx+Qt+evPmM1cbGM5eReIwmdvfx28rJFe
K2sVFMYiIi44K/hbot4UtmxVA93dSQOPg6fqNHIlJC68gCsa9ywUkn+oXysptiBIz9RxyCk76szv
iEaPkROzdDwWyAQpsMipkK7DH/fl76GPGTcPwIQVPPL8XuwwtsC0apGoieJQ2DDVEiYL6Xqa4lL4
Xe9YPBMnDdFgR8iTRkpwe/+zsBpxvVe8WQbsWWQDY6U4jNzssUP8tr50lbmgJb4H4btASKsKPh1v
bWCtpMgPv50tD/E+TqkvJuqZb7lGNi2n9kBs+JpeK/p4UKkWE+jKajyp72rGYWO6wBsbVMYsGIBJ
mkFafISstbP+uGt/VeqZ51uWkweyGtMNIGJ9hqdyNw8fqrd9h2i2sNfW2+ILoLlyiMwR+glN8xoI
M1wPv+2zN4Gfz6SGxXI7VKVLxYlENIbRS2CQ/WFf1JfkidB0wQRO+i0wpW2GVs8TLpZSMC/dd3qZ
9bbFSTFKOcYV0j/7v2llCN1fmTes7EFOprPqRYMId9Uj61FNelF1wzUUj7aVvNg04CUndWjaggVz
EqkclyFpCprF0G/bzGd52W81JubUlsuXtuBieF5vGQNDdXY4SgLt+iRCBDYuI0KASf0YcaJPpb88
iczE9j8fCWuiP8eTUUaYBHKvdwK/WjfV9L0YYvLJg0D/52lK97h8MTVCQPKFAqAVM4MuaICu4CT5
zyzBfUUxa1egjhtXdmpY8dJWw1xoN8jY57ZOv63LgOl2CqUs66lb8oZEsrIiTK2oURfq33cCJOaF
NUMYVQK6EYp+gq7DjM3SnE02iNzFI9+1NxSS/tON9ZTMyUajrjf72kRoxC/A81e80ZAM1h2E35Cq
m/gwTrETPhsy76ylbKxnxI6SqEInKVuaz5GnNrpABgSOEUoohxBOF04nv2GFwG47+9Q9KeTnQHMb
ViBr0cL6sOtAuLGf8KIiAY//rSTGMpMUIjQ60jAYjAc2XTUihYw3ARydE7hSdn6VQAPweiT79qO1
JvIs2Wx56440KM8yqx+LU7fDfselCE0RSksJga6l4EmUNHqUhZ8Vnh8iPr1Z2X84DybPyC+HPIe4
GWVJeSfC6V9vcqYB9lW9B5MOK3CpG9CV/w6nOYjAQeLZp/+lS1X9MjsYjmwXbi1Qly9Ta70sB3Ir
4JopEfC7k7ZzFm1Dz5+obkuNZ+W7viRwau3lYm/jLooWnbXxXAnLMq2KIOiE9qdZ9WMf+mMjriYv
f3AqgZfrqpU19UNy0/NULM942sKLNykryEYVaNdmNgqEennTuos512cqR0tEpoC9PGEni0kyQSbX
1bOkN59mZb6UO90wNYG1Wo8pmnZLURyKFwEQ1qBP04R7+y0vlWm6R3+DPF/aGSKy/ul62pYBhAud
XV4XHp7N51nOn2DGlZQ/Y+xZy2lr3QS6UxG6xLJT/bsbTmm9OLY2KrfFsOxn9v3jXRQ1u+0lyIi8
eCMWUCRrGm+r7o/IyfJ4iFcR4Tee1AvLbwd04jC9Ngq3Js3NehruXuGnRs+qEkfgKTwvB2ULBQyN
l6zLRdzI++ET6nliDSBiFxyVuVTdzkjh0OOHPq9Y7z++Hr2t5lSTuGDa7GZ/EcaWlEqr2K6Gi/km
aNXMIYDG0tO4ocljXrrTE7Kotl3z/vaQ9iEafFqXXGT8rapAa2cu5wBxNTJWmmhjht7MW77LcB79
aqm8e5C6TZ/LeaqKTDGy+Y/io+rckCbbq4UsZ1JU/ex5yer61+AY7sduU1yhWxfAB3Gi17Rk24xO
98QTU+Sil6XnddhqYLZcpPGoP/z/T+f6vBIEZ9DtmmULPOubWij064xqIar3mSHW23U1GBUGG4ZO
eyluLw8fKcSgkdPcntw/CJnvWkAMWRR0k2TeEKvJu1r/96Ie0TWTcybHFnYlI385FQfjPaRfFgiQ
O6emeM8ogyl3nx3YnFsxnsmXI28+yjvyuiGgUKNiluL20kLwHtgY7KUih+mnlou95Hiq+0Hw34uK
4pkC+0rCttD+ao/C7w04XrzOy7Bqt+WxYp8T9doedmWrxpZwkJli7SX5DozvdR7ffsdIIxm/Kx4S
PZ5KxegR7C+c+SU5U5ox0hHm8t2sCdez5oiXiXcvED6NJhVm6JaBQ7Jn8IO4yZZWJErpJuC9NjjH
FAxPVKujyZoveSJAW+CDi6dD4W7qatwxaRm9diqz7bCRSfZPlcnudegcigOO6jAQWOggO/pM2/ZK
qSiok6qVnDeFVbT25uKvtqdM/mxgozqbkC6Ot6srABHB+HUvjkWBEPmp+kntGSfU8x0O3OQR065g
aX8Xbpvv8fqGq5f7udA5Y1RthAPdia31tqksll1Of4JphSqG8VItCIq+rs5peShnoBkjICB+AtNM
Y1dW3Dv4sLXKQvYAn2oephf/q5IGybTS7pp3kQFoELHaoIk5lUiOneKSWGX6Oc7kkXf4CHv4txct
zfdS3SOfAosWnpqqs2tc0px8Wn2eMbxviq+5oR5R1TOGZ8e+EG7FxTd3LU7mncB4LhQcrqzQXJ40
E1H9r0elf5YBrT1tUQsfUWqHfo/p1eaFu2/3PTktmw/2+SyAGxNCJAHKTPIMwVyJI8N0FOg4VvH+
qLlAbxmBjTQe853k24DWq/RqRTkvLFs7I+o+cL3kqM7Bu2mVAzQIDBuFRZsG9dDXCVkliXC5gnND
Mvsi5w7YjAIy95JC4i9FVB/fej6zL8cPSWqR4ZmSt97lU7fIQkkI8+O171Ilw2u+ZFCM9whdIXMb
xIzDQ4sPEEkcMNdsTuHNXDdMzFJvykcB4fxTft3DIwkhB6XMPFae6QGZDXIxYfJzsEpk2OR/7G97
/KECLLljJBhuwCHuqwNR6YIiyWQkhshqpPT+4/NeaJ4bQJPbEgP0nF+jQbTC5Tw3sSvP8XTI9Ktx
gdvZqOvfS8rplPuEW5FqV/FQ8b6u4Kp+rG8rOqWvI6ZQLxQMT/ttQXj6NYjWbHdRMGcjNJh9+NFC
/8Y0+rQPv4fUnHgaP5Dw+/czY3Qc6AmNN/K+J2pVWgEoVMKTANXZjK9p4rqaGAsd/U64Yi9OfpMn
ObNbQnkdFyrJXlAyAv9PlyCxEg6hSudnZ4v7XWRa9QDjcD0kOT9x2f1OEd24g9JtVARftVUSG16j
HkmSVUbpv6goeANxhGFe4VB3uJELXf1/zjZ2UGvS9AFEOMvFIGhCJzP5/zRFONJRlMFoEWHSfPwc
w02dXZnOJNfNv2RMcy0t3Tb3RkKAQyQ78aqhEae8dEelKLK7xYDGIeY6fm/waUJEqN1BxnTacVRI
usHsv9KTs8bkvyEP1ENGyziCBghZJ82XO3wfjhyTMF4S0MtqZNwGkB6EZD+mLlzXHqxbV8eN3Qqf
Hgcv+Wgb0Bi4k52TaP9jOY5JGZqtRrHPpVRNXj6KHEg60mERwhqfiMxtUQR3pTeAThJvfHrZrAzx
DRIcE2e+jq1xeChfgX6uWKP80FsN8KvppP6AMhCyFgTFQJfuS/EX9N46TVjh/MuWl005HD1/vOIi
p8exIFAL2rZ4ezDj04zuR8iTOQPH9BtEXT/S7YWeFz2S+qHZDcXvC7Fnjh4yA9SGn7aCVb5A3dm1
+CAXwdHZAQ/ZtGfFvlpnJaCjlEizC4dlV9aCHrBqcMb8W+nCKf6Dr4DGL3Q2BqRYyZzuiRVuK/ac
piNPq8CHAPxKrseE2gmfjSSSoKQQD6qqe9kTDIp96m7tM6yt8/qNukbbVbgms0XRNcoXXyXrunEc
xINh+puZB2wLMiBl1yrKNMt/iOXrXS6RiuB+BRx82OHUNoLE4YOqU+7P4kMKsHms0jy+ZdwwR69s
o0o9QIDfqHwjkvxQALcNo/kzr4HhjGtsrD0XKqe+jhfFi14W5BDCR6N6FT19kClrqx+lw/e7NfP3
L69WNGkey0SfEMpg8IsF4RsaPwcEq158XJsbZJGq8bRxr0StAImZHvB5vkgrb7YpcMdv/xB17LIE
hQd2xe713G6rXscEZmfrExsBOPs1TsQhrJjaW++2eF+CtdQIFPpXfQuLwpUwfEvGTQ5pltjnmwaK
Sc38d+UvXM2VucFK7iwCDVWy2GJ0p6jeVYoy804k5TXQuPIFKn8xwjOXxUxqr2Q3vszhye98rRZq
Gng/x7pinGLOEEBEnUlXUm96lR8ztQY3rET6361qwEXVUMV5Nxo2zXwIHvWn4oZehIxyf7Mn+21v
5KOlMOVtVf+cgnqhw89cyaqj8+mumdO7F2TQTyl4cxyxXDff6ASZbKwXYCS7w1YhL1GbDEqQEd2v
MI/KmcW97PZu+MoUPcPKerpxZCIXL+eETZkpVH6XRMATTAFOjfkkLZU505ra9Tdci0gGGoNmMBaq
lkS5xvilagjE+/3q1YoYLTzS243jw+Kmg1tDrISWCqQLe0aYyMW5+ux+4IMf5HgbnT6QteXCV2Tf
0h/xZZjPP/Aa8CbjD7thQqUSKRcksO09eKTrkX8lPQcDgVz8u+CjpmodnF26ZUHgjcJetfajXyLQ
zLSYXBSYdgKqgRWGu2Fn4R0ypirl+ky6P0s7UCEIHQfPajmfvxwu/YDUIBebZPnGCc8hukThiM7k
RhOOMf2kxDhRLPZT3hXN7cdGtQdAG3UtBnPbB+axCuTZybklP2V/rcH+TPH/Le5s+4POiW7iKQ8C
6xm+iBa4jcuRKqV5K9wV1dHRa/Sj11lKEQEmMORJcJr/uDsJcwWlve7dH4seMJqx0y0RJtJ8OaoU
n3tUZj3+vtQFT706jBh4HeLHw+co+HV9FlHnamk/DebUI9U2Gyh6FVGC6Os1j8Gi1OKsrWHAzOHC
QbKhTtm4Y0TamPxXDTttiVmK/DnTLrHeuH7miIMPyIxiZK8nPXco73qzjJMObj7opN/vmndDG1Re
y8zSFnIn4bWAhDvttfiXBI8sBBSnMqder91EtLolc9CiZcXa2aq+GwyVk4RmFzIixvr8baE16rlF
VKIawwyg4qx/eYWYiS2jFSmQcGrkNSZqiRhsixH0Iwd81EsqLQ2jqer5nrb5YJYGKdcHBwq6qU1L
bdng0TrHUMZp94Sgk10yHA8lB6MVsR32ZL8JH3LvtxPL3JHp/ng/kt6CbdOvjdKi5UqPSqsotpZz
2Z5js8/fVu1YY+h155rC+cmjnnLTOMuLkVFBNDd81qFtRhaUEh+yD7Wpe6NSzpGnYoR0sjohyda/
WfhI7qH+yKlgEIOtdnQBvS68gCqqaR409MK0varDwzi2WY4B6R7Ht2pzHziK+I7MzbpTwcjVGT4y
Bl9u+TiSqZVawCCqCvJHhJ7G4UpsFwx6izCXjJjinXIKUFfcFcEhH5v+IYNQ+zBSbxEiRI5EJ9wM
IURylZqrka2oHN1i5qI2PaaFVGTp6OzTWJy5nNfJV56nhKvbcUGVunjaltxHIcJ0OkH++JC4ob6M
zJg8+U+QPDP3l5pAVqhv2H0szt8x+/TVem5nWq3ah2mw7qCsfLv054JSRQz/6waKYCmx0pRyrR5M
TW50GBfP7A+ch79uZFBTGPqOIOmWqjd/qHjIaGx1OaytWHWA1wXe+7beo2weMWOU9meOt8muGGDH
gFAtX/fZiHnjc9WwNkEFzpKsYllkL+HnRnVl01g4PYMb81Dm/Ph2XrkVin4StGu3u/9QOKOnpUQW
ezZVACTx1oHhK7u9x6nFXZq6d3l7Q7XHYqlUbyLn72vG+vH8usz6ipyKOcj8NMHDW0E0bjjH1O5+
I4I0abVYKAWofKcwDTggechGSEhnCMhvjYFoFBocLLOZ6OXaxthU8cYWBgbvRnTW4d0b6T/r4eeW
dXxDS1+AfCLSq+5zQ9rSmw9lcSwaQYqMBBSb61BorodRDCx+wn0vErT99eqKeLiFeNL3dSTHVOkK
2Fy0NyRS5qGAbZdGGEdDQ6wNk0VJa4n1SjePKQ5Q3UuMlvaZm/wvvus5dwuAO35YkaBxU/lzFai7
AV2sbVOXgXVEMS1F4OzzuXLTAzeo193MxMvbYtPKgI7uOMBkWuvV3f//z8tIp3V/QHSgPMH7FegJ
O8eJf81KxAboq3sEx0z5/nJFGB+l2EB0CEqGZEd+yHoO2uA0upZUXGCLD+klLbNfRcc6tSEJeha5
pWMhds2oMhFmVfmVr59Gx7DciK76LGCk5q/yyDRMoCOyTbzvCabS9sP9ZdeNwvePXsCB2iMOeaKK
F7SUvYQEXBLFCc+OUI99tbWglDRYLDQ24dtaMuC8TkSl3SboLQfKA09dUb7RLdd4HxBltYx47ea6
aLvr4/jKhdQb14P9lopoRjTL4Mabx5KyMVbn6tJfgi09NbTHLo9U8hlGYGrhRqYlzwitWcLb8SE8
RSHnbOb8ou7MOXar8yGzSL48zmFL8MUajbQpaEZbbr4lRbO7yHPp6gVekqMEfAP3IqszJVycKxjp
kzB6Zq86A2RJzT8KbQHi5FyhHTwDGfr/LVC0y+O4rbmIUXpQz8mDPbQbGeTUtJthCTMEgHd/8Q9h
0LWmNTXHErOIdSKbuV+6kTpSsSzNX+M6TXY3TxQnnezvi6TIe8Uxo/PPimN+hhdZ4qhOnDlC6SDa
ZqfBf4GGCsVE4bjEs+dZjX5G3pd9RX/5GsHJkeTs6VemuZn1JHTfsKFooglk9AxAnvmctBfEYbQL
FhakGJcmeG/3f2w1zZ9czdGtb1oJ0kNpewZYW7WCLHw1TwGb/Q8sMhduPKYL2uSiwnB3gDEtXkuk
kg7+nZDHC3D4sE6CG//mtSUX2Y2ZizhCyQczpdgYVi1FVQbtkgzSG0aFCIXGBBl5Se3N8LcN+QDi
2BrdMKfIS2pATA3fLkhFh5QN1VhZwGypByq2CTZfaO5Mb/GDkgAIbbK+hcc/xqcAr9G+9BG6H9PM
YORGIENuSEwuPt74ZooHaci6GxH3F0u3hOitDYwJ6Y9xbWyAAvGu/6Ut6Bi5dGWrnN2BuBBzZF+K
6AfOE34d0grDkoOzi39ts2aJajyXhKUmmCwqMT0K4z9Q43cqFqn9jLABS2mUYdXF1uYIthEcydBg
Yi8VT+2fnU9dSlfoKCAsqfkZvQ8U7x3DrB8O9ZnqB7YR8wO7vfzT3YAK7FwS5L6UI16QMbwjNn9Y
HN9FTd4BcBAtiQ5fJi8siWL5k6HqZxxvBe8+B/+zvkp2YTC/ro7xHObCXRK8l4jNCe67LD0KDUMi
2rqBS8ryx60gF49o5OHS+vIFjilHmgVRZGAE2BHp9b1N3K7/H8ecdSTRy2eZpneRzFaePT1tN4nP
ipe6SlkTZW15KxjqV9xSJt7I92K1j4SoedtVA+8eYHiaKYQMUxXe2kgJ3K5SCRZNBoqFn9iRMpza
Md6Z8fv5Y+4SruVFz4GYlfvHCcaOz+gQymEQHP7oHy6UrFh+osh9qeTwcFJBZr9qPfUKvcse0ner
8fhr52F2AbOTuknv7O9SE8MxqMOY3RE7DklmU6MTff6SykXT1MD67C0TkEtCgaF8jj+1Q7o1qIjI
WK9Xm3yYuVLpjgiLEnNUl+U9b58yQiZpC04L9x9SQBhUaQqkgXmhaxX0lKIBsysfEROqKEODAwZN
Vc3XFaSJmXVz6O1bkXIpUtbW6hZonysG384zlV3vA8lnrBscraSWbUwDg8sMW27KE9RkU/zNribB
Cmn0pdlbe+QpUkpJIkLVBu4AJ+k6ypjnMLyrs/uy4iMEW9WnmIu0agyGB8iP6RyF7Hv5T9dqVZ7N
9goSD6TQbsaQzjB4E8J6WePlIHNDzLP/+xlKjVlokQwVtgFXauLllozus+/2xEQwrgq3PP3A/Gc9
TlJHBPOTo1CO6xwFA9DdbfO6oQDLtDE49eRIBSTX7zpVGj3PrkOPLzTdB2KgQozfpFe37h+9uNFP
G1TTbqyqlXPTN3zVtROTro+QbkbmMIjoIEwyihmFdnuNfxSLaAVo+HfJXllITi1YD5koxmxBaxKl
B0GoIeH/ahf6YBK2lntoO5cDXOq0wIwR8CtamBYvIBpP+AM18giNy7J9t3z7UxnLAkr8xbSk78xL
xBUlkFon/UgTnhFflE17fqAjdB2Hd7+Xjg9oJXWNQP9ZYgMyGkhrSSLMFlUVHnUupcaidAAeVYlk
S9Z24ef37eC2gRIULgkYC85WX2/8CcRq7FVT6c85zUQMWdLpet6VJXlDTZbvPHt7iVR8XULDv99o
v9qgbMG6ytVIvI/krYsiivGWENdznQvpLMvnbrBN1rYoETtEntRiGGAlPmZOUrWGaiatkdPyOFkd
wYqqu/iPvHr2/o/bMVr9VbusqZXEfdhJImS1Ea8sDKKja3Dw0owBoFcgol1Vn/0fj4YYYemsDJQd
G4Ewg0IajHjtz3UoPqSjLVNAMO92dNcKqO5duBbutuJ5MlIC07SJlwTozCFH9/o+jtmbDeLIhwMC
aj9EwMoiuihOQJAvDMjawrtj3VlUp0y3/qok25OxOsZ2YPF7SWjUyjXnJVn8Vk3ZtvUF3m80BrWw
EsDqS71VAkE3QZIXiAh5yKgu9dqvCl98hBz37RyAmyIitF/TVmgSyrV16LatevNkK3RYyVQ8C1pq
DYeF0j5WkQJ3P8hMmRl0HML1Jrg2qZh4qUscGi+Tw+ZKEp7xF5Urltdl+bfQIVMdHUgXkLgyUxwK
X9TyyQqeA+vg4PyGghvia2OQn2mCxu4wuwKMt2oICxA/3l6cxBLPzuSYiB9472A8+uDCF/y/AnOn
DQx+Yo5CEr8sZjSf981uIyYcGBK3omiq2b6t9NjnveN0kvi63ESS3sJOWTS9/14p9+GH9xfm8BD2
qSqDArackOeoTjLVRV74UZ4wrtaTzPhg4N9O11u/Wrgb3EbvS3eLI/AkgeP8ftBtP+Evpb79okvz
GH3WjwvDVpS06JzQ2/j5BUlpyVR7R8PyUc1GlOcFZzU5ocpL7iZdPzylqnjP8fuw7vEn/eIcbulR
CLzLgYt9dPpqYn+iqAy3Fzzdd9K9KVgjc0MT9N5eKOelc8FDSRAEruQcviurM23bV9OpYk4/q8jE
+mMO3g+71LmrD/svKvTRlC1z59RdSZltmbw9Xt0ZZRYBKhDWIOzQhtRAkKfWK/Z6kE4Wsbu4ymO8
duKgVya4FYQtC/6vG7DNbRknevY3pc7wVlwXhibHkdGQaNzneAHjONxmrl02aT14/U0gwKOud4Tx
eSTy+GvSatRxaT+uAGBSx9jzU4EteZc8EHCnESeJtXc/5jXShT32VDmuFds72XilnIvAKlBD6B5E
ymznczxzZP+DsG0dG0wkPPCXrnkSnjsEfGQ40Y5vnBNRRIHzCkzdFbQJSMeyQNtMzAIUsh5zMcMi
Sb2YzRsVaV76qxXdh+Ww48BG+26H3lA/p1TVzBzEdNqK2/TAsbA38NjfWRYupYd7T56bQusrdSMI
C6Nk+uubYUJb3yJN1IKRIarvfTeGSwCl8c61x7tzdfdeVB+GhrYGn2+cMiFiYNx4FVaNaMVA9E60
rOhT8vFDbrNqO/3katBSUDi22J7QCTo02+QFK0O9jD0oWLnDAuGLonMcH0TgYh4MlM0dmtlGN4WC
i/tAMdr0p13N1bbrNCQYRDldUGh1Fqw+tjmGdoXV5A7JYKw7fSZRgOZINTBfQE0XI9ELdsfaX0KL
BsH9OTHUk500Mz2attCnok7RQEe+t4Vw/iDmyoxq2E8XYj5q1gUVbQNjADB1Vg6Dzy1731Am0M6v
A7TefEV9MMK9UM9CdUkfLQizU4NOEq3XED13lmz+Aj/XOX7lTVv0YDpqOQ0OeL3FzALVmbdy8S8y
/6vOQgVfozMhks09DAbXohZokRhOI+OZWJ/3zbQsALObSMnFVYwP9ecWO5Wq9ylBRBNEDLEhkisE
+H879Oq85o0gUMXzHM8W2wOW1HgMQOMhEsqN1lXuPshcpdVtQI2tsVMvDc9KgJN5C1hAofwxT4LY
ptYb2muRJMh4UMNmK+Uaso5pU3vrjj260lBUuoDOnXIDIP202dJjdl5Q02f2IYVwrP7HCOQr+szc
TZ4ZfhGWpfdKXWma360iWuorbhjFrWwhL8USLpjDguWJ27HPzF4aE+POD27EU86QP6zD2aJwdaf2
Zdi8JpfmDSQMEYPR+JUBReEFCzfjQLaZC6jnLxXVZFQH4xXWXG5ri9iH6F+KEqndPoManRtFRLGG
a12U88sTEdB9dOO8muImo00YNjDP/G+6mLotaLaoJ83BwGrxt6GR9HQoZPRdcb2wK5sIF113kIg1
dx+BT9ejin1ALx+2aLY9xBFLm2x/5bzNhYQkftbF3BuPJr4vXKf6kGTYnGTSRVzTNKtQZi7Lv+i6
WolnUo05M3BheWrTIkj5UZ/ug42RiP342oaOlVOKarR9aMIS/hi4dcdpUMZ2ww4aj8CSrYVMYbUj
1zuqO5Z/G0Mk7QzJppSoJ41qk0Zm/N2f5ruQmGVRLFDqUv5bDyUM3ALHLsgrcqO9QZjHrDDblZzr
Nud0t4MQe/myfqImKRdWrRwzRs52NdQHqnlED1l0SWlcLgWklwdks9NmHJZjdEyzfm/TUKUeQZ1+
8gBIFvcL8hbBfcG7019Kcs3fKvF0hw3liG7ax5PH3kZWPrqOgMA=
`protect end_protected

