------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   / 
-- /___/  \  /    Vendor: Xilinx 
-- \   \   \/     Version : 3.6
--  \   \         Application : 7 Series FPGAs Transceivers Wizard 
--  /   /         Filename : gtwizard_0_gt_usrclk_source.vhd
-- /___/   /\      
-- \   \  /  \ 
--  \___\/\___\ 
--
--
-- Module gtwizard_0_GT_USRCLK_SOURCE (for use with GTs)
-- Generated by Xilinx 7 Series FPGAs Transceivers 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;

--***********************************Entity Declaration*******************************
entity gtwizard_0_GT_USRCLK_SOURCE is
port
(
    txusrclk2_in : in std_logic;
    txusrclk_in : in std_logic;
    GT0_TXUSRCLK_OUT             : out std_logic;
    GT0_TXUSRCLK2_OUT            : out std_logic;
    GT0_TXOUTCLK_IN              : in  std_logic;
    GT0_TXCLK_LOCK_OUT           : out std_logic;
    GT0_TX_MMCM_RESET_IN         : in std_logic;
    GT0_RXUSRCLK_OUT             : out std_logic;
    GT0_RXUSRCLK2_OUT            : out std_logic;
    GT0_RXOUTCLK_IN              : in  std_logic;
    GT0_RXCLK_LOCK_OUT           : out std_logic;
    GT0_RX_MMCM_RESET_IN         : in std_logic;
 
    GT1_TXUSRCLK_OUT             : out std_logic;
    GT1_TXUSRCLK2_OUT            : out std_logic;
    GT1_TXOUTCLK_IN              : in  std_logic;
    GT1_TXCLK_LOCK_OUT           : out std_logic;
    GT1_TX_MMCM_RESET_IN         : in std_logic;
    GT1_RXUSRCLK_OUT             : out std_logic;
    GT1_RXUSRCLK2_OUT            : out std_logic;
    GT1_RXOUTCLK_IN              : in  std_logic;
    GT1_RXCLK_LOCK_OUT           : out std_logic;
    GT1_RX_MMCM_RESET_IN         : in std_logic;
 
    GT2_TXUSRCLK_OUT             : out std_logic;
    GT2_TXUSRCLK2_OUT            : out std_logic;
    GT2_TXOUTCLK_IN              : in  std_logic;
    GT2_TXCLK_LOCK_OUT           : out std_logic;
    GT2_TX_MMCM_RESET_IN         : in std_logic;
    GT2_RXUSRCLK_OUT             : out std_logic;
    GT2_RXUSRCLK2_OUT            : out std_logic;
    GT2_RXOUTCLK_IN              : in  std_logic;
    GT2_RXCLK_LOCK_OUT           : out std_logic;
    GT2_RX_MMCM_RESET_IN         : in std_logic;
 
    GT3_TXUSRCLK_OUT             : out std_logic;
    GT3_TXUSRCLK2_OUT            : out std_logic;
    GT3_TXOUTCLK_IN              : in  std_logic;
    GT3_TXCLK_LOCK_OUT           : out std_logic;
    GT3_TX_MMCM_RESET_IN         : in std_logic;
    GT3_RXUSRCLK_OUT             : out std_logic;
    GT3_RXUSRCLK2_OUT            : out std_logic;
    GT3_RXOUTCLK_IN              : in  std_logic;
    GT3_RXCLK_LOCK_OUT           : out std_logic;
    GT3_RX_MMCM_RESET_IN         : in std_logic;
 
    GT4_TXUSRCLK_OUT             : out std_logic;
    GT4_TXUSRCLK2_OUT            : out std_logic;
    GT4_TXOUTCLK_IN              : in  std_logic;
    GT4_TXCLK_LOCK_OUT           : out std_logic;
    GT4_TX_MMCM_RESET_IN         : in std_logic;
    GT4_RXUSRCLK_OUT             : out std_logic;
    GT4_RXUSRCLK2_OUT            : out std_logic;
    GT4_RXOUTCLK_IN              : in  std_logic;
    GT4_RXCLK_LOCK_OUT           : out std_logic;
    GT4_RX_MMCM_RESET_IN         : in std_logic;
 
    GT5_TXUSRCLK_OUT             : out std_logic;
    GT5_TXUSRCLK2_OUT            : out std_logic;
    GT5_TXOUTCLK_IN              : in  std_logic;
    GT5_TXCLK_LOCK_OUT           : out std_logic;
    GT5_TX_MMCM_RESET_IN         : in std_logic;
    GT5_RXUSRCLK_OUT             : out std_logic;
    GT5_RXUSRCLK2_OUT            : out std_logic;
    GT5_RXOUTCLK_IN              : in  std_logic;
    GT5_RXCLK_LOCK_OUT           : out std_logic;
    GT5_RX_MMCM_RESET_IN         : in std_logic;
 
    GT6_TXUSRCLK_OUT             : out std_logic;
    GT6_TXUSRCLK2_OUT            : out std_logic;
    GT6_TXOUTCLK_IN              : in  std_logic;
    GT6_TXCLK_LOCK_OUT           : out std_logic;
    GT6_TX_MMCM_RESET_IN         : in std_logic;
    GT6_RXUSRCLK_OUT             : out std_logic;
    GT6_RXUSRCLK2_OUT            : out std_logic;
    GT6_RXOUTCLK_IN              : in  std_logic;
    GT6_RXCLK_LOCK_OUT           : out std_logic;
    GT6_RX_MMCM_RESET_IN         : in std_logic;
 
    GT7_TXUSRCLK_OUT             : out std_logic;
    GT7_TXUSRCLK2_OUT            : out std_logic;
    GT7_TXOUTCLK_IN              : in  std_logic;
    GT7_TXCLK_LOCK_OUT           : out std_logic;
    GT7_TX_MMCM_RESET_IN         : in std_logic;
    GT7_RXUSRCLK_OUT             : out std_logic;
    GT7_RXUSRCLK2_OUT            : out std_logic;
    GT7_RXOUTCLK_IN              : in  std_logic;
    GT7_RXCLK_LOCK_OUT           : out std_logic;
    GT7_RX_MMCM_RESET_IN         : in std_logic;
 
    GT8_TXUSRCLK_OUT             : out std_logic;
    GT8_TXUSRCLK2_OUT            : out std_logic;
    GT8_TXOUTCLK_IN              : in  std_logic;
    GT8_TXCLK_LOCK_OUT           : out std_logic;
    GT8_TX_MMCM_RESET_IN         : in std_logic;
    GT8_RXUSRCLK_OUT             : out std_logic;
    GT8_RXUSRCLK2_OUT            : out std_logic;
    GT8_RXOUTCLK_IN              : in  std_logic;
    GT8_RXCLK_LOCK_OUT           : out std_logic;
    GT8_RX_MMCM_RESET_IN         : in std_logic;
 
    GT9_TXUSRCLK_OUT             : out std_logic;
    GT9_TXUSRCLK2_OUT            : out std_logic;
    GT9_TXOUTCLK_IN              : in  std_logic;
    GT9_TXCLK_LOCK_OUT           : out std_logic;
    GT9_TX_MMCM_RESET_IN         : in std_logic;
    GT9_RXUSRCLK_OUT             : out std_logic;
    GT9_RXUSRCLK2_OUT            : out std_logic;
    GT9_RXOUTCLK_IN              : in  std_logic;
    GT9_RXCLK_LOCK_OUT           : out std_logic;
    GT9_RX_MMCM_RESET_IN         : in std_logic;
 
    GT10_TXUSRCLK_OUT             : out std_logic;
    GT10_TXUSRCLK2_OUT            : out std_logic;
    GT10_TXOUTCLK_IN              : in  std_logic;
    GT10_TXCLK_LOCK_OUT           : out std_logic;
    GT10_TX_MMCM_RESET_IN         : in std_logic;
    GT10_RXUSRCLK_OUT             : out std_logic;
    GT10_RXUSRCLK2_OUT            : out std_logic;
    GT10_RXOUTCLK_IN              : in  std_logic;
    GT10_RXCLK_LOCK_OUT           : out std_logic;
    GT10_RX_MMCM_RESET_IN         : in std_logic;
 
    GT11_TXUSRCLK_OUT             : out std_logic;
    GT11_TXUSRCLK2_OUT            : out std_logic;
    GT11_TXOUTCLK_IN              : in  std_logic;
    GT11_TXCLK_LOCK_OUT           : out std_logic;
    GT11_TX_MMCM_RESET_IN         : in std_logic;
    GT11_RXUSRCLK_OUT             : out std_logic;
    GT11_RXUSRCLK2_OUT            : out std_logic;
    GT11_RXOUTCLK_IN              : in  std_logic;
    GT11_RXCLK_LOCK_OUT           : out std_logic;
    GT11_RX_MMCM_RESET_IN         : in std_logic;
 
    GT12_TXUSRCLK_OUT             : out std_logic;
    GT12_TXUSRCLK2_OUT            : out std_logic;
    GT12_TXOUTCLK_IN              : in  std_logic;
    GT12_TXCLK_LOCK_OUT           : out std_logic;
    GT12_TX_MMCM_RESET_IN         : in std_logic;
    GT12_RXUSRCLK_OUT             : out std_logic;
    GT12_RXUSRCLK2_OUT            : out std_logic;
    GT12_RXOUTCLK_IN              : in  std_logic;
    GT12_RXCLK_LOCK_OUT           : out std_logic;
    GT12_RX_MMCM_RESET_IN         : in std_logic;
 
    GT13_TXUSRCLK_OUT             : out std_logic;
    GT13_TXUSRCLK2_OUT            : out std_logic;
    GT13_TXOUTCLK_IN              : in  std_logic;
    GT13_TXCLK_LOCK_OUT           : out std_logic;
    GT13_TX_MMCM_RESET_IN         : in std_logic;
    GT13_RXUSRCLK_OUT             : out std_logic;
    GT13_RXUSRCLK2_OUT            : out std_logic;
    GT13_RXOUTCLK_IN              : in  std_logic;
    GT13_RXCLK_LOCK_OUT           : out std_logic;
    GT13_RX_MMCM_RESET_IN         : in std_logic;
 
    GT14_TXUSRCLK_OUT             : out std_logic;
    GT14_TXUSRCLK2_OUT            : out std_logic;
    GT14_TXOUTCLK_IN              : in  std_logic;
    GT14_TXCLK_LOCK_OUT           : out std_logic;
    GT14_TX_MMCM_RESET_IN         : in std_logic;
    GT14_RXUSRCLK_OUT             : out std_logic;
    GT14_RXUSRCLK2_OUT            : out std_logic;
    GT14_RXOUTCLK_IN              : in  std_logic;
    GT14_RXCLK_LOCK_OUT           : out std_logic;
    GT14_RX_MMCM_RESET_IN         : in std_logic;
 
    GT15_TXUSRCLK_OUT             : out std_logic;
    GT15_TXUSRCLK2_OUT            : out std_logic;
    GT15_TXOUTCLK_IN              : in  std_logic;
    GT15_TXCLK_LOCK_OUT           : out std_logic;
    GT15_TX_MMCM_RESET_IN         : in std_logic;
    GT15_RXUSRCLK_OUT             : out std_logic;
    GT15_RXUSRCLK2_OUT            : out std_logic;
    GT15_RXOUTCLK_IN              : in  std_logic;
    GT15_RXCLK_LOCK_OUT           : out std_logic;
    GT15_RX_MMCM_RESET_IN         : in std_logic;
 
    GT16_TXUSRCLK_OUT             : out std_logic;
    GT16_TXUSRCLK2_OUT            : out std_logic;
    GT16_TXOUTCLK_IN              : in  std_logic;
    GT16_TXCLK_LOCK_OUT           : out std_logic;
    GT16_TX_MMCM_RESET_IN         : in std_logic;
    GT16_RXUSRCLK_OUT             : out std_logic;
    GT16_RXUSRCLK2_OUT            : out std_logic;
    GT16_RXOUTCLK_IN              : in  std_logic;
    GT16_RXCLK_LOCK_OUT           : out std_logic;
    GT16_RX_MMCM_RESET_IN         : in std_logic;
 
    GT17_TXUSRCLK_OUT             : out std_logic;
    GT17_TXUSRCLK2_OUT            : out std_logic;
    GT17_TXOUTCLK_IN              : in  std_logic;
    GT17_TXCLK_LOCK_OUT           : out std_logic;
    GT17_TX_MMCM_RESET_IN         : in std_logic;
    GT17_RXUSRCLK_OUT             : out std_logic;
    GT17_RXUSRCLK2_OUT            : out std_logic;
    GT17_RXOUTCLK_IN              : in  std_logic;
    GT17_RXCLK_LOCK_OUT           : out std_logic;
    GT17_RX_MMCM_RESET_IN         : in std_logic;
 
    GT18_TXUSRCLK_OUT             : out std_logic;
    GT18_TXUSRCLK2_OUT            : out std_logic;
    GT18_TXOUTCLK_IN              : in  std_logic;
    GT18_TXCLK_LOCK_OUT           : out std_logic;
    GT18_TX_MMCM_RESET_IN         : in std_logic;
    GT18_RXUSRCLK_OUT             : out std_logic;
    GT18_RXUSRCLK2_OUT            : out std_logic;
    GT18_RXOUTCLK_IN              : in  std_logic;
    GT18_RXCLK_LOCK_OUT           : out std_logic;
    GT18_RX_MMCM_RESET_IN         : in std_logic;
 
    GT19_TXUSRCLK_OUT             : out std_logic;
    GT19_TXUSRCLK2_OUT            : out std_logic;
    GT19_TXOUTCLK_IN              : in  std_logic;
    GT19_TXCLK_LOCK_OUT           : out std_logic;
    GT19_TX_MMCM_RESET_IN         : in std_logic;
    GT19_RXUSRCLK_OUT             : out std_logic;
    GT19_RXUSRCLK2_OUT            : out std_logic;
    GT19_RXOUTCLK_IN              : in  std_logic;
    GT19_RXCLK_LOCK_OUT           : out std_logic;
    GT19_RX_MMCM_RESET_IN         : in std_logic;
 
    GT20_TXUSRCLK_OUT             : out std_logic;
    GT20_TXUSRCLK2_OUT            : out std_logic;
    GT20_TXOUTCLK_IN              : in  std_logic;
    GT20_TXCLK_LOCK_OUT           : out std_logic;
    GT20_TX_MMCM_RESET_IN         : in std_logic;
    GT20_RXUSRCLK_OUT             : out std_logic;
    GT20_RXUSRCLK2_OUT            : out std_logic;
    GT20_RXOUTCLK_IN              : in  std_logic;
    GT20_RXCLK_LOCK_OUT           : out std_logic;
    GT20_RX_MMCM_RESET_IN         : in std_logic;
 
    GT21_TXUSRCLK_OUT             : out std_logic;
    GT21_TXUSRCLK2_OUT            : out std_logic;
    GT21_TXOUTCLK_IN              : in  std_logic;
    GT21_TXCLK_LOCK_OUT           : out std_logic;
    GT21_TX_MMCM_RESET_IN         : in std_logic;
    GT21_RXUSRCLK_OUT             : out std_logic;
    GT21_RXUSRCLK2_OUT            : out std_logic;
    GT21_RXOUTCLK_IN              : in  std_logic;
    GT21_RXCLK_LOCK_OUT           : out std_logic;
    GT21_RX_MMCM_RESET_IN         : in std_logic;
 
    GT22_TXUSRCLK_OUT             : out std_logic;
    GT22_TXUSRCLK2_OUT            : out std_logic;
    GT22_TXOUTCLK_IN              : in  std_logic;
    GT22_TXCLK_LOCK_OUT           : out std_logic;
    GT22_TX_MMCM_RESET_IN         : in std_logic;
    GT22_RXUSRCLK_OUT             : out std_logic;
    GT22_RXUSRCLK2_OUT            : out std_logic;
    GT22_RXOUTCLK_IN              : in  std_logic;
    GT22_RXCLK_LOCK_OUT           : out std_logic;
    GT22_RX_MMCM_RESET_IN         : in std_logic;
 
    GT23_TXUSRCLK_OUT             : out std_logic;
    GT23_TXUSRCLK2_OUT            : out std_logic;
    GT23_TXOUTCLK_IN              : in  std_logic;
    GT23_TXCLK_LOCK_OUT           : out std_logic;
    GT23_TX_MMCM_RESET_IN         : in std_logic;
    GT23_RXUSRCLK_OUT             : out std_logic;
    GT23_RXUSRCLK2_OUT            : out std_logic;
    GT23_RXOUTCLK_IN              : in  std_logic;
    GT23_RXCLK_LOCK_OUT           : out std_logic;
    GT23_RX_MMCM_RESET_IN         : in std_logic;
 
    GT24_TXUSRCLK_OUT             : out std_logic;
    GT24_TXUSRCLK2_OUT            : out std_logic;
    GT24_TXOUTCLK_IN              : in  std_logic;
    GT24_TXCLK_LOCK_OUT           : out std_logic;
    GT24_TX_MMCM_RESET_IN         : in std_logic;
    GT24_RXUSRCLK_OUT             : out std_logic;
    GT24_RXUSRCLK2_OUT            : out std_logic;
    GT24_RXOUTCLK_IN              : in  std_logic;
    GT24_RXCLK_LOCK_OUT           : out std_logic;
    GT24_RX_MMCM_RESET_IN         : in std_logic;
 
    GT25_TXUSRCLK_OUT             : out std_logic;
    GT25_TXUSRCLK2_OUT            : out std_logic;
    GT25_TXOUTCLK_IN              : in  std_logic;
    GT25_TXCLK_LOCK_OUT           : out std_logic;
    GT25_TX_MMCM_RESET_IN         : in std_logic;
    GT25_RXUSRCLK_OUT             : out std_logic;
    GT25_RXUSRCLK2_OUT            : out std_logic;
    GT25_RXOUTCLK_IN              : in  std_logic;
    GT25_RXCLK_LOCK_OUT           : out std_logic;
    GT25_RX_MMCM_RESET_IN         : in std_logic;
 
    GT26_TXUSRCLK_OUT             : out std_logic;
    GT26_TXUSRCLK2_OUT            : out std_logic;
    GT26_TXOUTCLK_IN              : in  std_logic;
    GT26_TXCLK_LOCK_OUT           : out std_logic;
    GT26_TX_MMCM_RESET_IN         : in std_logic;
    GT26_RXUSRCLK_OUT             : out std_logic;
    GT26_RXUSRCLK2_OUT            : out std_logic;
    GT26_RXOUTCLK_IN              : in  std_logic;
    GT26_RXCLK_LOCK_OUT           : out std_logic;
    GT26_RX_MMCM_RESET_IN         : in std_logic;
 
    GT27_TXUSRCLK_OUT             : out std_logic;
    GT27_TXUSRCLK2_OUT            : out std_logic;
    GT27_TXOUTCLK_IN              : in  std_logic;
    GT27_TXCLK_LOCK_OUT           : out std_logic;
    GT27_TX_MMCM_RESET_IN         : in std_logic;
    GT27_RXUSRCLK_OUT             : out std_logic;
    GT27_RXUSRCLK2_OUT            : out std_logic;
    GT27_RXOUTCLK_IN              : in  std_logic;
    GT27_RXCLK_LOCK_OUT           : out std_logic;
    GT27_RX_MMCM_RESET_IN         : in std_logic;
 
    GT28_TXUSRCLK_OUT             : out std_logic;
    GT28_TXUSRCLK2_OUT            : out std_logic;
    GT28_TXOUTCLK_IN              : in  std_logic;
    GT28_TXCLK_LOCK_OUT           : out std_logic;
    GT28_TX_MMCM_RESET_IN         : in std_logic;
    GT28_RXUSRCLK_OUT             : out std_logic;
    GT28_RXUSRCLK2_OUT            : out std_logic;
    GT28_RXOUTCLK_IN              : in  std_logic;
    GT28_RXCLK_LOCK_OUT           : out std_logic;
    GT28_RX_MMCM_RESET_IN         : in std_logic;
 
    GT29_TXUSRCLK_OUT             : out std_logic;
    GT29_TXUSRCLK2_OUT            : out std_logic;
    GT29_TXOUTCLK_IN              : in  std_logic;
    GT29_TXCLK_LOCK_OUT           : out std_logic;
    GT29_TX_MMCM_RESET_IN         : in std_logic;
    GT29_RXUSRCLK_OUT             : out std_logic;
    GT29_RXUSRCLK2_OUT            : out std_logic;
    GT29_RXOUTCLK_IN              : in  std_logic;
    GT29_RXCLK_LOCK_OUT           : out std_logic;
    GT29_RX_MMCM_RESET_IN         : in std_logic;
 
    GT30_TXUSRCLK_OUT             : out std_logic;
    GT30_TXUSRCLK2_OUT            : out std_logic;
    GT30_TXOUTCLK_IN              : in  std_logic;
    GT30_TXCLK_LOCK_OUT           : out std_logic;
    GT30_TX_MMCM_RESET_IN         : in std_logic;
    GT30_RXUSRCLK_OUT             : out std_logic;
    GT30_RXUSRCLK2_OUT            : out std_logic;
    GT30_RXOUTCLK_IN              : in  std_logic;
    GT30_RXCLK_LOCK_OUT           : out std_logic;
    GT30_RX_MMCM_RESET_IN         : in std_logic;
 
    GT31_TXUSRCLK_OUT             : out std_logic;
    GT31_TXUSRCLK2_OUT            : out std_logic;
    GT31_TXOUTCLK_IN              : in  std_logic;
    GT31_TXCLK_LOCK_OUT           : out std_logic;
    GT31_TX_MMCM_RESET_IN         : in std_logic;
    GT31_RXUSRCLK_OUT             : out std_logic;
    GT31_RXUSRCLK2_OUT            : out std_logic;
    GT31_RXOUTCLK_IN              : in  std_logic;
    GT31_RXCLK_LOCK_OUT           : out std_logic;
    GT31_RX_MMCM_RESET_IN         : in std_logic;
    Q2_CLK0_GTREFCLK_PAD_N_IN               : in   std_logic;
    Q2_CLK0_GTREFCLK_PAD_P_IN               : in   std_logic;
    Q2_CLK0_GTREFCLK_OUT                    : out  std_logic;
    Q5_CLK0_GTREFCLK_PAD_N_IN               : in   std_logic;
    Q5_CLK0_GTREFCLK_PAD_P_IN               : in   std_logic;
    Q5_CLK0_GTREFCLK_OUT                    : out  std_logic;
    Q7_CLK0_GTREFCLK_PAD_N_IN               : in   std_logic;
    Q7_CLK0_GTREFCLK_PAD_P_IN               : in   std_logic;
    Q7_CLK0_GTREFCLK_OUT                    : out  std_logic
);


end gtwizard_0_GT_USRCLK_SOURCE;

architecture RTL of gtwizard_0_GT_USRCLK_SOURCE is

component GTWIZARD_0_CLOCK_MODULE is
generic
(
    MULT                : real              := 2.0;
    DIVIDE              : integer           := 2;    
    CLK_PERIOD          : real              := 6.4;    
    OUT0_DIVIDE         : real              := 2.0;
    OUT1_DIVIDE         : integer           := 2;
    OUT2_DIVIDE         : integer           := 2;
    OUT3_DIVIDE         : integer           := 2
);
port
 (-- Clock in ports
  CLK_IN           : in     std_logic;
  -- Clock out ports
  CLK0_OUT          : out    std_logic;
  CLK1_OUT          : out    std_logic;
  CLK2_OUT          : out    std_logic;
  CLK3_OUT          : out    std_logic;
  -- Status and control signals
  MMCM_RESET_IN     : in     std_logic;
  MMCM_LOCKED_OUT   : out    std_logic
 );
end component;

--*********************************Wire Declarations**********************************

    signal   tied_to_ground_i     :   std_logic;
    signal   tied_to_vcc_i        :   std_logic;
 
    signal   gt0_txoutclk_i :   std_logic;
    signal   gt0_rxoutclk_i :   std_logic;
 
    signal   gt1_txoutclk_i :   std_logic;
    signal   gt1_rxoutclk_i :   std_logic;
 
    signal   gt2_txoutclk_i :   std_logic;
    signal   gt2_rxoutclk_i :   std_logic;
 
    signal   gt3_txoutclk_i :   std_logic;
    signal   gt3_rxoutclk_i :   std_logic;
 
    signal   gt4_txoutclk_i :   std_logic;
    signal   gt4_rxoutclk_i :   std_logic;
 
    signal   gt5_txoutclk_i :   std_logic;
    signal   gt5_rxoutclk_i :   std_logic;
 
    signal   gt6_txoutclk_i :   std_logic;
    signal   gt6_rxoutclk_i :   std_logic;
 
    signal   gt7_txoutclk_i :   std_logic;
    signal   gt7_rxoutclk_i :   std_logic;
 
    signal   gt8_txoutclk_i :   std_logic;
    signal   gt8_rxoutclk_i :   std_logic;
 
    signal   gt9_txoutclk_i :   std_logic;
    signal   gt9_rxoutclk_i :   std_logic;
 
    signal   gt10_txoutclk_i :   std_logic;
    signal   gt10_rxoutclk_i :   std_logic;
 
    signal   gt11_txoutclk_i :   std_logic;
    signal   gt11_rxoutclk_i :   std_logic;
 
    signal   gt12_txoutclk_i :   std_logic;
    signal   gt12_rxoutclk_i :   std_logic;
 
    signal   gt13_txoutclk_i :   std_logic;
    signal   gt13_rxoutclk_i :   std_logic;
 
    signal   gt14_txoutclk_i :   std_logic;
    signal   gt14_rxoutclk_i :   std_logic;
 
    signal   gt15_txoutclk_i :   std_logic;
    signal   gt15_rxoutclk_i :   std_logic;
 
    signal   gt16_txoutclk_i :   std_logic;
    signal   gt16_rxoutclk_i :   std_logic;
 
    signal   gt17_txoutclk_i :   std_logic;
    signal   gt17_rxoutclk_i :   std_logic;
 
    signal   gt18_txoutclk_i :   std_logic;
    signal   gt18_rxoutclk_i :   std_logic;
 
    signal   gt19_txoutclk_i :   std_logic;
    signal   gt19_rxoutclk_i :   std_logic;
 
    signal   gt20_txoutclk_i :   std_logic;
    signal   gt20_rxoutclk_i :   std_logic;
 
    signal   gt21_txoutclk_i :   std_logic;
    signal   gt21_rxoutclk_i :   std_logic;
 
    signal   gt22_txoutclk_i :   std_logic;
    signal   gt22_rxoutclk_i :   std_logic;
 
    signal   gt23_txoutclk_i :   std_logic;
    signal   gt23_rxoutclk_i :   std_logic;
 
    signal   gt24_txoutclk_i :   std_logic;
    signal   gt24_rxoutclk_i :   std_logic;
 
    signal   gt25_txoutclk_i :   std_logic;
    signal   gt25_rxoutclk_i :   std_logic;
 
    signal   gt26_txoutclk_i :   std_logic;
    signal   gt26_rxoutclk_i :   std_logic;
 
    signal   gt27_txoutclk_i :   std_logic;
    signal   gt27_rxoutclk_i :   std_logic;
 
    signal   gt28_txoutclk_i :   std_logic;
    signal   gt28_rxoutclk_i :   std_logic;
 
    signal   gt29_txoutclk_i :   std_logic;
    signal   gt29_rxoutclk_i :   std_logic;
 
    signal   gt30_txoutclk_i :   std_logic;
    signal   gt30_rxoutclk_i :   std_logic;
 
    signal   gt31_txoutclk_i :   std_logic;
    signal   gt31_rxoutclk_i :   std_logic;

    attribute syn_noclockbuf : boolean;
    signal   q2_clk0_gtrefclk :   std_logic;
    attribute syn_noclockbuf of q2_clk0_gtrefclk : signal is true;
    signal   q5_clk0_gtrefclk :   std_logic;
    attribute syn_noclockbuf of q5_clk0_gtrefclk : signal is true;
    signal   q7_clk0_gtrefclk :   std_logic;
    attribute syn_noclockbuf of q7_clk0_gtrefclk : signal is true;

    signal  gt0_txusrclk_i                  : std_logic;
    signal  gt0_txusrclk2_i                 : std_logic;
    signal  gt0_rxusrclk_i                  : std_logic;
    signal  gt0_rxusrclk2_i                 : std_logic;
    signal  gt12_txusrclk_i                 : std_logic;
    signal  gt12_txusrclk2_i                : std_logic;
    signal  gt12_rxusrclk_i                 : std_logic;
    signal  gt12_rxusrclk2_i                : std_logic;
    signal  gt24_txusrclk_i                 : std_logic;
    signal  gt24_txusrclk2_i                : std_logic;
    signal  gt24_rxusrclk_i                 : std_logic;
    signal  gt24_rxusrclk2_i                : std_logic;
    signal  txoutclk_mmcm0_locked_i         : std_logic;
    signal  txoutclk_mmcm0_reset_i          : std_logic;
    signal  gt0_txoutclk_to_mmcm_i          : std_logic;
    signal  rxoutclk_mmcm1_locked_i         : std_logic;
    signal  rxoutclk_mmcm1_reset_i          : std_logic;
    signal  gt0_rxoutclk_to_mmcm_i          : std_logic;
    signal  txoutclk_mmcm2_locked_i         : std_logic;
    signal  txoutclk_mmcm2_reset_i          : std_logic;
    signal  gt12_txoutclk_to_mmcm_i         : std_logic;
    signal  rxoutclk_mmcm3_locked_i         : std_logic;
    signal  rxoutclk_mmcm3_reset_i          : std_logic;
    signal  gt12_rxoutclk_to_mmcm_i         : std_logic;
    signal  txoutclk_mmcm4_locked_i         : std_logic;
    signal  txoutclk_mmcm4_reset_i          : std_logic;
    signal  gt24_txoutclk_to_mmcm_i         : std_logic;
    signal  rxoutclk_mmcm5_locked_i         : std_logic;
    signal  rxoutclk_mmcm5_reset_i          : std_logic;
    signal  gt24_rxoutclk_to_mmcm_i         : std_logic;


begin

--*********************************** Beginning of Code *******************************

    --  Static signal Assigments    
    tied_to_ground_i         <= '0';
    tied_to_vcc_i            <= '1';
    gt0_txoutclk_i                               <= GT0_TXOUTCLK_IN;
    gt0_rxoutclk_i                               <= GT0_RXOUTCLK_IN;
    gt1_txoutclk_i                               <= GT1_TXOUTCLK_IN;
    gt1_rxoutclk_i                               <= GT1_RXOUTCLK_IN;
    gt2_txoutclk_i                               <= GT2_TXOUTCLK_IN;
    gt2_rxoutclk_i                               <= GT2_RXOUTCLK_IN;
    gt3_txoutclk_i                               <= GT3_TXOUTCLK_IN;
    gt3_rxoutclk_i                               <= GT3_RXOUTCLK_IN;
    gt4_txoutclk_i                               <= GT4_TXOUTCLK_IN;
    gt4_rxoutclk_i                               <= GT4_RXOUTCLK_IN;
    gt5_txoutclk_i                               <= GT5_TXOUTCLK_IN;
    gt5_rxoutclk_i                               <= GT5_RXOUTCLK_IN;
    gt6_txoutclk_i                               <= GT6_TXOUTCLK_IN;
    gt6_rxoutclk_i                               <= GT6_RXOUTCLK_IN;
    gt7_txoutclk_i                               <= GT7_TXOUTCLK_IN;
    gt7_rxoutclk_i                               <= GT7_RXOUTCLK_IN;
    gt8_txoutclk_i                               <= GT8_TXOUTCLK_IN;
    gt8_rxoutclk_i                               <= GT8_RXOUTCLK_IN;
    gt9_txoutclk_i                               <= GT9_TXOUTCLK_IN;
    gt9_rxoutclk_i                               <= GT9_RXOUTCLK_IN;
    gt10_txoutclk_i                              <= GT10_TXOUTCLK_IN;
    gt10_rxoutclk_i                              <= GT10_RXOUTCLK_IN;
    gt11_txoutclk_i                              <= GT11_TXOUTCLK_IN;
    gt11_rxoutclk_i                              <= GT11_RXOUTCLK_IN;
    gt12_txoutclk_i                              <= GT12_TXOUTCLK_IN;
    gt12_rxoutclk_i                              <= GT12_RXOUTCLK_IN;
    gt13_txoutclk_i                              <= GT13_TXOUTCLK_IN;
    gt13_rxoutclk_i                              <= GT13_RXOUTCLK_IN;
    gt14_txoutclk_i                              <= GT14_TXOUTCLK_IN;
    gt14_rxoutclk_i                              <= GT14_RXOUTCLK_IN;
    gt15_txoutclk_i                              <= GT15_TXOUTCLK_IN;
    gt15_rxoutclk_i                              <= GT15_RXOUTCLK_IN;
    gt16_txoutclk_i                              <= GT16_TXOUTCLK_IN;
    gt16_rxoutclk_i                              <= GT16_RXOUTCLK_IN;
    gt17_txoutclk_i                              <= GT17_TXOUTCLK_IN;
    gt17_rxoutclk_i                              <= GT17_RXOUTCLK_IN;
    gt18_txoutclk_i                              <= GT18_TXOUTCLK_IN;
    gt18_rxoutclk_i                              <= GT18_RXOUTCLK_IN;
    gt19_txoutclk_i                              <= GT19_TXOUTCLK_IN;
    gt19_rxoutclk_i                              <= GT19_RXOUTCLK_IN;
    gt20_txoutclk_i                              <= GT20_TXOUTCLK_IN;
    gt20_rxoutclk_i                              <= GT20_RXOUTCLK_IN;
    gt21_txoutclk_i                              <= GT21_TXOUTCLK_IN;
    gt21_rxoutclk_i                              <= GT21_RXOUTCLK_IN;
    gt22_txoutclk_i                              <= GT22_TXOUTCLK_IN;
    gt22_rxoutclk_i                              <= GT22_RXOUTCLK_IN;
    gt23_txoutclk_i                              <= GT23_TXOUTCLK_IN;
    gt23_rxoutclk_i                              <= GT23_RXOUTCLK_IN;
    gt24_txoutclk_i                              <= GT24_TXOUTCLK_IN;
    gt24_rxoutclk_i                              <= GT24_RXOUTCLK_IN;
    gt25_txoutclk_i                              <= GT25_TXOUTCLK_IN;
    gt25_rxoutclk_i                              <= GT25_RXOUTCLK_IN;
    gt26_txoutclk_i                              <= GT26_TXOUTCLK_IN;
    gt26_rxoutclk_i                              <= GT26_RXOUTCLK_IN;
    gt27_txoutclk_i                              <= GT27_TXOUTCLK_IN;
    gt27_rxoutclk_i                              <= GT27_RXOUTCLK_IN;
    gt28_txoutclk_i                              <= GT28_TXOUTCLK_IN;
    gt28_rxoutclk_i                              <= GT28_RXOUTCLK_IN;
    gt29_txoutclk_i                              <= GT29_TXOUTCLK_IN;
    gt29_rxoutclk_i                              <= GT29_RXOUTCLK_IN;
    gt30_txoutclk_i                              <= GT30_TXOUTCLK_IN;
    gt30_rxoutclk_i                              <= GT30_RXOUTCLK_IN;
    gt31_txoutclk_i                              <= GT31_TXOUTCLK_IN;
    gt31_rxoutclk_i                              <= GT31_RXOUTCLK_IN;

    Q2_CLK0_GTREFCLK_OUT                         <= q2_clk0_gtrefclk;
    Q5_CLK0_GTREFCLK_OUT                         <= q5_clk0_gtrefclk;
    Q7_CLK0_GTREFCLK_OUT                         <= q7_clk0_gtrefclk;

    --IBUFDS_GTE2
    ibufds_instq2_clk0 : IBUFDS_GTE2  
    port map
    (
        O               => 	q2_clk0_gtrefclk,
        ODIV2           =>    open,
        CEB             => 	tied_to_ground_i,
        I               => 	Q2_CLK0_GTREFCLK_PAD_P_IN,
        IB              => 	Q2_CLK0_GTREFCLK_PAD_N_IN
    );
    --IBUFDS_GTE2
    ibufds_instq5_clk0 : IBUFDS_GTE2  
    port map
    (
        O               => 	q5_clk0_gtrefclk,
        ODIV2           =>    open,
        CEB             => 	tied_to_ground_i,
        I               => 	Q5_CLK0_GTREFCLK_PAD_P_IN,
        IB              => 	Q5_CLK0_GTREFCLK_PAD_N_IN
    );
    --IBUFDS_GTE2
    ibufds_instq7_clk0 : IBUFDS_GTE2  
    port map
    (
        O               => 	q7_clk0_gtrefclk,
        ODIV2           =>    open,
        CEB             => 	tied_to_ground_i,
        I               => 	Q7_CLK0_GTREFCLK_PAD_P_IN,
        IB              => 	Q7_CLK0_GTREFCLK_PAD_N_IN
    );


    
    -- Instantiate a MMCM module to divide the reference clock. Uses internal feedback
    -- for improved jitter performance, and to avoid consuming an additional BUFG
    txoutclk_mmcm0_reset_i                       <= GT0_TX_MMCM_RESET_IN;
    -- txoutclk_mmcm0_i : gtwizard_0_CLOCK_MODULE
    -- generic map
    -- (
        -- MULT                            =>      10.0,
        -- DIVIDE                          =>      1,
        -- CLK_PERIOD                      =>      16.0,
        -- OUT0_DIVIDE                     =>      10.0,
        -- OUT1_DIVIDE                     =>      5,
        -- OUT2_DIVIDE                     =>      1,
        -- OUT3_DIVIDE                     =>      1
    -- )
    -- port map
    -- (
        -- CLK0_OUT                        =>      gt0_txusrclk2_i,
        -- CLK1_OUT                        =>      gt0_txusrclk_i,
        -- CLK2_OUT                        =>      open,
        -- CLK3_OUT                        =>      open,
        -- CLK_IN                          =>      gt0_txoutclk_i,
        -- MMCM_LOCKED_OUT                 =>      txoutclk_mmcm0_locked_i,
        -- MMCM_RESET_IN                   =>      txoutclk_mmcm0_reset_i
    -- );


    rxoutclk_mmcm1_reset_i                       <= GT0_RX_MMCM_RESET_IN;
    rxoutclk_mmcm1_i : gtwizard_0_CLOCK_MODULE
    generic map
    (
        MULT                            =>      5.0,
        DIVIDE                          =>      1,
        CLK_PERIOD                      =>      8.0,
        OUT0_DIVIDE                     =>      10.0,
        OUT1_DIVIDE                     =>      5,
        OUT2_DIVIDE                     =>      1,
        OUT3_DIVIDE                     =>      1
    )
    port map
    (
        CLK0_OUT                        =>      gt0_rxusrclk2_i,
        CLK1_OUT                        =>      gt0_rxusrclk_i,
        CLK2_OUT                        =>      open,
        CLK3_OUT                        =>      open,
        CLK_IN                          =>      gt0_rxoutclk_i,
        MMCM_LOCKED_OUT                 =>      rxoutclk_mmcm1_locked_i,
        MMCM_RESET_IN                   =>      rxoutclk_mmcm1_reset_i
    );


    txoutclk_mmcm2_reset_i                       <= GT12_TX_MMCM_RESET_IN;
    -- txoutclk_mmcm2_i : gtwizard_0_CLOCK_MODULE
    -- generic map
    -- (
        -- MULT                            =>      10.0,
        -- DIVIDE                          =>      1,
        -- CLK_PERIOD                      =>      16.0,
        -- OUT0_DIVIDE                     =>      10.0,
        -- OUT1_DIVIDE                     =>      5,
        -- OUT2_DIVIDE                     =>      1,
        -- OUT3_DIVIDE                     =>      1
    -- )
    -- port map
    -- (
        -- CLK0_OUT                        =>      gt12_txusrclk2_i,
        -- CLK1_OUT                        =>      gt12_txusrclk_i,
        -- CLK2_OUT                        =>      open,
        -- CLK3_OUT                        =>      open,
        -- CLK_IN                          =>      gt12_txoutclk_i,
        -- MMCM_LOCKED_OUT                 =>      txoutclk_mmcm2_locked_i,
        -- MMCM_RESET_IN                   =>      txoutclk_mmcm2_reset_i
    -- );


    rxoutclk_mmcm3_reset_i                       <= GT12_RX_MMCM_RESET_IN;
    rxoutclk_mmcm3_i : gtwizard_0_CLOCK_MODULE
    generic map
    (
        MULT                            =>      5.0,
        DIVIDE                          =>      1,
        CLK_PERIOD                      =>      8.0,
        OUT0_DIVIDE                     =>      10.0,
        OUT1_DIVIDE                     =>      5,
        OUT2_DIVIDE                     =>      1,
        OUT3_DIVIDE                     =>      1
    )
    port map
    (
        CLK0_OUT                        =>      gt12_rxusrclk2_i,
        CLK1_OUT                        =>      gt12_rxusrclk_i,
        CLK2_OUT                        =>      open,
        CLK3_OUT                        =>      open,
        CLK_IN                          =>      gt12_rxoutclk_i,
        MMCM_LOCKED_OUT                 =>      rxoutclk_mmcm3_locked_i,
        MMCM_RESET_IN                   =>      rxoutclk_mmcm3_reset_i
    );


    txoutclk_mmcm4_reset_i                       <= GT24_TX_MMCM_RESET_IN;
    -- txoutclk_mmcm4_i : gtwizard_0_CLOCK_MODULE
    -- generic map
    -- (
        -- MULT                            =>      10.0,
        -- DIVIDE                          =>      1,
        -- CLK_PERIOD                      =>      16.0,
        -- OUT0_DIVIDE                     =>      10.0,
        -- OUT1_DIVIDE                     =>      5,
        -- OUT2_DIVIDE                     =>      1,
        -- OUT3_DIVIDE                     =>      1
    -- )
    -- port map
    -- (
        -- CLK0_OUT                        =>      gt24_txusrclk2_i,
        -- CLK1_OUT                        =>      gt24_txusrclk_i,
        -- CLK2_OUT                        =>      open,
        -- CLK3_OUT                        =>      open,
        -- CLK_IN                          =>      gt24_txoutclk_i,
        -- MMCM_LOCKED_OUT                 =>      txoutclk_mmcm4_locked_i,
        -- MMCM_RESET_IN                   =>      txoutclk_mmcm4_reset_i
    -- );


    rxoutclk_mmcm5_reset_i                       <= GT24_RX_MMCM_RESET_IN;
    rxoutclk_mmcm5_i : gtwizard_0_CLOCK_MODULE
    generic map
    (
        MULT                            =>      5.0,
        DIVIDE                          =>      1,
        CLK_PERIOD                      =>      8.0,
        OUT0_DIVIDE                     =>      10.0,
        OUT1_DIVIDE                     =>      5,
        OUT2_DIVIDE                     =>      1,
        OUT3_DIVIDE                     =>      1
    )
    port map
    (
        CLK0_OUT                        =>      gt24_rxusrclk2_i,
        CLK1_OUT                        =>      gt24_rxusrclk_i,
        CLK2_OUT                        =>      open,
        CLK3_OUT                        =>      open,
        CLK_IN                          =>      gt24_rxoutclk_i,
        MMCM_LOCKED_OUT                 =>      rxoutclk_mmcm5_locked_i,
        MMCM_RESET_IN                   =>      rxoutclk_mmcm5_reset_i
    );



 
GT0_TXUSRCLK_OUT                             <= txusrclk_in;
GT0_TXUSRCLK2_OUT                            <= txusrclk2_in;
GT0_TXCLK_LOCK_OUT                           <= '1';
GT0_RXUSRCLK_OUT                             <= gt0_rxusrclk_i;
GT0_RXUSRCLK2_OUT                            <= gt0_rxusrclk2_i;
GT0_RXCLK_LOCK_OUT                           <= rxoutclk_mmcm1_locked_i;
 
GT1_TXUSRCLK_OUT                             <= txusrclk_in;
GT1_TXUSRCLK2_OUT                            <= txusrclk2_in;
GT1_TXCLK_LOCK_OUT                           <= '1';
GT1_RXUSRCLK_OUT                             <= gt0_rxusrclk_i;
GT1_RXUSRCLK2_OUT                            <= gt0_rxusrclk2_i;
GT1_RXCLK_LOCK_OUT                           <= rxoutclk_mmcm1_locked_i;
 
GT2_TXUSRCLK_OUT                             <= txusrclk_in;
GT2_TXUSRCLK2_OUT                            <= txusrclk2_in;
GT2_TXCLK_LOCK_OUT                           <= '1';
GT2_RXUSRCLK_OUT                             <= gt0_rxusrclk_i;
GT2_RXUSRCLK2_OUT                            <= gt0_rxusrclk2_i;
GT2_RXCLK_LOCK_OUT                           <= rxoutclk_mmcm1_locked_i;
 
GT3_TXUSRCLK_OUT                             <= txusrclk_in;
GT3_TXUSRCLK2_OUT                            <= txusrclk2_in;
GT3_TXCLK_LOCK_OUT                           <= '1';
GT3_RXUSRCLK_OUT                             <= gt0_rxusrclk_i;
GT3_RXUSRCLK2_OUT                            <= gt0_rxusrclk2_i;
GT3_RXCLK_LOCK_OUT                           <= rxoutclk_mmcm1_locked_i;
 
GT4_TXUSRCLK_OUT                             <= txusrclk_in;
GT4_TXUSRCLK2_OUT                            <= txusrclk2_in;
GT4_TXCLK_LOCK_OUT                           <= '1';
GT4_RXUSRCLK_OUT                             <= gt0_rxusrclk_i;
GT4_RXUSRCLK2_OUT                            <= gt0_rxusrclk2_i;
GT4_RXCLK_LOCK_OUT                           <= rxoutclk_mmcm1_locked_i;
 
GT5_TXUSRCLK_OUT                             <= txusrclk_in;
GT5_TXUSRCLK2_OUT                            <= txusrclk2_in;
GT5_TXCLK_LOCK_OUT                           <= '1';
GT5_RXUSRCLK_OUT                             <= gt0_rxusrclk_i;
GT5_RXUSRCLK2_OUT                            <= gt0_rxusrclk2_i;
GT5_RXCLK_LOCK_OUT                           <= rxoutclk_mmcm1_locked_i;
 
GT6_TXUSRCLK_OUT                             <= txusrclk_in;
GT6_TXUSRCLK2_OUT                            <= txusrclk2_in;
GT6_TXCLK_LOCK_OUT                           <= '1';
GT6_RXUSRCLK_OUT                             <= gt0_rxusrclk_i;
GT6_RXUSRCLK2_OUT                            <= gt0_rxusrclk2_i;
GT6_RXCLK_LOCK_OUT                           <= rxoutclk_mmcm1_locked_i;
 
GT7_TXUSRCLK_OUT                             <= txusrclk_in;
GT7_TXUSRCLK2_OUT                            <= txusrclk2_in;
GT7_TXCLK_LOCK_OUT                           <= '1';
GT7_RXUSRCLK_OUT                             <= gt0_rxusrclk_i;
GT7_RXUSRCLK2_OUT                            <= gt0_rxusrclk2_i;
GT7_RXCLK_LOCK_OUT                           <= rxoutclk_mmcm1_locked_i;
 
GT8_TXUSRCLK_OUT                             <= txusrclk_in;
GT8_TXUSRCLK2_OUT                            <= txusrclk2_in;
GT8_TXCLK_LOCK_OUT                           <= '1';
GT8_RXUSRCLK_OUT                             <= gt0_rxusrclk_i;
GT8_RXUSRCLK2_OUT                            <= gt0_rxusrclk2_i;
GT8_RXCLK_LOCK_OUT                           <= rxoutclk_mmcm1_locked_i;
 
GT9_TXUSRCLK_OUT                             <= txusrclk_in;
GT9_TXUSRCLK2_OUT                            <= txusrclk2_in;
GT9_TXCLK_LOCK_OUT                           <= '1';
GT9_RXUSRCLK_OUT                             <= gt0_rxusrclk_i;
GT9_RXUSRCLK2_OUT                            <= gt0_rxusrclk2_i;
GT9_RXCLK_LOCK_OUT                           <= rxoutclk_mmcm1_locked_i;
 
GT10_TXUSRCLK_OUT                            <= txusrclk_in;
GT10_TXUSRCLK2_OUT                           <= txusrclk2_in;
GT10_TXCLK_LOCK_OUT                          <= '1';
GT10_RXUSRCLK_OUT                            <= gt0_rxusrclk_i;
GT10_RXUSRCLK2_OUT                           <= gt0_rxusrclk2_i;
GT10_RXCLK_LOCK_OUT                          <= rxoutclk_mmcm1_locked_i;
 
GT11_TXUSRCLK_OUT                            <= txusrclk_in;
GT11_TXUSRCLK2_OUT                           <= txusrclk2_in;
GT11_TXCLK_LOCK_OUT                          <= '1';
GT11_RXUSRCLK_OUT                            <= gt0_rxusrclk_i;
GT11_RXUSRCLK2_OUT                           <= gt0_rxusrclk2_i;
GT11_RXCLK_LOCK_OUT                          <= rxoutclk_mmcm1_locked_i;
 
GT12_TXUSRCLK_OUT                            <= txusrclk_in;
GT12_TXUSRCLK2_OUT                           <= txusrclk2_in;
GT12_TXCLK_LOCK_OUT                          <= '1';
GT12_RXUSRCLK_OUT                            <= gt0_rxusrclk_i;
GT12_RXUSRCLK2_OUT                           <= gt0_rxusrclk2_i;
GT12_RXCLK_LOCK_OUT                          <= rxoutclk_mmcm1_locked_i;
 
GT13_TXUSRCLK_OUT                            <= txusrclk_in;
GT13_TXUSRCLK2_OUT                           <= txusrclk2_in;
GT13_TXCLK_LOCK_OUT                          <= '1';
GT13_RXUSRCLK_OUT                            <= gt0_rxusrclk_i;
GT13_RXUSRCLK2_OUT                           <= gt0_rxusrclk2_i;
GT13_RXCLK_LOCK_OUT                          <= rxoutclk_mmcm1_locked_i;
 
GT14_TXUSRCLK_OUT                            <= txusrclk_in;
GT14_TXUSRCLK2_OUT                           <= txusrclk2_in;
GT14_TXCLK_LOCK_OUT                          <= '1';
GT14_RXUSRCLK_OUT                            <= gt0_rxusrclk_i;
GT14_RXUSRCLK2_OUT                           <= gt0_rxusrclk2_i;
GT14_RXCLK_LOCK_OUT                          <= rxoutclk_mmcm1_locked_i;
 
GT15_TXUSRCLK_OUT                            <= txusrclk_in;
GT15_TXUSRCLK2_OUT                           <= txusrclk2_in;
GT15_TXCLK_LOCK_OUT                          <= '1';
GT15_RXUSRCLK_OUT                            <= gt0_rxusrclk_i;
GT15_RXUSRCLK2_OUT                           <= gt0_rxusrclk2_i;
GT15_RXCLK_LOCK_OUT                          <= rxoutclk_mmcm1_locked_i;
 
GT16_TXUSRCLK_OUT                            <= txusrclk_in;
GT16_TXUSRCLK2_OUT                           <= txusrclk2_in;
GT16_TXCLK_LOCK_OUT                          <= '1';
GT16_RXUSRCLK_OUT                            <= gt0_rxusrclk_i;
GT16_RXUSRCLK2_OUT                           <= gt0_rxusrclk2_i;
GT16_RXCLK_LOCK_OUT                          <= rxoutclk_mmcm1_locked_i;
 
GT17_TXUSRCLK_OUT                            <= txusrclk_in;
GT17_TXUSRCLK2_OUT                           <= txusrclk2_in;
GT17_TXCLK_LOCK_OUT                          <= '1';
GT17_RXUSRCLK_OUT                            <= gt0_rxusrclk_i;
GT17_RXUSRCLK2_OUT                           <= gt0_rxusrclk2_i;
GT17_RXCLK_LOCK_OUT                          <= rxoutclk_mmcm1_locked_i;
 
GT18_TXUSRCLK_OUT                            <= txusrclk_in;
GT18_TXUSRCLK2_OUT                           <= txusrclk2_in;
GT18_TXCLK_LOCK_OUT                          <= '1';
GT18_RXUSRCLK_OUT                            <= gt0_rxusrclk_i;
GT18_RXUSRCLK2_OUT                           <= gt0_rxusrclk2_i;
GT18_RXCLK_LOCK_OUT                          <= rxoutclk_mmcm1_locked_i;
 
GT19_TXUSRCLK_OUT                            <= txusrclk_in;
GT19_TXUSRCLK2_OUT                           <= txusrclk2_in;
GT19_TXCLK_LOCK_OUT                          <= '1';
GT19_RXUSRCLK_OUT                            <= gt0_rxusrclk_i;
GT19_RXUSRCLK2_OUT                           <= gt0_rxusrclk2_i;
GT19_RXCLK_LOCK_OUT                          <= rxoutclk_mmcm1_locked_i;
 
GT20_TXUSRCLK_OUT                            <= txusrclk_in;
GT20_TXUSRCLK2_OUT                           <= txusrclk2_in;
GT20_TXCLK_LOCK_OUT                          <= '1';
GT20_RXUSRCLK_OUT                            <= gt0_rxusrclk_i;
GT20_RXUSRCLK2_OUT                           <= gt0_rxusrclk2_i;
GT20_RXCLK_LOCK_OUT                          <= rxoutclk_mmcm1_locked_i;
 
GT21_TXUSRCLK_OUT                            <= txusrclk_in;
GT21_TXUSRCLK2_OUT                           <= txusrclk2_in;
GT21_TXCLK_LOCK_OUT                          <= '1';
GT21_RXUSRCLK_OUT                            <= gt0_rxusrclk_i;
GT21_RXUSRCLK2_OUT                           <= gt0_rxusrclk2_i;
GT21_RXCLK_LOCK_OUT                          <= rxoutclk_mmcm1_locked_i;
 
GT22_TXUSRCLK_OUT                            <= txusrclk_in;
GT22_TXUSRCLK2_OUT                           <= txusrclk2_in;
GT22_TXCLK_LOCK_OUT                          <= '1';
GT22_RXUSRCLK_OUT                            <= gt0_rxusrclk_i;
GT22_RXUSRCLK2_OUT                           <= gt0_rxusrclk2_i;
GT22_RXCLK_LOCK_OUT                          <= rxoutclk_mmcm1_locked_i;
 
GT23_TXUSRCLK_OUT                            <= txusrclk_in;
GT23_TXUSRCLK2_OUT                           <= txusrclk2_in;
GT23_TXCLK_LOCK_OUT                          <= '1';
GT23_RXUSRCLK_OUT                            <= gt0_rxusrclk_i;
GT23_RXUSRCLK2_OUT                           <= gt0_rxusrclk2_i;
GT23_RXCLK_LOCK_OUT                          <= rxoutclk_mmcm1_locked_i;
 
GT24_TXUSRCLK_OUT                            <= txusrclk_in;
GT24_TXUSRCLK2_OUT                           <= txusrclk2_in;
GT24_TXCLK_LOCK_OUT                          <= '1';
GT24_RXUSRCLK_OUT                            <= gt0_rxusrclk_i;
GT24_RXUSRCLK2_OUT                           <= gt0_rxusrclk2_i;
GT24_RXCLK_LOCK_OUT                          <= rxoutclk_mmcm1_locked_i;
 
GT25_TXUSRCLK_OUT                            <= txusrclk_in;
GT25_TXUSRCLK2_OUT                           <= txusrclk2_in;
GT25_TXCLK_LOCK_OUT                          <= '1';
GT25_RXUSRCLK_OUT                            <= gt0_rxusrclk_i;
GT25_RXUSRCLK2_OUT                           <= gt0_rxusrclk2_i;
GT25_RXCLK_LOCK_OUT                          <= rxoutclk_mmcm1_locked_i;
 
GT26_TXUSRCLK_OUT                            <= txusrclk_in;
GT26_TXUSRCLK2_OUT                           <= txusrclk2_in;
GT26_TXCLK_LOCK_OUT                          <= '1';
GT26_RXUSRCLK_OUT                            <= gt0_rxusrclk_i;
GT26_RXUSRCLK2_OUT                           <= gt0_rxusrclk2_i;
GT26_RXCLK_LOCK_OUT                          <= rxoutclk_mmcm1_locked_i;
 
GT27_TXUSRCLK_OUT                            <= txusrclk_in;
GT27_TXUSRCLK2_OUT                           <= txusrclk2_in;
GT27_TXCLK_LOCK_OUT                          <= '1';
GT27_RXUSRCLK_OUT                            <= gt0_rxusrclk_i;
GT27_RXUSRCLK2_OUT                           <= gt0_rxusrclk2_i;
GT27_RXCLK_LOCK_OUT                          <= rxoutclk_mmcm1_locked_i;
 
GT28_TXUSRCLK_OUT                            <= txusrclk_in;
GT28_TXUSRCLK2_OUT                           <= txusrclk2_in;
GT28_TXCLK_LOCK_OUT                          <= '1';
GT28_RXUSRCLK_OUT                            <= gt0_rxusrclk_i;
GT28_RXUSRCLK2_OUT                           <= gt0_rxusrclk2_i;
GT28_RXCLK_LOCK_OUT                          <= rxoutclk_mmcm1_locked_i;
 
GT29_TXUSRCLK_OUT                            <= txusrclk_in;
GT29_TXUSRCLK2_OUT                           <= txusrclk2_in;
GT29_TXCLK_LOCK_OUT                          <= '1';
GT29_RXUSRCLK_OUT                            <= gt0_rxusrclk_i;
GT29_RXUSRCLK2_OUT                           <= gt0_rxusrclk2_i;
GT29_RXCLK_LOCK_OUT                          <= rxoutclk_mmcm1_locked_i;
 
GT30_TXUSRCLK_OUT                            <= txusrclk_in;
GT30_TXUSRCLK2_OUT                           <= txusrclk2_in;
GT30_TXCLK_LOCK_OUT                          <= '1';
GT30_RXUSRCLK_OUT                            <= gt0_rxusrclk_i;
GT30_RXUSRCLK2_OUT                           <= gt0_rxusrclk2_i;
GT30_RXCLK_LOCK_OUT                          <= rxoutclk_mmcm1_locked_i;
 
GT31_TXUSRCLK_OUT                            <= txusrclk_in;
GT31_TXUSRCLK2_OUT                           <= txusrclk2_in;
GT31_TXCLK_LOCK_OUT                          <= '1';
GT31_RXUSRCLK_OUT                            <= gt0_rxusrclk_i;
GT31_RXUSRCLK2_OUT                           <= gt0_rxusrclk2_i;
GT31_RXCLK_LOCK_OUT                          <= rxoutclk_mmcm1_locked_i;
end RTL;

