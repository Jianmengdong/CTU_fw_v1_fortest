------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 3.6
--  \   \         Application : 7 Series FPGAs Transceivers Wizard 
--  /   /         Filename : gtwizard_0_init.vhd
-- /___/   /\      
-- \   \  /  \ 
--  \___\/\___\
--
--  Description : This module instantiates the modules required for
--                reset and initialisation of the Transceiver
--
-- Module gtwizard_0_init
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;

--***********************************Entity Declaration************************

entity gtwizard_0_init is
generic
(
    EXAMPLE_SIM_GTRESET_SPEEDUP             : string    := "FALSE";     -- simulation setting for GT SecureIP model
    EXAMPLE_SIMULATION                      : integer   := 0;          -- Set to 1 for simulation
 
 
    STABLE_CLOCK_PERIOD                     : integer   := 8;  
        -- Set to 1 for simulation
    EXAMPLE_USE_CHIPSCOPE                   : integer   := 0           -- Set to 1 to use Chipscope to drive resets

);
port
(
    SYSCLK_IN                               : in   std_logic;
    SOFT_RESET_TX_IN                        : in   std_logic;
    SOFT_RESET_RX_IN                        : in   std_logic;
    DONT_RESET_ON_DATA_ERROR_IN             : in   std_logic;
    GT0_DRP_BUSY_OUT                        : out  std_logic;
    GT0_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_DATA_VALID_IN                       : in   std_logic;
    GT0_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT0_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT0_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT0_RX_MMCM_RESET_OUT                   : out  std_logic;
    GT1_DRP_BUSY_OUT                        : out  std_logic;
    GT1_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT1_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT1_DATA_VALID_IN                       : in   std_logic;
    GT1_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT1_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT1_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT1_RX_MMCM_RESET_OUT                   : out  std_logic;
    GT2_DRP_BUSY_OUT                        : out  std_logic;
    GT2_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT2_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT2_DATA_VALID_IN                       : in   std_logic;
    GT2_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT2_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT2_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT2_RX_MMCM_RESET_OUT                   : out  std_logic;
    GT3_DRP_BUSY_OUT                        : out  std_logic;
    GT3_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT3_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT3_DATA_VALID_IN                       : in   std_logic;
    GT3_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT3_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT3_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT3_RX_MMCM_RESET_OUT                   : out  std_logic;
    GT4_DRP_BUSY_OUT                        : out  std_logic;
    GT4_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT4_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT4_DATA_VALID_IN                       : in   std_logic;
    GT4_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT4_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT4_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT4_RX_MMCM_RESET_OUT                   : out  std_logic;
    GT5_DRP_BUSY_OUT                        : out  std_logic;
    GT5_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT5_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT5_DATA_VALID_IN                       : in   std_logic;
    GT5_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT5_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT5_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT5_RX_MMCM_RESET_OUT                   : out  std_logic;
    GT6_DRP_BUSY_OUT                        : out  std_logic;
    GT6_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT6_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT6_DATA_VALID_IN                       : in   std_logic;
    GT6_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT6_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT6_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT6_RX_MMCM_RESET_OUT                   : out  std_logic;
    GT7_DRP_BUSY_OUT                        : out  std_logic;
    GT7_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT7_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT7_DATA_VALID_IN                       : in   std_logic;
    GT7_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT7_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT7_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT7_RX_MMCM_RESET_OUT                   : out  std_logic;
    GT8_DRP_BUSY_OUT                        : out  std_logic;
    GT8_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT8_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT8_DATA_VALID_IN                       : in   std_logic;
    GT8_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT8_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT8_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT8_RX_MMCM_RESET_OUT                   : out  std_logic;
    GT9_DRP_BUSY_OUT                        : out  std_logic;
    GT9_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT9_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT9_DATA_VALID_IN                       : in   std_logic;
    GT9_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT9_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT9_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT9_RX_MMCM_RESET_OUT                   : out  std_logic;
    GT10_DRP_BUSY_OUT                       : out  std_logic;
    GT10_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT10_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT10_DATA_VALID_IN                      : in   std_logic;
    GT10_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT10_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT10_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT10_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT11_DRP_BUSY_OUT                       : out  std_logic;
    GT11_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT11_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT11_DATA_VALID_IN                      : in   std_logic;
    GT11_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT11_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT11_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT11_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT12_DRP_BUSY_OUT                       : out  std_logic;
    GT12_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT12_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT12_DATA_VALID_IN                      : in   std_logic;
    GT12_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT12_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT12_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT12_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT13_DRP_BUSY_OUT                       : out  std_logic;
    GT13_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT13_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT13_DATA_VALID_IN                      : in   std_logic;
    GT13_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT13_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT13_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT13_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT14_DRP_BUSY_OUT                       : out  std_logic;
    GT14_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT14_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT14_DATA_VALID_IN                      : in   std_logic;
    GT14_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT14_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT14_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT14_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT15_DRP_BUSY_OUT                       : out  std_logic;
    GT15_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT15_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT15_DATA_VALID_IN                      : in   std_logic;
    GT15_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT15_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT15_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT15_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT16_DRP_BUSY_OUT                       : out  std_logic;
    GT16_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT16_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT16_DATA_VALID_IN                      : in   std_logic;
    GT16_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT16_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT16_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT16_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT17_DRP_BUSY_OUT                       : out  std_logic;
    GT17_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT17_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT17_DATA_VALID_IN                      : in   std_logic;
    GT17_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT17_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT17_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT17_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT18_DRP_BUSY_OUT                       : out  std_logic;
    GT18_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT18_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT18_DATA_VALID_IN                      : in   std_logic;
    GT18_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT18_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT18_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT18_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT19_DRP_BUSY_OUT                       : out  std_logic;
    GT19_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT19_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT19_DATA_VALID_IN                      : in   std_logic;
    GT19_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT19_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT19_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT19_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT20_DRP_BUSY_OUT                       : out  std_logic;
    GT20_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT20_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT20_DATA_VALID_IN                      : in   std_logic;
    GT20_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT20_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT20_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT20_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT21_DRP_BUSY_OUT                       : out  std_logic;
    GT21_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT21_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT21_DATA_VALID_IN                      : in   std_logic;
    GT21_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT21_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT21_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT21_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT22_DRP_BUSY_OUT                       : out  std_logic;
    GT22_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT22_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT22_DATA_VALID_IN                      : in   std_logic;
    GT22_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT22_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT22_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT22_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT23_DRP_BUSY_OUT                       : out  std_logic;
    GT23_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT23_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT23_DATA_VALID_IN                      : in   std_logic;
    GT23_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT23_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT23_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT23_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT24_DRP_BUSY_OUT                       : out  std_logic;
    GT24_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT24_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT24_DATA_VALID_IN                      : in   std_logic;
    GT24_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT24_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT24_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT24_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT25_DRP_BUSY_OUT                       : out  std_logic;
    GT25_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT25_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT25_DATA_VALID_IN                      : in   std_logic;
    GT25_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT25_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT25_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT25_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT26_DRP_BUSY_OUT                       : out  std_logic;
    GT26_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT26_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT26_DATA_VALID_IN                      : in   std_logic;
    GT26_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT26_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT26_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT26_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT27_DRP_BUSY_OUT                       : out  std_logic;
    GT27_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT27_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT27_DATA_VALID_IN                      : in   std_logic;
    GT27_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT27_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT27_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT27_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT28_DRP_BUSY_OUT                       : out  std_logic;
    GT28_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT28_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT28_DATA_VALID_IN                      : in   std_logic;
    GT28_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT28_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT28_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT28_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT29_DRP_BUSY_OUT                       : out  std_logic;
    GT29_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT29_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT29_DATA_VALID_IN                      : in   std_logic;
    GT29_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT29_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT29_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT29_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT30_DRP_BUSY_OUT                       : out  std_logic;
    GT30_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT30_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT30_DATA_VALID_IN                      : in   std_logic;
    GT30_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT30_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT30_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT30_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT31_DRP_BUSY_OUT                       : out  std_logic;
    GT31_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT31_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT31_DATA_VALID_IN                      : in   std_logic;
    GT31_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT31_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT31_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT31_RX_MMCM_RESET_OUT                  : out  std_logic;
    --_________________________________________________________________________
    --GT0  (X1Y4)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt0_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt0_drpclk_in                           : in   std_logic;
    gt0_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt0_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt0_drpen_in                            : in   std_logic;
    gt0_drprdy_out                          : out  std_logic;
    gt0_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt0_eyescanreset_in                     : in   std_logic;
    gt0_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt0_eyescandataerror_out                : out  std_logic;
    gt0_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt0_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt0_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt0_rxusrclk_in                         : in   std_logic;
    gt0_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt0_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt0_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt0_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt0_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt0_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt0_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt0_rxbyteisaligned_out                 : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt0_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt0_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt0_rxoutclk_out                        : out  std_logic;
    gt0_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt0_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt0_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt0_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt0_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt0_gttxreset_in                        : in   std_logic;
    gt0_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt0_txusrclk_in                         : in   std_logic;
    gt0_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt0_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt0_gthtxn_out                          : out  std_logic;
    gt0_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt0_txoutclk_out                        : out  std_logic;
    gt0_txoutclkfabric_out                  : out  std_logic;
    gt0_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt0_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt0_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT1  (X1Y5)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt1_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt1_drpclk_in                           : in   std_logic;
    gt1_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt1_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt1_drpen_in                            : in   std_logic;
    gt1_drprdy_out                          : out  std_logic;
    gt1_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt1_eyescanreset_in                     : in   std_logic;
    gt1_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt1_eyescandataerror_out                : out  std_logic;
    gt1_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt1_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt1_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt1_rxusrclk_in                         : in   std_logic;
    gt1_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt1_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt1_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt1_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt1_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt1_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt1_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt1_rxbyteisaligned_out                 : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt1_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt1_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt1_rxoutclk_out                        : out  std_logic;
    gt1_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt1_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt1_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt1_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt1_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt1_gttxreset_in                        : in   std_logic;
    gt1_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt1_txusrclk_in                         : in   std_logic;
    gt1_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt1_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt1_gthtxn_out                          : out  std_logic;
    gt1_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt1_txoutclk_out                        : out  std_logic;
    gt1_txoutclkfabric_out                  : out  std_logic;
    gt1_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt1_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt1_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT2  (X1Y6)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt2_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt2_drpclk_in                           : in   std_logic;
    gt2_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt2_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt2_drpen_in                            : in   std_logic;
    gt2_drprdy_out                          : out  std_logic;
    gt2_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt2_eyescanreset_in                     : in   std_logic;
    gt2_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt2_eyescandataerror_out                : out  std_logic;
    gt2_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt2_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt2_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt2_rxusrclk_in                         : in   std_logic;
    gt2_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt2_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt2_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt2_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt2_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt2_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt2_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt2_rxbyteisaligned_out                 : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt2_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt2_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt2_rxoutclk_out                        : out  std_logic;
    gt2_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt2_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt2_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt2_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt2_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt2_gttxreset_in                        : in   std_logic;
    gt2_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt2_txusrclk_in                         : in   std_logic;
    gt2_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt2_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt2_gthtxn_out                          : out  std_logic;
    gt2_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt2_txoutclk_out                        : out  std_logic;
    gt2_txoutclkfabric_out                  : out  std_logic;
    gt2_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt2_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt2_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT3  (X1Y7)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt3_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt3_drpclk_in                           : in   std_logic;
    gt3_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt3_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt3_drpen_in                            : in   std_logic;
    gt3_drprdy_out                          : out  std_logic;
    gt3_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt3_eyescanreset_in                     : in   std_logic;
    gt3_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt3_eyescandataerror_out                : out  std_logic;
    gt3_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt3_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt3_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt3_rxusrclk_in                         : in   std_logic;
    gt3_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt3_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt3_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt3_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt3_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt3_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt3_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt3_rxbyteisaligned_out                 : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt3_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt3_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt3_rxoutclk_out                        : out  std_logic;
    gt3_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt3_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt3_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt3_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt3_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt3_gttxreset_in                        : in   std_logic;
    gt3_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt3_txusrclk_in                         : in   std_logic;
    gt3_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt3_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt3_gthtxn_out                          : out  std_logic;
    gt3_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt3_txoutclk_out                        : out  std_logic;
    gt3_txoutclkfabric_out                  : out  std_logic;
    gt3_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt3_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt3_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT4  (X1Y8)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt4_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt4_drpclk_in                           : in   std_logic;
    gt4_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt4_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt4_drpen_in                            : in   std_logic;
    gt4_drprdy_out                          : out  std_logic;
    gt4_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt4_eyescanreset_in                     : in   std_logic;
    gt4_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt4_eyescandataerror_out                : out  std_logic;
    gt4_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt4_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt4_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt4_rxusrclk_in                         : in   std_logic;
    gt4_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt4_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt4_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt4_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt4_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt4_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt4_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt4_rxbyteisaligned_out                 : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt4_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt4_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt4_rxoutclk_out                        : out  std_logic;
    gt4_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt4_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt4_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt4_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt4_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt4_gttxreset_in                        : in   std_logic;
    gt4_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt4_txusrclk_in                         : in   std_logic;
    gt4_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt4_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt4_gthtxn_out                          : out  std_logic;
    gt4_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt4_txoutclk_out                        : out  std_logic;
    gt4_txoutclkfabric_out                  : out  std_logic;
    gt4_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt4_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt4_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT5  (X1Y9)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt5_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt5_drpclk_in                           : in   std_logic;
    gt5_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt5_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt5_drpen_in                            : in   std_logic;
    gt5_drprdy_out                          : out  std_logic;
    gt5_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt5_eyescanreset_in                     : in   std_logic;
    gt5_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt5_eyescandataerror_out                : out  std_logic;
    gt5_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt5_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt5_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt5_rxusrclk_in                         : in   std_logic;
    gt5_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt5_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt5_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt5_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt5_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt5_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt5_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt5_rxbyteisaligned_out                 : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt5_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt5_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt5_rxoutclk_out                        : out  std_logic;
    gt5_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt5_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt5_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt5_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt5_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt5_gttxreset_in                        : in   std_logic;
    gt5_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt5_txusrclk_in                         : in   std_logic;
    gt5_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt5_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt5_gthtxn_out                          : out  std_logic;
    gt5_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt5_txoutclk_out                        : out  std_logic;
    gt5_txoutclkfabric_out                  : out  std_logic;
    gt5_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt5_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt5_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT6  (X1Y10)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt6_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt6_drpclk_in                           : in   std_logic;
    gt6_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt6_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt6_drpen_in                            : in   std_logic;
    gt6_drprdy_out                          : out  std_logic;
    gt6_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt6_eyescanreset_in                     : in   std_logic;
    gt6_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt6_eyescandataerror_out                : out  std_logic;
    gt6_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt6_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt6_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt6_rxusrclk_in                         : in   std_logic;
    gt6_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt6_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt6_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt6_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt6_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt6_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt6_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt6_rxbyteisaligned_out                 : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt6_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt6_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt6_rxoutclk_out                        : out  std_logic;
    gt6_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt6_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt6_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt6_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt6_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt6_gttxreset_in                        : in   std_logic;
    gt6_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt6_txusrclk_in                         : in   std_logic;
    gt6_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt6_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt6_gthtxn_out                          : out  std_logic;
    gt6_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt6_txoutclk_out                        : out  std_logic;
    gt6_txoutclkfabric_out                  : out  std_logic;
    gt6_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt6_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt6_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT7  (X1Y11)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt7_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt7_drpclk_in                           : in   std_logic;
    gt7_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt7_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt7_drpen_in                            : in   std_logic;
    gt7_drprdy_out                          : out  std_logic;
    gt7_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt7_eyescanreset_in                     : in   std_logic;
    gt7_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt7_eyescandataerror_out                : out  std_logic;
    gt7_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt7_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt7_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt7_rxusrclk_in                         : in   std_logic;
    gt7_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt7_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt7_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt7_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt7_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt7_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt7_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt7_rxbyteisaligned_out                 : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt7_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt7_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt7_rxoutclk_out                        : out  std_logic;
    gt7_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt7_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt7_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt7_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt7_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt7_gttxreset_in                        : in   std_logic;
    gt7_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt7_txusrclk_in                         : in   std_logic;
    gt7_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt7_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt7_gthtxn_out                          : out  std_logic;
    gt7_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt7_txoutclk_out                        : out  std_logic;
    gt7_txoutclkfabric_out                  : out  std_logic;
    gt7_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt7_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt7_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT8  (X1Y12)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt8_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt8_drpclk_in                           : in   std_logic;
    gt8_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt8_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt8_drpen_in                            : in   std_logic;
    gt8_drprdy_out                          : out  std_logic;
    gt8_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt8_eyescanreset_in                     : in   std_logic;
    gt8_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt8_eyescandataerror_out                : out  std_logic;
    gt8_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt8_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt8_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt8_rxusrclk_in                         : in   std_logic;
    gt8_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt8_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt8_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt8_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt8_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt8_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt8_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt8_rxbyteisaligned_out                 : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt8_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt8_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt8_rxoutclk_out                        : out  std_logic;
    gt8_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt8_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt8_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt8_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt8_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt8_gttxreset_in                        : in   std_logic;
    gt8_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt8_txusrclk_in                         : in   std_logic;
    gt8_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt8_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt8_gthtxn_out                          : out  std_logic;
    gt8_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt8_txoutclk_out                        : out  std_logic;
    gt8_txoutclkfabric_out                  : out  std_logic;
    gt8_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt8_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt8_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT9  (X1Y13)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt9_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt9_drpclk_in                           : in   std_logic;
    gt9_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt9_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt9_drpen_in                            : in   std_logic;
    gt9_drprdy_out                          : out  std_logic;
    gt9_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt9_eyescanreset_in                     : in   std_logic;
    gt9_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt9_eyescandataerror_out                : out  std_logic;
    gt9_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt9_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt9_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt9_rxusrclk_in                         : in   std_logic;
    gt9_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt9_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt9_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt9_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt9_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt9_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt9_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt9_rxbyteisaligned_out                 : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt9_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt9_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt9_rxoutclk_out                        : out  std_logic;
    gt9_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt9_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt9_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt9_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt9_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt9_gttxreset_in                        : in   std_logic;
    gt9_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt9_txusrclk_in                         : in   std_logic;
    gt9_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt9_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt9_gthtxn_out                          : out  std_logic;
    gt9_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt9_txoutclk_out                        : out  std_logic;
    gt9_txoutclkfabric_out                  : out  std_logic;
    gt9_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt9_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt9_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT10  (X1Y14)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt10_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt10_drpclk_in                          : in   std_logic;
    gt10_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt10_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt10_drpen_in                           : in   std_logic;
    gt10_drprdy_out                         : out  std_logic;
    gt10_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt10_eyescanreset_in                    : in   std_logic;
    gt10_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt10_eyescandataerror_out               : out  std_logic;
    gt10_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt10_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt10_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt10_rxusrclk_in                        : in   std_logic;
    gt10_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt10_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt10_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt10_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt10_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt10_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt10_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt10_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt10_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt10_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt10_rxoutclk_out                       : out  std_logic;
    gt10_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt10_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt10_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt10_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt10_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt10_gttxreset_in                       : in   std_logic;
    gt10_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt10_txusrclk_in                        : in   std_logic;
    gt10_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt10_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt10_gthtxn_out                         : out  std_logic;
    gt10_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt10_txoutclk_out                       : out  std_logic;
    gt10_txoutclkfabric_out                 : out  std_logic;
    gt10_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt10_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt10_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT11  (X1Y15)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt11_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt11_drpclk_in                          : in   std_logic;
    gt11_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt11_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt11_drpen_in                           : in   std_logic;
    gt11_drprdy_out                         : out  std_logic;
    gt11_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt11_eyescanreset_in                    : in   std_logic;
    gt11_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt11_eyescandataerror_out               : out  std_logic;
    gt11_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt11_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt11_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt11_rxusrclk_in                        : in   std_logic;
    gt11_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt11_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt11_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt11_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt11_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt11_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt11_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt11_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt11_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt11_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt11_rxoutclk_out                       : out  std_logic;
    gt11_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt11_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt11_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt11_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt11_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt11_gttxreset_in                       : in   std_logic;
    gt11_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt11_txusrclk_in                        : in   std_logic;
    gt11_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt11_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt11_gthtxn_out                         : out  std_logic;
    gt11_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt11_txoutclk_out                       : out  std_logic;
    gt11_txoutclkfabric_out                 : out  std_logic;
    gt11_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt11_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt11_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT12  (X1Y16)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt12_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt12_drpclk_in                          : in   std_logic;
    gt12_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt12_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt12_drpen_in                           : in   std_logic;
    gt12_drprdy_out                         : out  std_logic;
    gt12_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt12_eyescanreset_in                    : in   std_logic;
    gt12_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt12_eyescandataerror_out               : out  std_logic;
    gt12_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt12_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt12_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt12_rxusrclk_in                        : in   std_logic;
    gt12_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt12_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt12_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt12_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt12_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt12_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt12_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt12_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt12_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt12_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt12_rxoutclk_out                       : out  std_logic;
    gt12_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt12_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt12_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt12_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt12_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt12_gttxreset_in                       : in   std_logic;
    gt12_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt12_txusrclk_in                        : in   std_logic;
    gt12_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt12_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt12_gthtxn_out                         : out  std_logic;
    gt12_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt12_txoutclk_out                       : out  std_logic;
    gt12_txoutclkfabric_out                 : out  std_logic;
    gt12_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt12_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt12_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT13  (X1Y17)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt13_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt13_drpclk_in                          : in   std_logic;
    gt13_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt13_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt13_drpen_in                           : in   std_logic;
    gt13_drprdy_out                         : out  std_logic;
    gt13_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt13_eyescanreset_in                    : in   std_logic;
    gt13_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt13_eyescandataerror_out               : out  std_logic;
    gt13_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt13_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt13_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt13_rxusrclk_in                        : in   std_logic;
    gt13_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt13_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt13_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt13_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt13_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt13_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt13_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt13_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt13_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt13_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt13_rxoutclk_out                       : out  std_logic;
    gt13_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt13_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt13_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt13_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt13_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt13_gttxreset_in                       : in   std_logic;
    gt13_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt13_txusrclk_in                        : in   std_logic;
    gt13_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt13_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt13_gthtxn_out                         : out  std_logic;
    gt13_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt13_txoutclk_out                       : out  std_logic;
    gt13_txoutclkfabric_out                 : out  std_logic;
    gt13_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt13_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt13_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT14  (X1Y18)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt14_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt14_drpclk_in                          : in   std_logic;
    gt14_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt14_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt14_drpen_in                           : in   std_logic;
    gt14_drprdy_out                         : out  std_logic;
    gt14_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt14_eyescanreset_in                    : in   std_logic;
    gt14_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt14_eyescandataerror_out               : out  std_logic;
    gt14_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt14_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt14_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt14_rxusrclk_in                        : in   std_logic;
    gt14_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt14_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt14_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt14_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt14_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt14_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt14_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt14_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt14_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt14_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt14_rxoutclk_out                       : out  std_logic;
    gt14_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt14_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt14_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt14_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt14_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt14_gttxreset_in                       : in   std_logic;
    gt14_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt14_txusrclk_in                        : in   std_logic;
    gt14_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt14_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt14_gthtxn_out                         : out  std_logic;
    gt14_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt14_txoutclk_out                       : out  std_logic;
    gt14_txoutclkfabric_out                 : out  std_logic;
    gt14_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt14_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt14_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT15  (X1Y19)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt15_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt15_drpclk_in                          : in   std_logic;
    gt15_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt15_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt15_drpen_in                           : in   std_logic;
    gt15_drprdy_out                         : out  std_logic;
    gt15_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt15_eyescanreset_in                    : in   std_logic;
    gt15_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt15_eyescandataerror_out               : out  std_logic;
    gt15_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt15_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt15_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt15_rxusrclk_in                        : in   std_logic;
    gt15_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt15_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt15_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt15_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt15_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt15_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt15_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt15_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt15_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt15_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt15_rxoutclk_out                       : out  std_logic;
    gt15_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt15_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt15_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt15_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt15_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt15_gttxreset_in                       : in   std_logic;
    gt15_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt15_txusrclk_in                        : in   std_logic;
    gt15_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt15_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt15_gthtxn_out                         : out  std_logic;
    gt15_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt15_txoutclk_out                       : out  std_logic;
    gt15_txoutclkfabric_out                 : out  std_logic;
    gt15_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt15_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt15_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT16  (X1Y20)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt16_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt16_drpclk_in                          : in   std_logic;
    gt16_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt16_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt16_drpen_in                           : in   std_logic;
    gt16_drprdy_out                         : out  std_logic;
    gt16_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt16_eyescanreset_in                    : in   std_logic;
    gt16_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt16_eyescandataerror_out               : out  std_logic;
    gt16_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt16_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt16_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt16_rxusrclk_in                        : in   std_logic;
    gt16_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt16_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt16_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt16_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt16_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt16_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt16_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt16_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt16_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt16_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt16_rxoutclk_out                       : out  std_logic;
    gt16_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt16_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt16_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt16_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt16_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt16_gttxreset_in                       : in   std_logic;
    gt16_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt16_txusrclk_in                        : in   std_logic;
    gt16_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt16_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt16_gthtxn_out                         : out  std_logic;
    gt16_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt16_txoutclk_out                       : out  std_logic;
    gt16_txoutclkfabric_out                 : out  std_logic;
    gt16_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt16_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt16_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT17  (X1Y21)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt17_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt17_drpclk_in                          : in   std_logic;
    gt17_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt17_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt17_drpen_in                           : in   std_logic;
    gt17_drprdy_out                         : out  std_logic;
    gt17_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt17_eyescanreset_in                    : in   std_logic;
    gt17_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt17_eyescandataerror_out               : out  std_logic;
    gt17_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt17_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt17_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt17_rxusrclk_in                        : in   std_logic;
    gt17_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt17_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt17_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt17_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt17_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt17_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt17_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt17_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt17_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt17_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt17_rxoutclk_out                       : out  std_logic;
    gt17_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt17_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt17_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt17_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt17_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt17_gttxreset_in                       : in   std_logic;
    gt17_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt17_txusrclk_in                        : in   std_logic;
    gt17_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt17_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt17_gthtxn_out                         : out  std_logic;
    gt17_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt17_txoutclk_out                       : out  std_logic;
    gt17_txoutclkfabric_out                 : out  std_logic;
    gt17_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt17_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt17_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT18  (X1Y22)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt18_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt18_drpclk_in                          : in   std_logic;
    gt18_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt18_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt18_drpen_in                           : in   std_logic;
    gt18_drprdy_out                         : out  std_logic;
    gt18_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt18_eyescanreset_in                    : in   std_logic;
    gt18_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt18_eyescandataerror_out               : out  std_logic;
    gt18_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt18_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt18_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt18_rxusrclk_in                        : in   std_logic;
    gt18_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt18_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt18_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt18_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt18_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt18_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt18_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt18_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt18_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt18_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt18_rxoutclk_out                       : out  std_logic;
    gt18_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt18_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt18_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt18_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt18_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt18_gttxreset_in                       : in   std_logic;
    gt18_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt18_txusrclk_in                        : in   std_logic;
    gt18_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt18_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt18_gthtxn_out                         : out  std_logic;
    gt18_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt18_txoutclk_out                       : out  std_logic;
    gt18_txoutclkfabric_out                 : out  std_logic;
    gt18_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt18_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt18_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT19  (X1Y23)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt19_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt19_drpclk_in                          : in   std_logic;
    gt19_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt19_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt19_drpen_in                           : in   std_logic;
    gt19_drprdy_out                         : out  std_logic;
    gt19_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt19_eyescanreset_in                    : in   std_logic;
    gt19_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt19_eyescandataerror_out               : out  std_logic;
    gt19_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt19_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt19_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt19_rxusrclk_in                        : in   std_logic;
    gt19_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt19_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt19_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt19_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt19_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt19_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt19_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt19_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt19_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt19_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt19_rxoutclk_out                       : out  std_logic;
    gt19_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt19_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt19_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt19_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt19_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt19_gttxreset_in                       : in   std_logic;
    gt19_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt19_txusrclk_in                        : in   std_logic;
    gt19_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt19_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt19_gthtxn_out                         : out  std_logic;
    gt19_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt19_txoutclk_out                       : out  std_logic;
    gt19_txoutclkfabric_out                 : out  std_logic;
    gt19_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt19_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt19_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT20  (X1Y24)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt20_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt20_drpclk_in                          : in   std_logic;
    gt20_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt20_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt20_drpen_in                           : in   std_logic;
    gt20_drprdy_out                         : out  std_logic;
    gt20_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt20_eyescanreset_in                    : in   std_logic;
    gt20_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt20_eyescandataerror_out               : out  std_logic;
    gt20_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt20_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt20_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt20_rxusrclk_in                        : in   std_logic;
    gt20_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt20_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt20_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt20_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt20_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt20_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt20_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt20_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt20_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt20_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt20_rxoutclk_out                       : out  std_logic;
    gt20_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt20_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt20_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt20_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt20_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt20_gttxreset_in                       : in   std_logic;
    gt20_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt20_txusrclk_in                        : in   std_logic;
    gt20_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt20_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt20_gthtxn_out                         : out  std_logic;
    gt20_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt20_txoutclk_out                       : out  std_logic;
    gt20_txoutclkfabric_out                 : out  std_logic;
    gt20_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt20_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt20_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT21  (X1Y25)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt21_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt21_drpclk_in                          : in   std_logic;
    gt21_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt21_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt21_drpen_in                           : in   std_logic;
    gt21_drprdy_out                         : out  std_logic;
    gt21_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt21_eyescanreset_in                    : in   std_logic;
    gt21_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt21_eyescandataerror_out               : out  std_logic;
    gt21_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt21_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt21_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt21_rxusrclk_in                        : in   std_logic;
    gt21_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt21_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt21_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt21_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt21_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt21_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt21_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt21_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt21_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt21_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt21_rxoutclk_out                       : out  std_logic;
    gt21_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt21_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt21_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt21_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt21_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt21_gttxreset_in                       : in   std_logic;
    gt21_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt21_txusrclk_in                        : in   std_logic;
    gt21_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt21_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt21_gthtxn_out                         : out  std_logic;
    gt21_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt21_txoutclk_out                       : out  std_logic;
    gt21_txoutclkfabric_out                 : out  std_logic;
    gt21_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt21_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt21_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT22  (X1Y26)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt22_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt22_drpclk_in                          : in   std_logic;
    gt22_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt22_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt22_drpen_in                           : in   std_logic;
    gt22_drprdy_out                         : out  std_logic;
    gt22_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt22_eyescanreset_in                    : in   std_logic;
    gt22_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt22_eyescandataerror_out               : out  std_logic;
    gt22_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt22_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt22_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt22_rxusrclk_in                        : in   std_logic;
    gt22_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt22_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt22_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt22_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt22_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt22_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt22_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt22_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt22_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt22_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt22_rxoutclk_out                       : out  std_logic;
    gt22_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt22_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt22_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt22_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt22_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt22_gttxreset_in                       : in   std_logic;
    gt22_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt22_txusrclk_in                        : in   std_logic;
    gt22_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt22_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt22_gthtxn_out                         : out  std_logic;
    gt22_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt22_txoutclk_out                       : out  std_logic;
    gt22_txoutclkfabric_out                 : out  std_logic;
    gt22_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt22_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt22_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT23  (X1Y27)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt23_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt23_drpclk_in                          : in   std_logic;
    gt23_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt23_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt23_drpen_in                           : in   std_logic;
    gt23_drprdy_out                         : out  std_logic;
    gt23_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt23_eyescanreset_in                    : in   std_logic;
    gt23_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt23_eyescandataerror_out               : out  std_logic;
    gt23_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt23_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt23_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt23_rxusrclk_in                        : in   std_logic;
    gt23_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt23_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt23_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt23_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt23_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt23_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt23_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt23_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt23_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt23_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt23_rxoutclk_out                       : out  std_logic;
    gt23_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt23_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt23_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt23_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt23_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt23_gttxreset_in                       : in   std_logic;
    gt23_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt23_txusrclk_in                        : in   std_logic;
    gt23_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt23_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt23_gthtxn_out                         : out  std_logic;
    gt23_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt23_txoutclk_out                       : out  std_logic;
    gt23_txoutclkfabric_out                 : out  std_logic;
    gt23_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt23_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt23_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT24  (X1Y28)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt24_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt24_drpclk_in                          : in   std_logic;
    gt24_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt24_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt24_drpen_in                           : in   std_logic;
    gt24_drprdy_out                         : out  std_logic;
    gt24_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt24_eyescanreset_in                    : in   std_logic;
    gt24_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt24_eyescandataerror_out               : out  std_logic;
    gt24_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt24_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt24_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt24_rxusrclk_in                        : in   std_logic;
    gt24_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt24_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt24_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt24_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt24_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt24_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt24_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt24_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt24_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt24_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt24_rxoutclk_out                       : out  std_logic;
    gt24_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt24_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt24_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt24_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt24_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt24_gttxreset_in                       : in   std_logic;
    gt24_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt24_txusrclk_in                        : in   std_logic;
    gt24_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt24_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt24_gthtxn_out                         : out  std_logic;
    gt24_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt24_txoutclk_out                       : out  std_logic;
    gt24_txoutclkfabric_out                 : out  std_logic;
    gt24_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt24_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt24_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT25  (X1Y29)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt25_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt25_drpclk_in                          : in   std_logic;
    gt25_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt25_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt25_drpen_in                           : in   std_logic;
    gt25_drprdy_out                         : out  std_logic;
    gt25_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt25_eyescanreset_in                    : in   std_logic;
    gt25_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt25_eyescandataerror_out               : out  std_logic;
    gt25_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt25_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt25_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt25_rxusrclk_in                        : in   std_logic;
    gt25_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt25_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt25_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt25_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt25_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt25_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt25_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt25_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt25_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt25_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt25_rxoutclk_out                       : out  std_logic;
    gt25_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt25_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt25_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt25_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt25_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt25_gttxreset_in                       : in   std_logic;
    gt25_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt25_txusrclk_in                        : in   std_logic;
    gt25_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt25_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt25_gthtxn_out                         : out  std_logic;
    gt25_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt25_txoutclk_out                       : out  std_logic;
    gt25_txoutclkfabric_out                 : out  std_logic;
    gt25_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt25_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt25_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT26  (X1Y30)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt26_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt26_drpclk_in                          : in   std_logic;
    gt26_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt26_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt26_drpen_in                           : in   std_logic;
    gt26_drprdy_out                         : out  std_logic;
    gt26_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt26_eyescanreset_in                    : in   std_logic;
    gt26_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt26_eyescandataerror_out               : out  std_logic;
    gt26_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt26_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt26_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt26_rxusrclk_in                        : in   std_logic;
    gt26_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt26_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt26_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt26_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt26_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt26_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt26_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt26_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt26_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt26_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt26_rxoutclk_out                       : out  std_logic;
    gt26_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt26_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt26_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt26_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt26_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt26_gttxreset_in                       : in   std_logic;
    gt26_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt26_txusrclk_in                        : in   std_logic;
    gt26_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt26_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt26_gthtxn_out                         : out  std_logic;
    gt26_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt26_txoutclk_out                       : out  std_logic;
    gt26_txoutclkfabric_out                 : out  std_logic;
    gt26_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt26_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt26_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT27  (X1Y31)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt27_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt27_drpclk_in                          : in   std_logic;
    gt27_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt27_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt27_drpen_in                           : in   std_logic;
    gt27_drprdy_out                         : out  std_logic;
    gt27_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt27_eyescanreset_in                    : in   std_logic;
    gt27_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt27_eyescandataerror_out               : out  std_logic;
    gt27_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt27_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt27_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt27_rxusrclk_in                        : in   std_logic;
    gt27_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt27_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt27_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt27_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt27_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt27_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt27_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt27_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt27_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt27_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt27_rxoutclk_out                       : out  std_logic;
    gt27_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt27_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt27_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt27_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt27_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt27_gttxreset_in                       : in   std_logic;
    gt27_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt27_txusrclk_in                        : in   std_logic;
    gt27_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt27_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt27_gthtxn_out                         : out  std_logic;
    gt27_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt27_txoutclk_out                       : out  std_logic;
    gt27_txoutclkfabric_out                 : out  std_logic;
    gt27_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt27_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt27_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT28  (X1Y32)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt28_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt28_drpclk_in                          : in   std_logic;
    gt28_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt28_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt28_drpen_in                           : in   std_logic;
    gt28_drprdy_out                         : out  std_logic;
    gt28_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt28_eyescanreset_in                    : in   std_logic;
    gt28_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt28_eyescandataerror_out               : out  std_logic;
    gt28_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt28_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt28_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt28_rxusrclk_in                        : in   std_logic;
    gt28_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt28_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt28_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt28_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt28_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt28_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt28_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt28_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt28_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt28_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt28_rxoutclk_out                       : out  std_logic;
    gt28_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt28_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt28_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt28_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt28_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt28_gttxreset_in                       : in   std_logic;
    gt28_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt28_txusrclk_in                        : in   std_logic;
    gt28_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt28_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt28_gthtxn_out                         : out  std_logic;
    gt28_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt28_txoutclk_out                       : out  std_logic;
    gt28_txoutclkfabric_out                 : out  std_logic;
    gt28_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt28_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt28_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT29  (X1Y33)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt29_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt29_drpclk_in                          : in   std_logic;
    gt29_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt29_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt29_drpen_in                           : in   std_logic;
    gt29_drprdy_out                         : out  std_logic;
    gt29_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt29_eyescanreset_in                    : in   std_logic;
    gt29_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt29_eyescandataerror_out               : out  std_logic;
    gt29_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt29_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt29_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt29_rxusrclk_in                        : in   std_logic;
    gt29_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt29_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt29_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt29_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt29_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt29_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt29_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt29_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt29_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt29_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt29_rxoutclk_out                       : out  std_logic;
    gt29_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt29_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt29_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt29_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt29_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt29_gttxreset_in                       : in   std_logic;
    gt29_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt29_txusrclk_in                        : in   std_logic;
    gt29_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt29_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt29_gthtxn_out                         : out  std_logic;
    gt29_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt29_txoutclk_out                       : out  std_logic;
    gt29_txoutclkfabric_out                 : out  std_logic;
    gt29_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt29_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt29_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT30  (X1Y34)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt30_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt30_drpclk_in                          : in   std_logic;
    gt30_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt30_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt30_drpen_in                           : in   std_logic;
    gt30_drprdy_out                         : out  std_logic;
    gt30_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt30_eyescanreset_in                    : in   std_logic;
    gt30_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt30_eyescandataerror_out               : out  std_logic;
    gt30_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt30_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt30_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt30_rxusrclk_in                        : in   std_logic;
    gt30_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt30_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt30_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt30_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt30_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt30_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt30_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt30_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt30_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt30_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt30_rxoutclk_out                       : out  std_logic;
    gt30_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt30_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt30_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt30_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt30_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt30_gttxreset_in                       : in   std_logic;
    gt30_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt30_txusrclk_in                        : in   std_logic;
    gt30_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt30_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt30_gthtxn_out                         : out  std_logic;
    gt30_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt30_txoutclk_out                       : out  std_logic;
    gt30_txoutclkfabric_out                 : out  std_logic;
    gt30_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt30_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt30_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT31  (X1Y35)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt31_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt31_drpclk_in                          : in   std_logic;
    gt31_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt31_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt31_drpen_in                           : in   std_logic;
    gt31_drprdy_out                         : out  std_logic;
    gt31_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt31_eyescanreset_in                    : in   std_logic;
    gt31_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt31_eyescandataerror_out               : out  std_logic;
    gt31_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt31_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt31_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt31_rxusrclk_in                        : in   std_logic;
    gt31_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt31_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt31_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt31_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt31_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt31_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt31_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt31_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt31_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt31_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt31_rxoutclk_out                       : out  std_logic;
    gt31_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt31_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt31_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt31_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt31_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt31_gttxreset_in                       : in   std_logic;
    gt31_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt31_txusrclk_in                        : in   std_logic;
    gt31_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt31_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt31_gthtxn_out                         : out  std_logic;
    gt31_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt31_txoutclk_out                       : out  std_logic;
    gt31_txoutclkfabric_out                 : out  std_logic;
    gt31_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt31_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt31_txcharisk_in                       : in   std_logic_vector(7 downto 0);


    --____________________________COMMON PORTS________________________________
    GT0_QPLLLOCK_IN : in std_logic;
    GT0_QPLLREFCLKLOST_IN  : in std_logic;
    GT0_QPLLRESET_OUT  : out std_logic;
     GT0_QPLLOUTCLK_IN  : in std_logic;
     GT0_QPLLOUTREFCLK_IN : in std_logic;
    --____________________________COMMON PORTS________________________________
    GT1_QPLLLOCK_IN : in std_logic;
    GT1_QPLLREFCLKLOST_IN  : in std_logic;
    GT1_QPLLRESET_OUT  : out std_logic;
     GT1_QPLLOUTCLK_IN  : in std_logic;
     GT1_QPLLOUTREFCLK_IN : in std_logic;
    --____________________________COMMON PORTS________________________________
    GT2_QPLLLOCK_IN : in std_logic;
    GT2_QPLLREFCLKLOST_IN  : in std_logic;
    GT2_QPLLRESET_OUT  : out std_logic;
     GT2_QPLLOUTCLK_IN  : in std_logic;
     GT2_QPLLOUTREFCLK_IN : in std_logic;
    --____________________________COMMON PORTS________________________________
    GT3_QPLLLOCK_IN : in std_logic;
    GT3_QPLLREFCLKLOST_IN  : in std_logic;
    GT3_QPLLRESET_OUT  : out std_logic;
     GT3_QPLLOUTCLK_IN  : in std_logic;
     GT3_QPLLOUTREFCLK_IN : in std_logic;
    --____________________________COMMON PORTS________________________________
    GT4_QPLLLOCK_IN : in std_logic;
    GT4_QPLLREFCLKLOST_IN  : in std_logic;
    GT4_QPLLRESET_OUT  : out std_logic;
     GT4_QPLLOUTCLK_IN  : in std_logic;
     GT4_QPLLOUTREFCLK_IN : in std_logic;
    --____________________________COMMON PORTS________________________________
    GT5_QPLLLOCK_IN : in std_logic;
    GT5_QPLLREFCLKLOST_IN  : in std_logic;
    GT5_QPLLRESET_OUT  : out std_logic;
     GT5_QPLLOUTCLK_IN  : in std_logic;
     GT5_QPLLOUTREFCLK_IN : in std_logic;
    --____________________________COMMON PORTS________________________________
    GT6_QPLLLOCK_IN : in std_logic;
    GT6_QPLLREFCLKLOST_IN  : in std_logic;
    GT6_QPLLRESET_OUT  : out std_logic;
     GT6_QPLLOUTCLK_IN  : in std_logic;
     GT6_QPLLOUTREFCLK_IN : in std_logic;
    --____________________________COMMON PORTS________________________________
    GT7_QPLLLOCK_IN : in std_logic;
    GT7_QPLLREFCLKLOST_IN  : in std_logic;
    GT7_QPLLRESET_OUT  : out std_logic;
     GT7_QPLLOUTCLK_IN  : in std_logic;
     GT7_QPLLOUTREFCLK_IN : in std_logic

);

end gtwizard_0_init;
    
architecture RTL of gtwizard_0_init is
attribute DowngradeIPIdentifiedWarnings: string;
attribute DowngradeIPIdentifiedWarnings of RTL : architecture is "yes";

--**************************Component Declarations*****************************


component gtwizard_0_multi_gt 
generic
(
    -- Simulation attributes
    EXAMPLE_SIMULATION             : integer   := 0;      -- Set to 1 for simulation
    WRAPPER_SIM_GTRESET_SPEEDUP    : string    := "FALSE" -- Set to "TRUE" to speed up sim reset

);
port
(

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT0  (X1Y4)
    --____________________________CHANNEL PORTS________________________________
    GT0_DRP_BUSY_OUT                        : out  std_logic;
    GT0_RXPMARESETDONE_OUT                        : out  std_logic;
    GT0_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt0_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt0_drpclk_in                           : in   std_logic;
    gt0_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt0_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt0_drpen_in                            : in   std_logic;
    gt0_drprdy_out                          : out  std_logic;
    gt0_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt0_eyescanreset_in                     : in   std_logic;
    gt0_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt0_eyescandataerror_out                : out  std_logic;
    gt0_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt0_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt0_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt0_rxusrclk_in                         : in   std_logic;
    gt0_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt0_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt0_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt0_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt0_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt0_rxdlyen_in                          : in   std_logic;
    gt0_rxdlysreset_in                      : in   std_logic;
    gt0_rxdlysresetdone_out                 : out  std_logic;
    gt0_rxphalign_in                        : in   std_logic;
    gt0_rxphaligndone_out                   : out  std_logic;
    gt0_rxphalignen_in                      : in   std_logic;
    gt0_rxphdlyreset_in                     : in   std_logic;
    gt0_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt0_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    gt0_rxsyncallin_in                      : in   std_logic;
    gt0_rxsyncdone_out                      : out  std_logic;
    gt0_rxsyncin_in                         : in   std_logic;
    gt0_rxsyncmode_in                       : in   std_logic;
    gt0_rxsyncout_out                       : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt0_rxbyteisaligned_out                 : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt0_rxlpmhfhold_in                      : in   std_logic;
    gt0_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt0_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt0_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt0_rxoutclk_out                        : out  std_logic;
    gt0_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt0_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt0_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt0_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt0_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt0_gttxreset_in                        : in   std_logic;
    gt0_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt0_txusrclk_in                         : in   std_logic;
    gt0_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt0_txdlyen_in                          : in   std_logic;
    gt0_txdlysreset_in                      : in   std_logic;
    gt0_txdlysresetdone_out                 : out  std_logic;
    gt0_txphalign_in                        : in   std_logic;
    gt0_txphaligndone_out                   : out  std_logic;
    gt0_txphalignen_in                      : in   std_logic;
    gt0_txphdlyreset_in                     : in   std_logic;
    gt0_txphinit_in                         : in   std_logic;
    gt0_txphinitdone_out                    : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt0_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt0_gthtxn_out                          : out  std_logic;
    gt0_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt0_txoutclk_out                        : out  std_logic;
    gt0_txoutclkfabric_out                  : out  std_logic;
    gt0_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt0_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt0_txcharisk_in                        : in   std_logic_vector(7 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT1  (X1Y5)
    --____________________________CHANNEL PORTS________________________________
    GT1_DRP_BUSY_OUT                        : out  std_logic;
    GT1_RXPMARESETDONE_OUT                        : out  std_logic;
    GT1_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt1_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt1_drpclk_in                           : in   std_logic;
    gt1_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt1_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt1_drpen_in                            : in   std_logic;
    gt1_drprdy_out                          : out  std_logic;
    gt1_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt1_eyescanreset_in                     : in   std_logic;
    gt1_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt1_eyescandataerror_out                : out  std_logic;
    gt1_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt1_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt1_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt1_rxusrclk_in                         : in   std_logic;
    gt1_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt1_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt1_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt1_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt1_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt1_rxdlyen_in                          : in   std_logic;
    gt1_rxdlysreset_in                      : in   std_logic;
    gt1_rxdlysresetdone_out                 : out  std_logic;
    gt1_rxphalign_in                        : in   std_logic;
    gt1_rxphaligndone_out                   : out  std_logic;
    gt1_rxphalignen_in                      : in   std_logic;
    gt1_rxphdlyreset_in                     : in   std_logic;
    gt1_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt1_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    gt1_rxsyncallin_in                      : in   std_logic;
    gt1_rxsyncdone_out                      : out  std_logic;
    gt1_rxsyncin_in                         : in   std_logic;
    gt1_rxsyncmode_in                       : in   std_logic;
    gt1_rxsyncout_out                       : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt1_rxbyteisaligned_out                 : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt1_rxlpmhfhold_in                      : in   std_logic;
    gt1_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt1_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt1_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt1_rxoutclk_out                        : out  std_logic;
    gt1_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt1_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt1_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt1_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt1_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt1_gttxreset_in                        : in   std_logic;
    gt1_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt1_txusrclk_in                         : in   std_logic;
    gt1_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt1_txdlyen_in                          : in   std_logic;
    gt1_txdlysreset_in                      : in   std_logic;
    gt1_txdlysresetdone_out                 : out  std_logic;
    gt1_txphalign_in                        : in   std_logic;
    gt1_txphaligndone_out                   : out  std_logic;
    gt1_txphalignen_in                      : in   std_logic;
    gt1_txphdlyreset_in                     : in   std_logic;
    gt1_txphinit_in                         : in   std_logic;
    gt1_txphinitdone_out                    : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt1_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt1_gthtxn_out                          : out  std_logic;
    gt1_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt1_txoutclk_out                        : out  std_logic;
    gt1_txoutclkfabric_out                  : out  std_logic;
    gt1_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt1_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt1_txcharisk_in                        : in   std_logic_vector(7 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT2  (X1Y6)
    --____________________________CHANNEL PORTS________________________________
    GT2_DRP_BUSY_OUT                        : out  std_logic;
    GT2_RXPMARESETDONE_OUT                        : out  std_logic;
    GT2_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt2_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt2_drpclk_in                           : in   std_logic;
    gt2_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt2_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt2_drpen_in                            : in   std_logic;
    gt2_drprdy_out                          : out  std_logic;
    gt2_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt2_eyescanreset_in                     : in   std_logic;
    gt2_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt2_eyescandataerror_out                : out  std_logic;
    gt2_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt2_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt2_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt2_rxusrclk_in                         : in   std_logic;
    gt2_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt2_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt2_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt2_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt2_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt2_rxdlyen_in                          : in   std_logic;
    gt2_rxdlysreset_in                      : in   std_logic;
    gt2_rxdlysresetdone_out                 : out  std_logic;
    gt2_rxphalign_in                        : in   std_logic;
    gt2_rxphaligndone_out                   : out  std_logic;
    gt2_rxphalignen_in                      : in   std_logic;
    gt2_rxphdlyreset_in                     : in   std_logic;
    gt2_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt2_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    gt2_rxsyncallin_in                      : in   std_logic;
    gt2_rxsyncdone_out                      : out  std_logic;
    gt2_rxsyncin_in                         : in   std_logic;
    gt2_rxsyncmode_in                       : in   std_logic;
    gt2_rxsyncout_out                       : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt2_rxbyteisaligned_out                 : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt2_rxlpmhfhold_in                      : in   std_logic;
    gt2_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt2_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt2_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt2_rxoutclk_out                        : out  std_logic;
    gt2_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt2_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt2_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt2_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt2_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt2_gttxreset_in                        : in   std_logic;
    gt2_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt2_txusrclk_in                         : in   std_logic;
    gt2_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt2_txdlyen_in                          : in   std_logic;
    gt2_txdlysreset_in                      : in   std_logic;
    gt2_txdlysresetdone_out                 : out  std_logic;
    gt2_txphalign_in                        : in   std_logic;
    gt2_txphaligndone_out                   : out  std_logic;
    gt2_txphalignen_in                      : in   std_logic;
    gt2_txphdlyreset_in                     : in   std_logic;
    gt2_txphinit_in                         : in   std_logic;
    gt2_txphinitdone_out                    : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt2_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt2_gthtxn_out                          : out  std_logic;
    gt2_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt2_txoutclk_out                        : out  std_logic;
    gt2_txoutclkfabric_out                  : out  std_logic;
    gt2_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt2_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt2_txcharisk_in                        : in   std_logic_vector(7 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT3  (X1Y7)
    --____________________________CHANNEL PORTS________________________________
    GT3_DRP_BUSY_OUT                        : out  std_logic;
    GT3_RXPMARESETDONE_OUT                        : out  std_logic;
    GT3_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt3_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt3_drpclk_in                           : in   std_logic;
    gt3_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt3_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt3_drpen_in                            : in   std_logic;
    gt3_drprdy_out                          : out  std_logic;
    gt3_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt3_eyescanreset_in                     : in   std_logic;
    gt3_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt3_eyescandataerror_out                : out  std_logic;
    gt3_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt3_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt3_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt3_rxusrclk_in                         : in   std_logic;
    gt3_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt3_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt3_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt3_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt3_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt3_rxdlyen_in                          : in   std_logic;
    gt3_rxdlysreset_in                      : in   std_logic;
    gt3_rxdlysresetdone_out                 : out  std_logic;
    gt3_rxphalign_in                        : in   std_logic;
    gt3_rxphaligndone_out                   : out  std_logic;
    gt3_rxphalignen_in                      : in   std_logic;
    gt3_rxphdlyreset_in                     : in   std_logic;
    gt3_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt3_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    gt3_rxsyncallin_in                      : in   std_logic;
    gt3_rxsyncdone_out                      : out  std_logic;
    gt3_rxsyncin_in                         : in   std_logic;
    gt3_rxsyncmode_in                       : in   std_logic;
    gt3_rxsyncout_out                       : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt3_rxbyteisaligned_out                 : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt3_rxlpmhfhold_in                      : in   std_logic;
    gt3_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt3_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt3_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt3_rxoutclk_out                        : out  std_logic;
    gt3_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt3_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt3_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt3_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt3_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt3_gttxreset_in                        : in   std_logic;
    gt3_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt3_txusrclk_in                         : in   std_logic;
    gt3_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt3_txdlyen_in                          : in   std_logic;
    gt3_txdlysreset_in                      : in   std_logic;
    gt3_txdlysresetdone_out                 : out  std_logic;
    gt3_txphalign_in                        : in   std_logic;
    gt3_txphaligndone_out                   : out  std_logic;
    gt3_txphalignen_in                      : in   std_logic;
    gt3_txphdlyreset_in                     : in   std_logic;
    gt3_txphinit_in                         : in   std_logic;
    gt3_txphinitdone_out                    : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt3_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt3_gthtxn_out                          : out  std_logic;
    gt3_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt3_txoutclk_out                        : out  std_logic;
    gt3_txoutclkfabric_out                  : out  std_logic;
    gt3_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt3_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt3_txcharisk_in                        : in   std_logic_vector(7 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT4  (X1Y8)
    --____________________________CHANNEL PORTS________________________________
    GT4_DRP_BUSY_OUT                        : out  std_logic;
    GT4_RXPMARESETDONE_OUT                        : out  std_logic;
    GT4_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt4_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt4_drpclk_in                           : in   std_logic;
    gt4_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt4_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt4_drpen_in                            : in   std_logic;
    gt4_drprdy_out                          : out  std_logic;
    gt4_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt4_eyescanreset_in                     : in   std_logic;
    gt4_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt4_eyescandataerror_out                : out  std_logic;
    gt4_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt4_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt4_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt4_rxusrclk_in                         : in   std_logic;
    gt4_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt4_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt4_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt4_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt4_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt4_rxdlyen_in                          : in   std_logic;
    gt4_rxdlysreset_in                      : in   std_logic;
    gt4_rxdlysresetdone_out                 : out  std_logic;
    gt4_rxphalign_in                        : in   std_logic;
    gt4_rxphaligndone_out                   : out  std_logic;
    gt4_rxphalignen_in                      : in   std_logic;
    gt4_rxphdlyreset_in                     : in   std_logic;
    gt4_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt4_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    gt4_rxsyncallin_in                      : in   std_logic;
    gt4_rxsyncdone_out                      : out  std_logic;
    gt4_rxsyncin_in                         : in   std_logic;
    gt4_rxsyncmode_in                       : in   std_logic;
    gt4_rxsyncout_out                       : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt4_rxbyteisaligned_out                 : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt4_rxlpmhfhold_in                      : in   std_logic;
    gt4_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt4_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt4_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt4_rxoutclk_out                        : out  std_logic;
    gt4_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt4_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt4_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt4_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt4_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt4_gttxreset_in                        : in   std_logic;
    gt4_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt4_txusrclk_in                         : in   std_logic;
    gt4_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt4_txdlyen_in                          : in   std_logic;
    gt4_txdlysreset_in                      : in   std_logic;
    gt4_txdlysresetdone_out                 : out  std_logic;
    gt4_txphalign_in                        : in   std_logic;
    gt4_txphaligndone_out                   : out  std_logic;
    gt4_txphalignen_in                      : in   std_logic;
    gt4_txphdlyreset_in                     : in   std_logic;
    gt4_txphinit_in                         : in   std_logic;
    gt4_txphinitdone_out                    : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt4_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt4_gthtxn_out                          : out  std_logic;
    gt4_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt4_txoutclk_out                        : out  std_logic;
    gt4_txoutclkfabric_out                  : out  std_logic;
    gt4_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt4_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt4_txcharisk_in                        : in   std_logic_vector(7 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT5  (X1Y9)
    --____________________________CHANNEL PORTS________________________________
    GT5_DRP_BUSY_OUT                        : out  std_logic;
    GT5_RXPMARESETDONE_OUT                        : out  std_logic;
    GT5_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt5_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt5_drpclk_in                           : in   std_logic;
    gt5_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt5_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt5_drpen_in                            : in   std_logic;
    gt5_drprdy_out                          : out  std_logic;
    gt5_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt5_eyescanreset_in                     : in   std_logic;
    gt5_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt5_eyescandataerror_out                : out  std_logic;
    gt5_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt5_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt5_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt5_rxusrclk_in                         : in   std_logic;
    gt5_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt5_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt5_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt5_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt5_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt5_rxdlyen_in                          : in   std_logic;
    gt5_rxdlysreset_in                      : in   std_logic;
    gt5_rxdlysresetdone_out                 : out  std_logic;
    gt5_rxphalign_in                        : in   std_logic;
    gt5_rxphaligndone_out                   : out  std_logic;
    gt5_rxphalignen_in                      : in   std_logic;
    gt5_rxphdlyreset_in                     : in   std_logic;
    gt5_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt5_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    gt5_rxsyncallin_in                      : in   std_logic;
    gt5_rxsyncdone_out                      : out  std_logic;
    gt5_rxsyncin_in                         : in   std_logic;
    gt5_rxsyncmode_in                       : in   std_logic;
    gt5_rxsyncout_out                       : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt5_rxbyteisaligned_out                 : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt5_rxlpmhfhold_in                      : in   std_logic;
    gt5_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt5_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt5_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt5_rxoutclk_out                        : out  std_logic;
    gt5_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt5_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt5_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt5_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt5_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt5_gttxreset_in                        : in   std_logic;
    gt5_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt5_txusrclk_in                         : in   std_logic;
    gt5_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt5_txdlyen_in                          : in   std_logic;
    gt5_txdlysreset_in                      : in   std_logic;
    gt5_txdlysresetdone_out                 : out  std_logic;
    gt5_txphalign_in                        : in   std_logic;
    gt5_txphaligndone_out                   : out  std_logic;
    gt5_txphalignen_in                      : in   std_logic;
    gt5_txphdlyreset_in                     : in   std_logic;
    gt5_txphinit_in                         : in   std_logic;
    gt5_txphinitdone_out                    : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt5_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt5_gthtxn_out                          : out  std_logic;
    gt5_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt5_txoutclk_out                        : out  std_logic;
    gt5_txoutclkfabric_out                  : out  std_logic;
    gt5_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt5_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt5_txcharisk_in                        : in   std_logic_vector(7 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT6  (X1Y10)
    --____________________________CHANNEL PORTS________________________________
    GT6_DRP_BUSY_OUT                        : out  std_logic;
    GT6_RXPMARESETDONE_OUT                        : out  std_logic;
    GT6_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt6_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt6_drpclk_in                           : in   std_logic;
    gt6_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt6_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt6_drpen_in                            : in   std_logic;
    gt6_drprdy_out                          : out  std_logic;
    gt6_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt6_eyescanreset_in                     : in   std_logic;
    gt6_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt6_eyescandataerror_out                : out  std_logic;
    gt6_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt6_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt6_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt6_rxusrclk_in                         : in   std_logic;
    gt6_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt6_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt6_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt6_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt6_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt6_rxdlyen_in                          : in   std_logic;
    gt6_rxdlysreset_in                      : in   std_logic;
    gt6_rxdlysresetdone_out                 : out  std_logic;
    gt6_rxphalign_in                        : in   std_logic;
    gt6_rxphaligndone_out                   : out  std_logic;
    gt6_rxphalignen_in                      : in   std_logic;
    gt6_rxphdlyreset_in                     : in   std_logic;
    gt6_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt6_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    gt6_rxsyncallin_in                      : in   std_logic;
    gt6_rxsyncdone_out                      : out  std_logic;
    gt6_rxsyncin_in                         : in   std_logic;
    gt6_rxsyncmode_in                       : in   std_logic;
    gt6_rxsyncout_out                       : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt6_rxbyteisaligned_out                 : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt6_rxlpmhfhold_in                      : in   std_logic;
    gt6_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt6_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt6_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt6_rxoutclk_out                        : out  std_logic;
    gt6_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt6_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt6_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt6_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt6_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt6_gttxreset_in                        : in   std_logic;
    gt6_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt6_txusrclk_in                         : in   std_logic;
    gt6_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt6_txdlyen_in                          : in   std_logic;
    gt6_txdlysreset_in                      : in   std_logic;
    gt6_txdlysresetdone_out                 : out  std_logic;
    gt6_txphalign_in                        : in   std_logic;
    gt6_txphaligndone_out                   : out  std_logic;
    gt6_txphalignen_in                      : in   std_logic;
    gt6_txphdlyreset_in                     : in   std_logic;
    gt6_txphinit_in                         : in   std_logic;
    gt6_txphinitdone_out                    : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt6_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt6_gthtxn_out                          : out  std_logic;
    gt6_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt6_txoutclk_out                        : out  std_logic;
    gt6_txoutclkfabric_out                  : out  std_logic;
    gt6_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt6_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt6_txcharisk_in                        : in   std_logic_vector(7 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT7  (X1Y11)
    --____________________________CHANNEL PORTS________________________________
    GT7_DRP_BUSY_OUT                        : out  std_logic;
    GT7_RXPMARESETDONE_OUT                        : out  std_logic;
    GT7_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt7_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt7_drpclk_in                           : in   std_logic;
    gt7_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt7_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt7_drpen_in                            : in   std_logic;
    gt7_drprdy_out                          : out  std_logic;
    gt7_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt7_eyescanreset_in                     : in   std_logic;
    gt7_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt7_eyescandataerror_out                : out  std_logic;
    gt7_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt7_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt7_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt7_rxusrclk_in                         : in   std_logic;
    gt7_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt7_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt7_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt7_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt7_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt7_rxdlyen_in                          : in   std_logic;
    gt7_rxdlysreset_in                      : in   std_logic;
    gt7_rxdlysresetdone_out                 : out  std_logic;
    gt7_rxphalign_in                        : in   std_logic;
    gt7_rxphaligndone_out                   : out  std_logic;
    gt7_rxphalignen_in                      : in   std_logic;
    gt7_rxphdlyreset_in                     : in   std_logic;
    gt7_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt7_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    gt7_rxsyncallin_in                      : in   std_logic;
    gt7_rxsyncdone_out                      : out  std_logic;
    gt7_rxsyncin_in                         : in   std_logic;
    gt7_rxsyncmode_in                       : in   std_logic;
    gt7_rxsyncout_out                       : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt7_rxbyteisaligned_out                 : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt7_rxlpmhfhold_in                      : in   std_logic;
    gt7_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt7_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt7_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt7_rxoutclk_out                        : out  std_logic;
    gt7_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt7_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt7_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt7_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt7_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt7_gttxreset_in                        : in   std_logic;
    gt7_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt7_txusrclk_in                         : in   std_logic;
    gt7_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt7_txdlyen_in                          : in   std_logic;
    gt7_txdlysreset_in                      : in   std_logic;
    gt7_txdlysresetdone_out                 : out  std_logic;
    gt7_txphalign_in                        : in   std_logic;
    gt7_txphaligndone_out                   : out  std_logic;
    gt7_txphalignen_in                      : in   std_logic;
    gt7_txphdlyreset_in                     : in   std_logic;
    gt7_txphinit_in                         : in   std_logic;
    gt7_txphinitdone_out                    : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt7_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt7_gthtxn_out                          : out  std_logic;
    gt7_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt7_txoutclk_out                        : out  std_logic;
    gt7_txoutclkfabric_out                  : out  std_logic;
    gt7_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt7_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt7_txcharisk_in                        : in   std_logic_vector(7 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT8  (X1Y12)
    --____________________________CHANNEL PORTS________________________________
    GT8_DRP_BUSY_OUT                        : out  std_logic;
    GT8_RXPMARESETDONE_OUT                        : out  std_logic;
    GT8_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt8_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt8_drpclk_in                           : in   std_logic;
    gt8_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt8_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt8_drpen_in                            : in   std_logic;
    gt8_drprdy_out                          : out  std_logic;
    gt8_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt8_eyescanreset_in                     : in   std_logic;
    gt8_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt8_eyescandataerror_out                : out  std_logic;
    gt8_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt8_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt8_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt8_rxusrclk_in                         : in   std_logic;
    gt8_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt8_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt8_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt8_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt8_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt8_rxdlyen_in                          : in   std_logic;
    gt8_rxdlysreset_in                      : in   std_logic;
    gt8_rxdlysresetdone_out                 : out  std_logic;
    gt8_rxphalign_in                        : in   std_logic;
    gt8_rxphaligndone_out                   : out  std_logic;
    gt8_rxphalignen_in                      : in   std_logic;
    gt8_rxphdlyreset_in                     : in   std_logic;
    gt8_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt8_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    gt8_rxsyncallin_in                      : in   std_logic;
    gt8_rxsyncdone_out                      : out  std_logic;
    gt8_rxsyncin_in                         : in   std_logic;
    gt8_rxsyncmode_in                       : in   std_logic;
    gt8_rxsyncout_out                       : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt8_rxbyteisaligned_out                 : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt8_rxlpmhfhold_in                      : in   std_logic;
    gt8_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt8_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt8_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt8_rxoutclk_out                        : out  std_logic;
    gt8_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt8_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt8_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt8_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt8_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt8_gttxreset_in                        : in   std_logic;
    gt8_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt8_txusrclk_in                         : in   std_logic;
    gt8_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt8_txdlyen_in                          : in   std_logic;
    gt8_txdlysreset_in                      : in   std_logic;
    gt8_txdlysresetdone_out                 : out  std_logic;
    gt8_txphalign_in                        : in   std_logic;
    gt8_txphaligndone_out                   : out  std_logic;
    gt8_txphalignen_in                      : in   std_logic;
    gt8_txphdlyreset_in                     : in   std_logic;
    gt8_txphinit_in                         : in   std_logic;
    gt8_txphinitdone_out                    : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt8_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt8_gthtxn_out                          : out  std_logic;
    gt8_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt8_txoutclk_out                        : out  std_logic;
    gt8_txoutclkfabric_out                  : out  std_logic;
    gt8_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt8_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt8_txcharisk_in                        : in   std_logic_vector(7 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT9  (X1Y13)
    --____________________________CHANNEL PORTS________________________________
    GT9_DRP_BUSY_OUT                        : out  std_logic;
    GT9_RXPMARESETDONE_OUT                        : out  std_logic;
    GT9_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt9_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt9_drpclk_in                           : in   std_logic;
    gt9_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt9_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt9_drpen_in                            : in   std_logic;
    gt9_drprdy_out                          : out  std_logic;
    gt9_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt9_eyescanreset_in                     : in   std_logic;
    gt9_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt9_eyescandataerror_out                : out  std_logic;
    gt9_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt9_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt9_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt9_rxusrclk_in                         : in   std_logic;
    gt9_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt9_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt9_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt9_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt9_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt9_rxdlyen_in                          : in   std_logic;
    gt9_rxdlysreset_in                      : in   std_logic;
    gt9_rxdlysresetdone_out                 : out  std_logic;
    gt9_rxphalign_in                        : in   std_logic;
    gt9_rxphaligndone_out                   : out  std_logic;
    gt9_rxphalignen_in                      : in   std_logic;
    gt9_rxphdlyreset_in                     : in   std_logic;
    gt9_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt9_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    gt9_rxsyncallin_in                      : in   std_logic;
    gt9_rxsyncdone_out                      : out  std_logic;
    gt9_rxsyncin_in                         : in   std_logic;
    gt9_rxsyncmode_in                       : in   std_logic;
    gt9_rxsyncout_out                       : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt9_rxbyteisaligned_out                 : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt9_rxlpmhfhold_in                      : in   std_logic;
    gt9_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt9_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt9_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt9_rxoutclk_out                        : out  std_logic;
    gt9_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt9_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt9_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt9_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt9_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt9_gttxreset_in                        : in   std_logic;
    gt9_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt9_txusrclk_in                         : in   std_logic;
    gt9_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt9_txdlyen_in                          : in   std_logic;
    gt9_txdlysreset_in                      : in   std_logic;
    gt9_txdlysresetdone_out                 : out  std_logic;
    gt9_txphalign_in                        : in   std_logic;
    gt9_txphaligndone_out                   : out  std_logic;
    gt9_txphalignen_in                      : in   std_logic;
    gt9_txphdlyreset_in                     : in   std_logic;
    gt9_txphinit_in                         : in   std_logic;
    gt9_txphinitdone_out                    : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt9_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt9_gthtxn_out                          : out  std_logic;
    gt9_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt9_txoutclk_out                        : out  std_logic;
    gt9_txoutclkfabric_out                  : out  std_logic;
    gt9_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt9_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt9_txcharisk_in                        : in   std_logic_vector(7 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT10  (X1Y14)
    --____________________________CHANNEL PORTS________________________________
    GT10_DRP_BUSY_OUT                        : out  std_logic;
    GT10_RXPMARESETDONE_OUT                        : out  std_logic;
    GT10_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt10_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt10_drpclk_in                          : in   std_logic;
    gt10_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt10_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt10_drpen_in                           : in   std_logic;
    gt10_drprdy_out                         : out  std_logic;
    gt10_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt10_eyescanreset_in                    : in   std_logic;
    gt10_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt10_eyescandataerror_out               : out  std_logic;
    gt10_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt10_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt10_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt10_rxusrclk_in                        : in   std_logic;
    gt10_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt10_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt10_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt10_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt10_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt10_rxdlyen_in                         : in   std_logic;
    gt10_rxdlysreset_in                     : in   std_logic;
    gt10_rxdlysresetdone_out                : out  std_logic;
    gt10_rxphalign_in                       : in   std_logic;
    gt10_rxphaligndone_out                  : out  std_logic;
    gt10_rxphalignen_in                     : in   std_logic;
    gt10_rxphdlyreset_in                    : in   std_logic;
    gt10_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt10_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt10_rxsyncallin_in                     : in   std_logic;
    gt10_rxsyncdone_out                     : out  std_logic;
    gt10_rxsyncin_in                        : in   std_logic;
    gt10_rxsyncmode_in                      : in   std_logic;
    gt10_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt10_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt10_rxlpmhfhold_in                     : in   std_logic;
    gt10_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt10_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt10_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt10_rxoutclk_out                       : out  std_logic;
    gt10_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt10_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt10_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt10_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt10_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt10_gttxreset_in                       : in   std_logic;
    gt10_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt10_txusrclk_in                        : in   std_logic;
    gt10_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt10_txdlyen_in                         : in   std_logic;
    gt10_txdlysreset_in                     : in   std_logic;
    gt10_txdlysresetdone_out                : out  std_logic;
    gt10_txphalign_in                       : in   std_logic;
    gt10_txphaligndone_out                  : out  std_logic;
    gt10_txphalignen_in                     : in   std_logic;
    gt10_txphdlyreset_in                    : in   std_logic;
    gt10_txphinit_in                        : in   std_logic;
    gt10_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt10_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt10_gthtxn_out                         : out  std_logic;
    gt10_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt10_txoutclk_out                       : out  std_logic;
    gt10_txoutclkfabric_out                 : out  std_logic;
    gt10_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt10_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt10_txcharisk_in                       : in   std_logic_vector(7 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT11  (X1Y15)
    --____________________________CHANNEL PORTS________________________________
    GT11_DRP_BUSY_OUT                        : out  std_logic;
    GT11_RXPMARESETDONE_OUT                        : out  std_logic;
    GT11_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt11_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt11_drpclk_in                          : in   std_logic;
    gt11_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt11_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt11_drpen_in                           : in   std_logic;
    gt11_drprdy_out                         : out  std_logic;
    gt11_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt11_eyescanreset_in                    : in   std_logic;
    gt11_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt11_eyescandataerror_out               : out  std_logic;
    gt11_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt11_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt11_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt11_rxusrclk_in                        : in   std_logic;
    gt11_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt11_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt11_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt11_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt11_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt11_rxdlyen_in                         : in   std_logic;
    gt11_rxdlysreset_in                     : in   std_logic;
    gt11_rxdlysresetdone_out                : out  std_logic;
    gt11_rxphalign_in                       : in   std_logic;
    gt11_rxphaligndone_out                  : out  std_logic;
    gt11_rxphalignen_in                     : in   std_logic;
    gt11_rxphdlyreset_in                    : in   std_logic;
    gt11_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt11_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt11_rxsyncallin_in                     : in   std_logic;
    gt11_rxsyncdone_out                     : out  std_logic;
    gt11_rxsyncin_in                        : in   std_logic;
    gt11_rxsyncmode_in                      : in   std_logic;
    gt11_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt11_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt11_rxlpmhfhold_in                     : in   std_logic;
    gt11_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt11_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt11_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt11_rxoutclk_out                       : out  std_logic;
    gt11_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt11_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt11_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt11_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt11_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt11_gttxreset_in                       : in   std_logic;
    gt11_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt11_txusrclk_in                        : in   std_logic;
    gt11_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt11_txdlyen_in                         : in   std_logic;
    gt11_txdlysreset_in                     : in   std_logic;
    gt11_txdlysresetdone_out                : out  std_logic;
    gt11_txphalign_in                       : in   std_logic;
    gt11_txphaligndone_out                  : out  std_logic;
    gt11_txphalignen_in                     : in   std_logic;
    gt11_txphdlyreset_in                    : in   std_logic;
    gt11_txphinit_in                        : in   std_logic;
    gt11_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt11_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt11_gthtxn_out                         : out  std_logic;
    gt11_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt11_txoutclk_out                       : out  std_logic;
    gt11_txoutclkfabric_out                 : out  std_logic;
    gt11_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt11_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt11_txcharisk_in                       : in   std_logic_vector(7 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT12  (X1Y16)
    --____________________________CHANNEL PORTS________________________________
    GT12_DRP_BUSY_OUT                        : out  std_logic;
    GT12_RXPMARESETDONE_OUT                        : out  std_logic;
    GT12_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt12_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt12_drpclk_in                          : in   std_logic;
    gt12_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt12_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt12_drpen_in                           : in   std_logic;
    gt12_drprdy_out                         : out  std_logic;
    gt12_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt12_eyescanreset_in                    : in   std_logic;
    gt12_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt12_eyescandataerror_out               : out  std_logic;
    gt12_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt12_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt12_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt12_rxusrclk_in                        : in   std_logic;
    gt12_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt12_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt12_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt12_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt12_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt12_rxdlyen_in                         : in   std_logic;
    gt12_rxdlysreset_in                     : in   std_logic;
    gt12_rxdlysresetdone_out                : out  std_logic;
    gt12_rxphalign_in                       : in   std_logic;
    gt12_rxphaligndone_out                  : out  std_logic;
    gt12_rxphalignen_in                     : in   std_logic;
    gt12_rxphdlyreset_in                    : in   std_logic;
    gt12_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt12_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt12_rxsyncallin_in                     : in   std_logic;
    gt12_rxsyncdone_out                     : out  std_logic;
    gt12_rxsyncin_in                        : in   std_logic;
    gt12_rxsyncmode_in                      : in   std_logic;
    gt12_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt12_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt12_rxlpmhfhold_in                     : in   std_logic;
    gt12_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt12_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt12_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt12_rxoutclk_out                       : out  std_logic;
    gt12_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt12_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt12_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt12_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt12_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt12_gttxreset_in                       : in   std_logic;
    gt12_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt12_txusrclk_in                        : in   std_logic;
    gt12_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt12_txdlyen_in                         : in   std_logic;
    gt12_txdlysreset_in                     : in   std_logic;
    gt12_txdlysresetdone_out                : out  std_logic;
    gt12_txphalign_in                       : in   std_logic;
    gt12_txphaligndone_out                  : out  std_logic;
    gt12_txphalignen_in                     : in   std_logic;
    gt12_txphdlyreset_in                    : in   std_logic;
    gt12_txphinit_in                        : in   std_logic;
    gt12_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt12_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt12_gthtxn_out                         : out  std_logic;
    gt12_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt12_txoutclk_out                       : out  std_logic;
    gt12_txoutclkfabric_out                 : out  std_logic;
    gt12_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt12_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt12_txcharisk_in                       : in   std_logic_vector(7 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT13  (X1Y17)
    --____________________________CHANNEL PORTS________________________________
    GT13_DRP_BUSY_OUT                        : out  std_logic;
    GT13_RXPMARESETDONE_OUT                        : out  std_logic;
    GT13_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt13_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt13_drpclk_in                          : in   std_logic;
    gt13_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt13_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt13_drpen_in                           : in   std_logic;
    gt13_drprdy_out                         : out  std_logic;
    gt13_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt13_eyescanreset_in                    : in   std_logic;
    gt13_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt13_eyescandataerror_out               : out  std_logic;
    gt13_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt13_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt13_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt13_rxusrclk_in                        : in   std_logic;
    gt13_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt13_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt13_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt13_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt13_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt13_rxdlyen_in                         : in   std_logic;
    gt13_rxdlysreset_in                     : in   std_logic;
    gt13_rxdlysresetdone_out                : out  std_logic;
    gt13_rxphalign_in                       : in   std_logic;
    gt13_rxphaligndone_out                  : out  std_logic;
    gt13_rxphalignen_in                     : in   std_logic;
    gt13_rxphdlyreset_in                    : in   std_logic;
    gt13_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt13_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt13_rxsyncallin_in                     : in   std_logic;
    gt13_rxsyncdone_out                     : out  std_logic;
    gt13_rxsyncin_in                        : in   std_logic;
    gt13_rxsyncmode_in                      : in   std_logic;
    gt13_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt13_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt13_rxlpmhfhold_in                     : in   std_logic;
    gt13_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt13_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt13_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt13_rxoutclk_out                       : out  std_logic;
    gt13_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt13_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt13_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt13_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt13_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt13_gttxreset_in                       : in   std_logic;
    gt13_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt13_txusrclk_in                        : in   std_logic;
    gt13_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt13_txdlyen_in                         : in   std_logic;
    gt13_txdlysreset_in                     : in   std_logic;
    gt13_txdlysresetdone_out                : out  std_logic;
    gt13_txphalign_in                       : in   std_logic;
    gt13_txphaligndone_out                  : out  std_logic;
    gt13_txphalignen_in                     : in   std_logic;
    gt13_txphdlyreset_in                    : in   std_logic;
    gt13_txphinit_in                        : in   std_logic;
    gt13_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt13_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt13_gthtxn_out                         : out  std_logic;
    gt13_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt13_txoutclk_out                       : out  std_logic;
    gt13_txoutclkfabric_out                 : out  std_logic;
    gt13_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt13_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt13_txcharisk_in                       : in   std_logic_vector(7 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT14  (X1Y18)
    --____________________________CHANNEL PORTS________________________________
    GT14_DRP_BUSY_OUT                        : out  std_logic;
    GT14_RXPMARESETDONE_OUT                        : out  std_logic;
    GT14_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt14_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt14_drpclk_in                          : in   std_logic;
    gt14_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt14_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt14_drpen_in                           : in   std_logic;
    gt14_drprdy_out                         : out  std_logic;
    gt14_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt14_eyescanreset_in                    : in   std_logic;
    gt14_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt14_eyescandataerror_out               : out  std_logic;
    gt14_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt14_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt14_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt14_rxusrclk_in                        : in   std_logic;
    gt14_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt14_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt14_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt14_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt14_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt14_rxdlyen_in                         : in   std_logic;
    gt14_rxdlysreset_in                     : in   std_logic;
    gt14_rxdlysresetdone_out                : out  std_logic;
    gt14_rxphalign_in                       : in   std_logic;
    gt14_rxphaligndone_out                  : out  std_logic;
    gt14_rxphalignen_in                     : in   std_logic;
    gt14_rxphdlyreset_in                    : in   std_logic;
    gt14_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt14_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt14_rxsyncallin_in                     : in   std_logic;
    gt14_rxsyncdone_out                     : out  std_logic;
    gt14_rxsyncin_in                        : in   std_logic;
    gt14_rxsyncmode_in                      : in   std_logic;
    gt14_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt14_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt14_rxlpmhfhold_in                     : in   std_logic;
    gt14_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt14_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt14_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt14_rxoutclk_out                       : out  std_logic;
    gt14_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt14_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt14_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt14_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt14_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt14_gttxreset_in                       : in   std_logic;
    gt14_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt14_txusrclk_in                        : in   std_logic;
    gt14_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt14_txdlyen_in                         : in   std_logic;
    gt14_txdlysreset_in                     : in   std_logic;
    gt14_txdlysresetdone_out                : out  std_logic;
    gt14_txphalign_in                       : in   std_logic;
    gt14_txphaligndone_out                  : out  std_logic;
    gt14_txphalignen_in                     : in   std_logic;
    gt14_txphdlyreset_in                    : in   std_logic;
    gt14_txphinit_in                        : in   std_logic;
    gt14_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt14_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt14_gthtxn_out                         : out  std_logic;
    gt14_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt14_txoutclk_out                       : out  std_logic;
    gt14_txoutclkfabric_out                 : out  std_logic;
    gt14_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt14_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt14_txcharisk_in                       : in   std_logic_vector(7 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT15  (X1Y19)
    --____________________________CHANNEL PORTS________________________________
    GT15_DRP_BUSY_OUT                        : out  std_logic;
    GT15_RXPMARESETDONE_OUT                        : out  std_logic;
    GT15_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt15_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt15_drpclk_in                          : in   std_logic;
    gt15_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt15_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt15_drpen_in                           : in   std_logic;
    gt15_drprdy_out                         : out  std_logic;
    gt15_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt15_eyescanreset_in                    : in   std_logic;
    gt15_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt15_eyescandataerror_out               : out  std_logic;
    gt15_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt15_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt15_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt15_rxusrclk_in                        : in   std_logic;
    gt15_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt15_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt15_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt15_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt15_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt15_rxdlyen_in                         : in   std_logic;
    gt15_rxdlysreset_in                     : in   std_logic;
    gt15_rxdlysresetdone_out                : out  std_logic;
    gt15_rxphalign_in                       : in   std_logic;
    gt15_rxphaligndone_out                  : out  std_logic;
    gt15_rxphalignen_in                     : in   std_logic;
    gt15_rxphdlyreset_in                    : in   std_logic;
    gt15_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt15_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt15_rxsyncallin_in                     : in   std_logic;
    gt15_rxsyncdone_out                     : out  std_logic;
    gt15_rxsyncin_in                        : in   std_logic;
    gt15_rxsyncmode_in                      : in   std_logic;
    gt15_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt15_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt15_rxlpmhfhold_in                     : in   std_logic;
    gt15_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt15_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt15_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt15_rxoutclk_out                       : out  std_logic;
    gt15_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt15_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt15_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt15_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt15_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt15_gttxreset_in                       : in   std_logic;
    gt15_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt15_txusrclk_in                        : in   std_logic;
    gt15_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt15_txdlyen_in                         : in   std_logic;
    gt15_txdlysreset_in                     : in   std_logic;
    gt15_txdlysresetdone_out                : out  std_logic;
    gt15_txphalign_in                       : in   std_logic;
    gt15_txphaligndone_out                  : out  std_logic;
    gt15_txphalignen_in                     : in   std_logic;
    gt15_txphdlyreset_in                    : in   std_logic;
    gt15_txphinit_in                        : in   std_logic;
    gt15_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt15_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt15_gthtxn_out                         : out  std_logic;
    gt15_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt15_txoutclk_out                       : out  std_logic;
    gt15_txoutclkfabric_out                 : out  std_logic;
    gt15_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt15_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt15_txcharisk_in                       : in   std_logic_vector(7 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT16  (X1Y20)
    --____________________________CHANNEL PORTS________________________________
    GT16_DRP_BUSY_OUT                        : out  std_logic;
    GT16_RXPMARESETDONE_OUT                        : out  std_logic;
    GT16_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt16_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt16_drpclk_in                          : in   std_logic;
    gt16_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt16_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt16_drpen_in                           : in   std_logic;
    gt16_drprdy_out                         : out  std_logic;
    gt16_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt16_eyescanreset_in                    : in   std_logic;
    gt16_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt16_eyescandataerror_out               : out  std_logic;
    gt16_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt16_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt16_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt16_rxusrclk_in                        : in   std_logic;
    gt16_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt16_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt16_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt16_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt16_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt16_rxdlyen_in                         : in   std_logic;
    gt16_rxdlysreset_in                     : in   std_logic;
    gt16_rxdlysresetdone_out                : out  std_logic;
    gt16_rxphalign_in                       : in   std_logic;
    gt16_rxphaligndone_out                  : out  std_logic;
    gt16_rxphalignen_in                     : in   std_logic;
    gt16_rxphdlyreset_in                    : in   std_logic;
    gt16_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt16_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt16_rxsyncallin_in                     : in   std_logic;
    gt16_rxsyncdone_out                     : out  std_logic;
    gt16_rxsyncin_in                        : in   std_logic;
    gt16_rxsyncmode_in                      : in   std_logic;
    gt16_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt16_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt16_rxlpmhfhold_in                     : in   std_logic;
    gt16_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt16_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt16_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt16_rxoutclk_out                       : out  std_logic;
    gt16_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt16_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt16_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt16_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt16_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt16_gttxreset_in                       : in   std_logic;
    gt16_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt16_txusrclk_in                        : in   std_logic;
    gt16_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt16_txdlyen_in                         : in   std_logic;
    gt16_txdlysreset_in                     : in   std_logic;
    gt16_txdlysresetdone_out                : out  std_logic;
    gt16_txphalign_in                       : in   std_logic;
    gt16_txphaligndone_out                  : out  std_logic;
    gt16_txphalignen_in                     : in   std_logic;
    gt16_txphdlyreset_in                    : in   std_logic;
    gt16_txphinit_in                        : in   std_logic;
    gt16_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt16_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt16_gthtxn_out                         : out  std_logic;
    gt16_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt16_txoutclk_out                       : out  std_logic;
    gt16_txoutclkfabric_out                 : out  std_logic;
    gt16_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt16_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt16_txcharisk_in                       : in   std_logic_vector(7 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT17  (X1Y21)
    --____________________________CHANNEL PORTS________________________________
    GT17_DRP_BUSY_OUT                        : out  std_logic;
    GT17_RXPMARESETDONE_OUT                        : out  std_logic;
    GT17_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt17_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt17_drpclk_in                          : in   std_logic;
    gt17_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt17_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt17_drpen_in                           : in   std_logic;
    gt17_drprdy_out                         : out  std_logic;
    gt17_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt17_eyescanreset_in                    : in   std_logic;
    gt17_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt17_eyescandataerror_out               : out  std_logic;
    gt17_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt17_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt17_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt17_rxusrclk_in                        : in   std_logic;
    gt17_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt17_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt17_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt17_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt17_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt17_rxdlyen_in                         : in   std_logic;
    gt17_rxdlysreset_in                     : in   std_logic;
    gt17_rxdlysresetdone_out                : out  std_logic;
    gt17_rxphalign_in                       : in   std_logic;
    gt17_rxphaligndone_out                  : out  std_logic;
    gt17_rxphalignen_in                     : in   std_logic;
    gt17_rxphdlyreset_in                    : in   std_logic;
    gt17_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt17_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt17_rxsyncallin_in                     : in   std_logic;
    gt17_rxsyncdone_out                     : out  std_logic;
    gt17_rxsyncin_in                        : in   std_logic;
    gt17_rxsyncmode_in                      : in   std_logic;
    gt17_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt17_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt17_rxlpmhfhold_in                     : in   std_logic;
    gt17_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt17_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt17_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt17_rxoutclk_out                       : out  std_logic;
    gt17_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt17_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt17_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt17_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt17_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt17_gttxreset_in                       : in   std_logic;
    gt17_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt17_txusrclk_in                        : in   std_logic;
    gt17_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt17_txdlyen_in                         : in   std_logic;
    gt17_txdlysreset_in                     : in   std_logic;
    gt17_txdlysresetdone_out                : out  std_logic;
    gt17_txphalign_in                       : in   std_logic;
    gt17_txphaligndone_out                  : out  std_logic;
    gt17_txphalignen_in                     : in   std_logic;
    gt17_txphdlyreset_in                    : in   std_logic;
    gt17_txphinit_in                        : in   std_logic;
    gt17_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt17_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt17_gthtxn_out                         : out  std_logic;
    gt17_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt17_txoutclk_out                       : out  std_logic;
    gt17_txoutclkfabric_out                 : out  std_logic;
    gt17_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt17_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt17_txcharisk_in                       : in   std_logic_vector(7 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT18  (X1Y22)
    --____________________________CHANNEL PORTS________________________________
    GT18_DRP_BUSY_OUT                        : out  std_logic;
    GT18_RXPMARESETDONE_OUT                        : out  std_logic;
    GT18_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt18_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt18_drpclk_in                          : in   std_logic;
    gt18_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt18_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt18_drpen_in                           : in   std_logic;
    gt18_drprdy_out                         : out  std_logic;
    gt18_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt18_eyescanreset_in                    : in   std_logic;
    gt18_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt18_eyescandataerror_out               : out  std_logic;
    gt18_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt18_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt18_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt18_rxusrclk_in                        : in   std_logic;
    gt18_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt18_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt18_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt18_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt18_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt18_rxdlyen_in                         : in   std_logic;
    gt18_rxdlysreset_in                     : in   std_logic;
    gt18_rxdlysresetdone_out                : out  std_logic;
    gt18_rxphalign_in                       : in   std_logic;
    gt18_rxphaligndone_out                  : out  std_logic;
    gt18_rxphalignen_in                     : in   std_logic;
    gt18_rxphdlyreset_in                    : in   std_logic;
    gt18_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt18_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt18_rxsyncallin_in                     : in   std_logic;
    gt18_rxsyncdone_out                     : out  std_logic;
    gt18_rxsyncin_in                        : in   std_logic;
    gt18_rxsyncmode_in                      : in   std_logic;
    gt18_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt18_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt18_rxlpmhfhold_in                     : in   std_logic;
    gt18_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt18_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt18_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt18_rxoutclk_out                       : out  std_logic;
    gt18_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt18_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt18_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt18_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt18_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt18_gttxreset_in                       : in   std_logic;
    gt18_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt18_txusrclk_in                        : in   std_logic;
    gt18_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt18_txdlyen_in                         : in   std_logic;
    gt18_txdlysreset_in                     : in   std_logic;
    gt18_txdlysresetdone_out                : out  std_logic;
    gt18_txphalign_in                       : in   std_logic;
    gt18_txphaligndone_out                  : out  std_logic;
    gt18_txphalignen_in                     : in   std_logic;
    gt18_txphdlyreset_in                    : in   std_logic;
    gt18_txphinit_in                        : in   std_logic;
    gt18_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt18_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt18_gthtxn_out                         : out  std_logic;
    gt18_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt18_txoutclk_out                       : out  std_logic;
    gt18_txoutclkfabric_out                 : out  std_logic;
    gt18_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt18_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt18_txcharisk_in                       : in   std_logic_vector(7 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT19  (X1Y23)
    --____________________________CHANNEL PORTS________________________________
    GT19_DRP_BUSY_OUT                        : out  std_logic;
    GT19_RXPMARESETDONE_OUT                        : out  std_logic;
    GT19_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt19_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt19_drpclk_in                          : in   std_logic;
    gt19_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt19_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt19_drpen_in                           : in   std_logic;
    gt19_drprdy_out                         : out  std_logic;
    gt19_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt19_eyescanreset_in                    : in   std_logic;
    gt19_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt19_eyescandataerror_out               : out  std_logic;
    gt19_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt19_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt19_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt19_rxusrclk_in                        : in   std_logic;
    gt19_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt19_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt19_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt19_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt19_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt19_rxdlyen_in                         : in   std_logic;
    gt19_rxdlysreset_in                     : in   std_logic;
    gt19_rxdlysresetdone_out                : out  std_logic;
    gt19_rxphalign_in                       : in   std_logic;
    gt19_rxphaligndone_out                  : out  std_logic;
    gt19_rxphalignen_in                     : in   std_logic;
    gt19_rxphdlyreset_in                    : in   std_logic;
    gt19_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt19_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt19_rxsyncallin_in                     : in   std_logic;
    gt19_rxsyncdone_out                     : out  std_logic;
    gt19_rxsyncin_in                        : in   std_logic;
    gt19_rxsyncmode_in                      : in   std_logic;
    gt19_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt19_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt19_rxlpmhfhold_in                     : in   std_logic;
    gt19_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt19_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt19_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt19_rxoutclk_out                       : out  std_logic;
    gt19_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt19_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt19_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt19_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt19_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt19_gttxreset_in                       : in   std_logic;
    gt19_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt19_txusrclk_in                        : in   std_logic;
    gt19_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt19_txdlyen_in                         : in   std_logic;
    gt19_txdlysreset_in                     : in   std_logic;
    gt19_txdlysresetdone_out                : out  std_logic;
    gt19_txphalign_in                       : in   std_logic;
    gt19_txphaligndone_out                  : out  std_logic;
    gt19_txphalignen_in                     : in   std_logic;
    gt19_txphdlyreset_in                    : in   std_logic;
    gt19_txphinit_in                        : in   std_logic;
    gt19_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt19_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt19_gthtxn_out                         : out  std_logic;
    gt19_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt19_txoutclk_out                       : out  std_logic;
    gt19_txoutclkfabric_out                 : out  std_logic;
    gt19_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt19_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt19_txcharisk_in                       : in   std_logic_vector(7 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT20  (X1Y24)
    --____________________________CHANNEL PORTS________________________________
    GT20_DRP_BUSY_OUT                        : out  std_logic;
    GT20_RXPMARESETDONE_OUT                        : out  std_logic;
    GT20_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt20_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt20_drpclk_in                          : in   std_logic;
    gt20_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt20_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt20_drpen_in                           : in   std_logic;
    gt20_drprdy_out                         : out  std_logic;
    gt20_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt20_eyescanreset_in                    : in   std_logic;
    gt20_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt20_eyescandataerror_out               : out  std_logic;
    gt20_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt20_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt20_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt20_rxusrclk_in                        : in   std_logic;
    gt20_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt20_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt20_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt20_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt20_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt20_rxdlyen_in                         : in   std_logic;
    gt20_rxdlysreset_in                     : in   std_logic;
    gt20_rxdlysresetdone_out                : out  std_logic;
    gt20_rxphalign_in                       : in   std_logic;
    gt20_rxphaligndone_out                  : out  std_logic;
    gt20_rxphalignen_in                     : in   std_logic;
    gt20_rxphdlyreset_in                    : in   std_logic;
    gt20_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt20_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt20_rxsyncallin_in                     : in   std_logic;
    gt20_rxsyncdone_out                     : out  std_logic;
    gt20_rxsyncin_in                        : in   std_logic;
    gt20_rxsyncmode_in                      : in   std_logic;
    gt20_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt20_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt20_rxlpmhfhold_in                     : in   std_logic;
    gt20_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt20_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt20_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt20_rxoutclk_out                       : out  std_logic;
    gt20_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt20_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt20_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt20_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt20_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt20_gttxreset_in                       : in   std_logic;
    gt20_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt20_txusrclk_in                        : in   std_logic;
    gt20_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt20_txdlyen_in                         : in   std_logic;
    gt20_txdlysreset_in                     : in   std_logic;
    gt20_txdlysresetdone_out                : out  std_logic;
    gt20_txphalign_in                       : in   std_logic;
    gt20_txphaligndone_out                  : out  std_logic;
    gt20_txphalignen_in                     : in   std_logic;
    gt20_txphdlyreset_in                    : in   std_logic;
    gt20_txphinit_in                        : in   std_logic;
    gt20_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt20_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt20_gthtxn_out                         : out  std_logic;
    gt20_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt20_txoutclk_out                       : out  std_logic;
    gt20_txoutclkfabric_out                 : out  std_logic;
    gt20_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt20_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt20_txcharisk_in                       : in   std_logic_vector(7 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT21  (X1Y25)
    --____________________________CHANNEL PORTS________________________________
    GT21_DRP_BUSY_OUT                        : out  std_logic;
    GT21_RXPMARESETDONE_OUT                        : out  std_logic;
    GT21_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt21_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt21_drpclk_in                          : in   std_logic;
    gt21_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt21_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt21_drpen_in                           : in   std_logic;
    gt21_drprdy_out                         : out  std_logic;
    gt21_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt21_eyescanreset_in                    : in   std_logic;
    gt21_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt21_eyescandataerror_out               : out  std_logic;
    gt21_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt21_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt21_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt21_rxusrclk_in                        : in   std_logic;
    gt21_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt21_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt21_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt21_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt21_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt21_rxdlyen_in                         : in   std_logic;
    gt21_rxdlysreset_in                     : in   std_logic;
    gt21_rxdlysresetdone_out                : out  std_logic;
    gt21_rxphalign_in                       : in   std_logic;
    gt21_rxphaligndone_out                  : out  std_logic;
    gt21_rxphalignen_in                     : in   std_logic;
    gt21_rxphdlyreset_in                    : in   std_logic;
    gt21_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt21_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt21_rxsyncallin_in                     : in   std_logic;
    gt21_rxsyncdone_out                     : out  std_logic;
    gt21_rxsyncin_in                        : in   std_logic;
    gt21_rxsyncmode_in                      : in   std_logic;
    gt21_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt21_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt21_rxlpmhfhold_in                     : in   std_logic;
    gt21_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt21_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt21_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt21_rxoutclk_out                       : out  std_logic;
    gt21_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt21_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt21_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt21_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt21_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt21_gttxreset_in                       : in   std_logic;
    gt21_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt21_txusrclk_in                        : in   std_logic;
    gt21_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt21_txdlyen_in                         : in   std_logic;
    gt21_txdlysreset_in                     : in   std_logic;
    gt21_txdlysresetdone_out                : out  std_logic;
    gt21_txphalign_in                       : in   std_logic;
    gt21_txphaligndone_out                  : out  std_logic;
    gt21_txphalignen_in                     : in   std_logic;
    gt21_txphdlyreset_in                    : in   std_logic;
    gt21_txphinit_in                        : in   std_logic;
    gt21_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt21_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt21_gthtxn_out                         : out  std_logic;
    gt21_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt21_txoutclk_out                       : out  std_logic;
    gt21_txoutclkfabric_out                 : out  std_logic;
    gt21_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt21_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt21_txcharisk_in                       : in   std_logic_vector(7 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT22  (X1Y26)
    --____________________________CHANNEL PORTS________________________________
    GT22_DRP_BUSY_OUT                        : out  std_logic;
    GT22_RXPMARESETDONE_OUT                        : out  std_logic;
    GT22_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt22_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt22_drpclk_in                          : in   std_logic;
    gt22_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt22_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt22_drpen_in                           : in   std_logic;
    gt22_drprdy_out                         : out  std_logic;
    gt22_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt22_eyescanreset_in                    : in   std_logic;
    gt22_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt22_eyescandataerror_out               : out  std_logic;
    gt22_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt22_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt22_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt22_rxusrclk_in                        : in   std_logic;
    gt22_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt22_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt22_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt22_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt22_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt22_rxdlyen_in                         : in   std_logic;
    gt22_rxdlysreset_in                     : in   std_logic;
    gt22_rxdlysresetdone_out                : out  std_logic;
    gt22_rxphalign_in                       : in   std_logic;
    gt22_rxphaligndone_out                  : out  std_logic;
    gt22_rxphalignen_in                     : in   std_logic;
    gt22_rxphdlyreset_in                    : in   std_logic;
    gt22_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt22_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt22_rxsyncallin_in                     : in   std_logic;
    gt22_rxsyncdone_out                     : out  std_logic;
    gt22_rxsyncin_in                        : in   std_logic;
    gt22_rxsyncmode_in                      : in   std_logic;
    gt22_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt22_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt22_rxlpmhfhold_in                     : in   std_logic;
    gt22_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt22_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt22_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt22_rxoutclk_out                       : out  std_logic;
    gt22_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt22_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt22_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt22_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt22_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt22_gttxreset_in                       : in   std_logic;
    gt22_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt22_txusrclk_in                        : in   std_logic;
    gt22_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt22_txdlyen_in                         : in   std_logic;
    gt22_txdlysreset_in                     : in   std_logic;
    gt22_txdlysresetdone_out                : out  std_logic;
    gt22_txphalign_in                       : in   std_logic;
    gt22_txphaligndone_out                  : out  std_logic;
    gt22_txphalignen_in                     : in   std_logic;
    gt22_txphdlyreset_in                    : in   std_logic;
    gt22_txphinit_in                        : in   std_logic;
    gt22_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt22_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt22_gthtxn_out                         : out  std_logic;
    gt22_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt22_txoutclk_out                       : out  std_logic;
    gt22_txoutclkfabric_out                 : out  std_logic;
    gt22_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt22_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt22_txcharisk_in                       : in   std_logic_vector(7 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT23  (X1Y27)
    --____________________________CHANNEL PORTS________________________________
    GT23_DRP_BUSY_OUT                        : out  std_logic;
    GT23_RXPMARESETDONE_OUT                        : out  std_logic;
    GT23_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt23_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt23_drpclk_in                          : in   std_logic;
    gt23_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt23_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt23_drpen_in                           : in   std_logic;
    gt23_drprdy_out                         : out  std_logic;
    gt23_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt23_eyescanreset_in                    : in   std_logic;
    gt23_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt23_eyescandataerror_out               : out  std_logic;
    gt23_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt23_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt23_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt23_rxusrclk_in                        : in   std_logic;
    gt23_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt23_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt23_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt23_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt23_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt23_rxdlyen_in                         : in   std_logic;
    gt23_rxdlysreset_in                     : in   std_logic;
    gt23_rxdlysresetdone_out                : out  std_logic;
    gt23_rxphalign_in                       : in   std_logic;
    gt23_rxphaligndone_out                  : out  std_logic;
    gt23_rxphalignen_in                     : in   std_logic;
    gt23_rxphdlyreset_in                    : in   std_logic;
    gt23_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt23_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt23_rxsyncallin_in                     : in   std_logic;
    gt23_rxsyncdone_out                     : out  std_logic;
    gt23_rxsyncin_in                        : in   std_logic;
    gt23_rxsyncmode_in                      : in   std_logic;
    gt23_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt23_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt23_rxlpmhfhold_in                     : in   std_logic;
    gt23_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt23_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt23_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt23_rxoutclk_out                       : out  std_logic;
    gt23_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt23_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt23_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt23_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt23_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt23_gttxreset_in                       : in   std_logic;
    gt23_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt23_txusrclk_in                        : in   std_logic;
    gt23_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt23_txdlyen_in                         : in   std_logic;
    gt23_txdlysreset_in                     : in   std_logic;
    gt23_txdlysresetdone_out                : out  std_logic;
    gt23_txphalign_in                       : in   std_logic;
    gt23_txphaligndone_out                  : out  std_logic;
    gt23_txphalignen_in                     : in   std_logic;
    gt23_txphdlyreset_in                    : in   std_logic;
    gt23_txphinit_in                        : in   std_logic;
    gt23_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt23_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt23_gthtxn_out                         : out  std_logic;
    gt23_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt23_txoutclk_out                       : out  std_logic;
    gt23_txoutclkfabric_out                 : out  std_logic;
    gt23_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt23_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt23_txcharisk_in                       : in   std_logic_vector(7 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT24  (X1Y28)
    --____________________________CHANNEL PORTS________________________________
    GT24_DRP_BUSY_OUT                        : out  std_logic;
    GT24_RXPMARESETDONE_OUT                        : out  std_logic;
    GT24_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt24_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt24_drpclk_in                          : in   std_logic;
    gt24_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt24_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt24_drpen_in                           : in   std_logic;
    gt24_drprdy_out                         : out  std_logic;
    gt24_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt24_eyescanreset_in                    : in   std_logic;
    gt24_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt24_eyescandataerror_out               : out  std_logic;
    gt24_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt24_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt24_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt24_rxusrclk_in                        : in   std_logic;
    gt24_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt24_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt24_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt24_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt24_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt24_rxdlyen_in                         : in   std_logic;
    gt24_rxdlysreset_in                     : in   std_logic;
    gt24_rxdlysresetdone_out                : out  std_logic;
    gt24_rxphalign_in                       : in   std_logic;
    gt24_rxphaligndone_out                  : out  std_logic;
    gt24_rxphalignen_in                     : in   std_logic;
    gt24_rxphdlyreset_in                    : in   std_logic;
    gt24_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt24_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt24_rxsyncallin_in                     : in   std_logic;
    gt24_rxsyncdone_out                     : out  std_logic;
    gt24_rxsyncin_in                        : in   std_logic;
    gt24_rxsyncmode_in                      : in   std_logic;
    gt24_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt24_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt24_rxlpmhfhold_in                     : in   std_logic;
    gt24_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt24_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt24_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt24_rxoutclk_out                       : out  std_logic;
    gt24_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt24_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt24_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt24_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt24_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt24_gttxreset_in                       : in   std_logic;
    gt24_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt24_txusrclk_in                        : in   std_logic;
    gt24_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt24_txdlyen_in                         : in   std_logic;
    gt24_txdlysreset_in                     : in   std_logic;
    gt24_txdlysresetdone_out                : out  std_logic;
    gt24_txphalign_in                       : in   std_logic;
    gt24_txphaligndone_out                  : out  std_logic;
    gt24_txphalignen_in                     : in   std_logic;
    gt24_txphdlyreset_in                    : in   std_logic;
    gt24_txphinit_in                        : in   std_logic;
    gt24_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt24_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt24_gthtxn_out                         : out  std_logic;
    gt24_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt24_txoutclk_out                       : out  std_logic;
    gt24_txoutclkfabric_out                 : out  std_logic;
    gt24_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt24_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt24_txcharisk_in                       : in   std_logic_vector(7 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT25  (X1Y29)
    --____________________________CHANNEL PORTS________________________________
    GT25_DRP_BUSY_OUT                        : out  std_logic;
    GT25_RXPMARESETDONE_OUT                        : out  std_logic;
    GT25_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt25_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt25_drpclk_in                          : in   std_logic;
    gt25_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt25_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt25_drpen_in                           : in   std_logic;
    gt25_drprdy_out                         : out  std_logic;
    gt25_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt25_eyescanreset_in                    : in   std_logic;
    gt25_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt25_eyescandataerror_out               : out  std_logic;
    gt25_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt25_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt25_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt25_rxusrclk_in                        : in   std_logic;
    gt25_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt25_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt25_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt25_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt25_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt25_rxdlyen_in                         : in   std_logic;
    gt25_rxdlysreset_in                     : in   std_logic;
    gt25_rxdlysresetdone_out                : out  std_logic;
    gt25_rxphalign_in                       : in   std_logic;
    gt25_rxphaligndone_out                  : out  std_logic;
    gt25_rxphalignen_in                     : in   std_logic;
    gt25_rxphdlyreset_in                    : in   std_logic;
    gt25_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt25_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt25_rxsyncallin_in                     : in   std_logic;
    gt25_rxsyncdone_out                     : out  std_logic;
    gt25_rxsyncin_in                        : in   std_logic;
    gt25_rxsyncmode_in                      : in   std_logic;
    gt25_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt25_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt25_rxlpmhfhold_in                     : in   std_logic;
    gt25_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt25_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt25_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt25_rxoutclk_out                       : out  std_logic;
    gt25_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt25_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt25_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt25_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt25_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt25_gttxreset_in                       : in   std_logic;
    gt25_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt25_txusrclk_in                        : in   std_logic;
    gt25_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt25_txdlyen_in                         : in   std_logic;
    gt25_txdlysreset_in                     : in   std_logic;
    gt25_txdlysresetdone_out                : out  std_logic;
    gt25_txphalign_in                       : in   std_logic;
    gt25_txphaligndone_out                  : out  std_logic;
    gt25_txphalignen_in                     : in   std_logic;
    gt25_txphdlyreset_in                    : in   std_logic;
    gt25_txphinit_in                        : in   std_logic;
    gt25_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt25_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt25_gthtxn_out                         : out  std_logic;
    gt25_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt25_txoutclk_out                       : out  std_logic;
    gt25_txoutclkfabric_out                 : out  std_logic;
    gt25_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt25_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt25_txcharisk_in                       : in   std_logic_vector(7 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT26  (X1Y30)
    --____________________________CHANNEL PORTS________________________________
    GT26_DRP_BUSY_OUT                        : out  std_logic;
    GT26_RXPMARESETDONE_OUT                        : out  std_logic;
    GT26_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt26_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt26_drpclk_in                          : in   std_logic;
    gt26_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt26_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt26_drpen_in                           : in   std_logic;
    gt26_drprdy_out                         : out  std_logic;
    gt26_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt26_eyescanreset_in                    : in   std_logic;
    gt26_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt26_eyescandataerror_out               : out  std_logic;
    gt26_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt26_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt26_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt26_rxusrclk_in                        : in   std_logic;
    gt26_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt26_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt26_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt26_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt26_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt26_rxdlyen_in                         : in   std_logic;
    gt26_rxdlysreset_in                     : in   std_logic;
    gt26_rxdlysresetdone_out                : out  std_logic;
    gt26_rxphalign_in                       : in   std_logic;
    gt26_rxphaligndone_out                  : out  std_logic;
    gt26_rxphalignen_in                     : in   std_logic;
    gt26_rxphdlyreset_in                    : in   std_logic;
    gt26_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt26_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt26_rxsyncallin_in                     : in   std_logic;
    gt26_rxsyncdone_out                     : out  std_logic;
    gt26_rxsyncin_in                        : in   std_logic;
    gt26_rxsyncmode_in                      : in   std_logic;
    gt26_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt26_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt26_rxlpmhfhold_in                     : in   std_logic;
    gt26_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt26_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt26_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt26_rxoutclk_out                       : out  std_logic;
    gt26_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt26_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt26_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt26_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt26_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt26_gttxreset_in                       : in   std_logic;
    gt26_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt26_txusrclk_in                        : in   std_logic;
    gt26_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt26_txdlyen_in                         : in   std_logic;
    gt26_txdlysreset_in                     : in   std_logic;
    gt26_txdlysresetdone_out                : out  std_logic;
    gt26_txphalign_in                       : in   std_logic;
    gt26_txphaligndone_out                  : out  std_logic;
    gt26_txphalignen_in                     : in   std_logic;
    gt26_txphdlyreset_in                    : in   std_logic;
    gt26_txphinit_in                        : in   std_logic;
    gt26_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt26_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt26_gthtxn_out                         : out  std_logic;
    gt26_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt26_txoutclk_out                       : out  std_logic;
    gt26_txoutclkfabric_out                 : out  std_logic;
    gt26_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt26_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt26_txcharisk_in                       : in   std_logic_vector(7 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT27  (X1Y31)
    --____________________________CHANNEL PORTS________________________________
    GT27_DRP_BUSY_OUT                        : out  std_logic;
    GT27_RXPMARESETDONE_OUT                        : out  std_logic;
    GT27_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt27_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt27_drpclk_in                          : in   std_logic;
    gt27_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt27_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt27_drpen_in                           : in   std_logic;
    gt27_drprdy_out                         : out  std_logic;
    gt27_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt27_eyescanreset_in                    : in   std_logic;
    gt27_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt27_eyescandataerror_out               : out  std_logic;
    gt27_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt27_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt27_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt27_rxusrclk_in                        : in   std_logic;
    gt27_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt27_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt27_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt27_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt27_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt27_rxdlyen_in                         : in   std_logic;
    gt27_rxdlysreset_in                     : in   std_logic;
    gt27_rxdlysresetdone_out                : out  std_logic;
    gt27_rxphalign_in                       : in   std_logic;
    gt27_rxphaligndone_out                  : out  std_logic;
    gt27_rxphalignen_in                     : in   std_logic;
    gt27_rxphdlyreset_in                    : in   std_logic;
    gt27_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt27_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt27_rxsyncallin_in                     : in   std_logic;
    gt27_rxsyncdone_out                     : out  std_logic;
    gt27_rxsyncin_in                        : in   std_logic;
    gt27_rxsyncmode_in                      : in   std_logic;
    gt27_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt27_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt27_rxlpmhfhold_in                     : in   std_logic;
    gt27_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt27_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt27_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt27_rxoutclk_out                       : out  std_logic;
    gt27_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt27_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt27_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt27_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt27_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt27_gttxreset_in                       : in   std_logic;
    gt27_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt27_txusrclk_in                        : in   std_logic;
    gt27_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt27_txdlyen_in                         : in   std_logic;
    gt27_txdlysreset_in                     : in   std_logic;
    gt27_txdlysresetdone_out                : out  std_logic;
    gt27_txphalign_in                       : in   std_logic;
    gt27_txphaligndone_out                  : out  std_logic;
    gt27_txphalignen_in                     : in   std_logic;
    gt27_txphdlyreset_in                    : in   std_logic;
    gt27_txphinit_in                        : in   std_logic;
    gt27_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt27_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt27_gthtxn_out                         : out  std_logic;
    gt27_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt27_txoutclk_out                       : out  std_logic;
    gt27_txoutclkfabric_out                 : out  std_logic;
    gt27_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt27_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt27_txcharisk_in                       : in   std_logic_vector(7 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT28  (X1Y32)
    --____________________________CHANNEL PORTS________________________________
    GT28_DRP_BUSY_OUT                        : out  std_logic;
    GT28_RXPMARESETDONE_OUT                        : out  std_logic;
    GT28_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt28_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt28_drpclk_in                          : in   std_logic;
    gt28_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt28_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt28_drpen_in                           : in   std_logic;
    gt28_drprdy_out                         : out  std_logic;
    gt28_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt28_eyescanreset_in                    : in   std_logic;
    gt28_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt28_eyescandataerror_out               : out  std_logic;
    gt28_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt28_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt28_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt28_rxusrclk_in                        : in   std_logic;
    gt28_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt28_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt28_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt28_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt28_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt28_rxdlyen_in                         : in   std_logic;
    gt28_rxdlysreset_in                     : in   std_logic;
    gt28_rxdlysresetdone_out                : out  std_logic;
    gt28_rxphalign_in                       : in   std_logic;
    gt28_rxphaligndone_out                  : out  std_logic;
    gt28_rxphalignen_in                     : in   std_logic;
    gt28_rxphdlyreset_in                    : in   std_logic;
    gt28_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt28_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt28_rxsyncallin_in                     : in   std_logic;
    gt28_rxsyncdone_out                     : out  std_logic;
    gt28_rxsyncin_in                        : in   std_logic;
    gt28_rxsyncmode_in                      : in   std_logic;
    gt28_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt28_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt28_rxlpmhfhold_in                     : in   std_logic;
    gt28_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt28_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt28_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt28_rxoutclk_out                       : out  std_logic;
    gt28_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt28_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt28_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt28_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt28_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt28_gttxreset_in                       : in   std_logic;
    gt28_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt28_txusrclk_in                        : in   std_logic;
    gt28_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt28_txdlyen_in                         : in   std_logic;
    gt28_txdlysreset_in                     : in   std_logic;
    gt28_txdlysresetdone_out                : out  std_logic;
    gt28_txphalign_in                       : in   std_logic;
    gt28_txphaligndone_out                  : out  std_logic;
    gt28_txphalignen_in                     : in   std_logic;
    gt28_txphdlyreset_in                    : in   std_logic;
    gt28_txphinit_in                        : in   std_logic;
    gt28_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt28_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt28_gthtxn_out                         : out  std_logic;
    gt28_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt28_txoutclk_out                       : out  std_logic;
    gt28_txoutclkfabric_out                 : out  std_logic;
    gt28_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt28_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt28_txcharisk_in                       : in   std_logic_vector(7 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT29  (X1Y33)
    --____________________________CHANNEL PORTS________________________________
    GT29_DRP_BUSY_OUT                        : out  std_logic;
    GT29_RXPMARESETDONE_OUT                        : out  std_logic;
    GT29_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt29_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt29_drpclk_in                          : in   std_logic;
    gt29_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt29_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt29_drpen_in                           : in   std_logic;
    gt29_drprdy_out                         : out  std_logic;
    gt29_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt29_eyescanreset_in                    : in   std_logic;
    gt29_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt29_eyescandataerror_out               : out  std_logic;
    gt29_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt29_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt29_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt29_rxusrclk_in                        : in   std_logic;
    gt29_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt29_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt29_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt29_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt29_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt29_rxdlyen_in                         : in   std_logic;
    gt29_rxdlysreset_in                     : in   std_logic;
    gt29_rxdlysresetdone_out                : out  std_logic;
    gt29_rxphalign_in                       : in   std_logic;
    gt29_rxphaligndone_out                  : out  std_logic;
    gt29_rxphalignen_in                     : in   std_logic;
    gt29_rxphdlyreset_in                    : in   std_logic;
    gt29_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt29_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt29_rxsyncallin_in                     : in   std_logic;
    gt29_rxsyncdone_out                     : out  std_logic;
    gt29_rxsyncin_in                        : in   std_logic;
    gt29_rxsyncmode_in                      : in   std_logic;
    gt29_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt29_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt29_rxlpmhfhold_in                     : in   std_logic;
    gt29_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt29_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt29_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt29_rxoutclk_out                       : out  std_logic;
    gt29_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt29_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt29_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt29_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt29_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt29_gttxreset_in                       : in   std_logic;
    gt29_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt29_txusrclk_in                        : in   std_logic;
    gt29_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt29_txdlyen_in                         : in   std_logic;
    gt29_txdlysreset_in                     : in   std_logic;
    gt29_txdlysresetdone_out                : out  std_logic;
    gt29_txphalign_in                       : in   std_logic;
    gt29_txphaligndone_out                  : out  std_logic;
    gt29_txphalignen_in                     : in   std_logic;
    gt29_txphdlyreset_in                    : in   std_logic;
    gt29_txphinit_in                        : in   std_logic;
    gt29_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt29_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt29_gthtxn_out                         : out  std_logic;
    gt29_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt29_txoutclk_out                       : out  std_logic;
    gt29_txoutclkfabric_out                 : out  std_logic;
    gt29_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt29_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt29_txcharisk_in                       : in   std_logic_vector(7 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT30  (X1Y34)
    --____________________________CHANNEL PORTS________________________________
    GT30_DRP_BUSY_OUT                        : out  std_logic;
    GT30_RXPMARESETDONE_OUT                        : out  std_logic;
    GT30_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt30_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt30_drpclk_in                          : in   std_logic;
    gt30_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt30_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt30_drpen_in                           : in   std_logic;
    gt30_drprdy_out                         : out  std_logic;
    gt30_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt30_eyescanreset_in                    : in   std_logic;
    gt30_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt30_eyescandataerror_out               : out  std_logic;
    gt30_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt30_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt30_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt30_rxusrclk_in                        : in   std_logic;
    gt30_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt30_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt30_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt30_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt30_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt30_rxdlyen_in                         : in   std_logic;
    gt30_rxdlysreset_in                     : in   std_logic;
    gt30_rxdlysresetdone_out                : out  std_logic;
    gt30_rxphalign_in                       : in   std_logic;
    gt30_rxphaligndone_out                  : out  std_logic;
    gt30_rxphalignen_in                     : in   std_logic;
    gt30_rxphdlyreset_in                    : in   std_logic;
    gt30_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt30_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt30_rxsyncallin_in                     : in   std_logic;
    gt30_rxsyncdone_out                     : out  std_logic;
    gt30_rxsyncin_in                        : in   std_logic;
    gt30_rxsyncmode_in                      : in   std_logic;
    gt30_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt30_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt30_rxlpmhfhold_in                     : in   std_logic;
    gt30_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt30_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt30_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt30_rxoutclk_out                       : out  std_logic;
    gt30_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt30_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt30_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt30_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt30_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt30_gttxreset_in                       : in   std_logic;
    gt30_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt30_txusrclk_in                        : in   std_logic;
    gt30_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt30_txdlyen_in                         : in   std_logic;
    gt30_txdlysreset_in                     : in   std_logic;
    gt30_txdlysresetdone_out                : out  std_logic;
    gt30_txphalign_in                       : in   std_logic;
    gt30_txphaligndone_out                  : out  std_logic;
    gt30_txphalignen_in                     : in   std_logic;
    gt30_txphdlyreset_in                    : in   std_logic;
    gt30_txphinit_in                        : in   std_logic;
    gt30_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt30_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt30_gthtxn_out                         : out  std_logic;
    gt30_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt30_txoutclk_out                       : out  std_logic;
    gt30_txoutclkfabric_out                 : out  std_logic;
    gt30_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt30_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt30_txcharisk_in                       : in   std_logic_vector(7 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT31  (X1Y35)
    --____________________________CHANNEL PORTS________________________________
    GT31_DRP_BUSY_OUT                        : out  std_logic;
    GT31_RXPMARESETDONE_OUT                        : out  std_logic;
    GT31_TXPMARESETDONE_OUT                        : out  std_logic;

    ---------------------------- Channel - DRP Ports  --------------------------
    gt31_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt31_drpclk_in                          : in   std_logic;
    gt31_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt31_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt31_drpen_in                           : in   std_logic;
    gt31_drprdy_out                         : out  std_logic;
    gt31_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt31_eyescanreset_in                    : in   std_logic;
    gt31_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt31_eyescandataerror_out               : out  std_logic;
    gt31_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt31_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt31_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt31_rxusrclk_in                        : in   std_logic;
    gt31_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt31_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt31_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt31_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt31_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt31_rxdlyen_in                         : in   std_logic;
    gt31_rxdlysreset_in                     : in   std_logic;
    gt31_rxdlysresetdone_out                : out  std_logic;
    gt31_rxphalign_in                       : in   std_logic;
    gt31_rxphaligndone_out                  : out  std_logic;
    gt31_rxphalignen_in                     : in   std_logic;
    gt31_rxphdlyreset_in                    : in   std_logic;
    gt31_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt31_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt31_rxsyncallin_in                     : in   std_logic;
    gt31_rxsyncdone_out                     : out  std_logic;
    gt31_rxsyncin_in                        : in   std_logic;
    gt31_rxsyncmode_in                      : in   std_logic;
    gt31_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt31_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt31_rxlpmhfhold_in                     : in   std_logic;
    gt31_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt31_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt31_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt31_rxoutclk_out                       : out  std_logic;
    gt31_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt31_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt31_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt31_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt31_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt31_gttxreset_in                       : in   std_logic;
    gt31_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt31_txusrclk_in                        : in   std_logic;
    gt31_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt31_txdlyen_in                         : in   std_logic;
    gt31_txdlysreset_in                     : in   std_logic;
    gt31_txdlysresetdone_out                : out  std_logic;
    gt31_txphalign_in                       : in   std_logic;
    gt31_txphaligndone_out                  : out  std_logic;
    gt31_txphalignen_in                     : in   std_logic;
    gt31_txphdlyreset_in                    : in   std_logic;
    gt31_txphinit_in                        : in   std_logic;
    gt31_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt31_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt31_gthtxn_out                         : out  std_logic;
    gt31_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt31_txoutclk_out                       : out  std_logic;
    gt31_txoutclkfabric_out                 : out  std_logic;
    gt31_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt31_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt31_txcharisk_in                       : in   std_logic_vector(7 downto 0);
   

    --____________________________COMMON PORTS________________________________
     GT0_QPLLOUTCLK_IN   : in std_logic;
     GT0_QPLLRESET_IN  : in std_logic;
     GT0_QPLLOUTREFCLK_IN   : in std_logic;
    --____________________________COMMON PORTS________________________________
     GT1_QPLLOUTCLK_IN   : in std_logic;
     GT1_QPLLRESET_IN  : in std_logic;
     GT1_QPLLOUTREFCLK_IN   : in std_logic;
    --____________________________COMMON PORTS________________________________
     GT2_QPLLOUTCLK_IN   : in std_logic;
     GT2_QPLLRESET_IN  : in std_logic;
     GT2_QPLLOUTREFCLK_IN   : in std_logic;
    --____________________________COMMON PORTS________________________________
     GT3_QPLLOUTCLK_IN   : in std_logic;
     GT3_QPLLRESET_IN  : in std_logic;
     GT3_QPLLOUTREFCLK_IN   : in std_logic;
    --____________________________COMMON PORTS________________________________
     GT4_QPLLOUTCLK_IN   : in std_logic;
     GT4_QPLLRESET_IN  : in std_logic;
     GT4_QPLLOUTREFCLK_IN   : in std_logic;
    --____________________________COMMON PORTS________________________________
     GT5_QPLLOUTCLK_IN   : in std_logic;
     GT5_QPLLRESET_IN  : in std_logic;
     GT5_QPLLOUTREFCLK_IN   : in std_logic;
    --____________________________COMMON PORTS________________________________
     GT6_QPLLOUTCLK_IN   : in std_logic;
     GT6_QPLLRESET_IN  : in std_logic;
     GT6_QPLLOUTREFCLK_IN   : in std_logic;
    --____________________________COMMON PORTS________________________________
     GT7_QPLLOUTCLK_IN   : in std_logic;
     GT7_QPLLRESET_IN  : in std_logic;
     GT7_QPLLOUTREFCLK_IN   : in std_logic

);
end component;

component gtwizard_0_TX_STARTUP_FSM
  Generic(
           EXAMPLE_SIMULATION       : integer := 0;
           STABLE_CLOCK_PERIOD      : integer range 4 to 250 := 8; --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   : integer range 2 to 8  := 8; 
           TX_QPLL_USED             : boolean := False;           -- the TX and RX Reset FSMs must
           RX_QPLL_USED             : boolean := False;           -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   : boolean := True             -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                  -- is enough. For single-lane applications the automatic alignment is 
                                                                  -- sufficient              
         );     
    Port ( STABLE_CLOCK             : in  STD_LOGIC;              --Stable Clock, either a stable clock from the PCB
                                                                  --or reference-clock present at startup.
           TXUSERCLK                : in  STD_LOGIC;              --TXUSERCLK as used in the design
           SOFT_RESET               : in  STD_LOGIC;              --User Reset, can be pulled any time
           QPLLREFCLKLOST           : in  STD_LOGIC;              --QPLL Reference-clock for the GT is lost
           CPLLREFCLKLOST           : in  STD_LOGIC;              --CPLL Reference-clock for the GT is lost
           QPLLLOCK                 : in  STD_LOGIC;              --Lock Detect from the QPLL of the GT
           CPLLLOCK                 : in  STD_LOGIC;              --Lock Detect from the CPLL of the GT
           TXRESETDONE              : in  STD_LOGIC;      
           MMCM_LOCK                : in  STD_LOGIC;      
           GTTXRESET                : out STD_LOGIC:='0';      
           MMCM_RESET               : out STD_LOGIC:='0';      
           QPLL_RESET               : out STD_LOGIC:='0';        --Reset QPLL
           CPLL_RESET               : out STD_LOGIC:='0';        --Reset CPLL
           TX_FSM_RESET_DONE        : out STD_LOGIC:='0';        --Reset-sequence has sucessfully been finished.
           TXUSERRDY                : out STD_LOGIC:='0';
           RUN_PHALIGNMENT          : out STD_LOGIC:='0';
           RESET_PHALIGNMENT        : out STD_LOGIC:='0';
           PHALIGNMENT_DONE         : in  STD_LOGIC;
           
           RETRY_COUNTER            : out  STD_LOGIC_VECTOR (RETRY_COUNTER_BITWIDTH-1 downto 0):=(others=>'0')-- Number of 
                                                            -- Retries it took to get the transceiver up and running
           );
end component;

component gtwizard_0_RX_STARTUP_FSM
  Generic(
           EXAMPLE_SIMULATION       : integer := 0;
           EQ_MODE                  : string := "DFE";
           STABLE_CLOCK_PERIOD      : integer range 4 to 250 := 8; --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   : integer range 2 to 8  := 8; 
           TX_QPLL_USED             : boolean := False;           -- the TX and RX Reset FSMs must
           RX_QPLL_USED             : boolean := False;           -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   : boolean := True             -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                  -- is enough. For single-lane applications the automatic alignment is 
                                                                  -- sufficient                         
         );     
    Port ( STABLE_CLOCK             : in  STD_LOGIC;        --Stable Clock, either a stable clock from the PCB
                                                            --or reference-clock present at startup.
           RXUSERCLK                : in  STD_LOGIC;        --RXUSERCLK as used in the design
           SOFT_RESET               : in  STD_LOGIC;        --User Reset, can be pulled any time
           RXPMARESETDONE               : in  STD_LOGIC;              
           RXOUTCLK               : in  STD_LOGIC; 
             
           QPLLREFCLKLOST           : in  STD_LOGIC;        --QPLL Reference-clock for the GT is lost
           CPLLREFCLKLOST           : in  STD_LOGIC;        --CPLL Reference-clock for the GT is lost
           QPLLLOCK                 : in  STD_LOGIC;        --Lock Detect from the QPLL of the GT
           CPLLLOCK                 : in  STD_LOGIC;        --Lock Detect from the CPLL of the GT
           RXRESETDONE              : in  STD_LOGIC;
           MMCM_LOCK                : in  STD_LOGIC;
           RECCLK_STABLE            : in  STD_LOGIC;
           RECCLK_MONITOR_RESTART   : in  STD_LOGIC;
           DATA_VALID               : in  STD_LOGIC;
           TXUSERRDY                : in  STD_LOGIC;       --TXUSERRDY from GT 
           DONT_RESET_ON_DATA_ERROR : in  STD_LOGIC;
           GTRXRESET                : out STD_LOGIC:='0';
           MMCM_RESET               : out STD_LOGIC:='0';
           QPLL_RESET               : out STD_LOGIC:='0';  --Reset QPLL (only if RX uses QPLL)
           CPLL_RESET               : out STD_LOGIC:='0';  --Reset CPLL (only if RX uses CPLL)
           RX_FSM_RESET_DONE        : out STD_LOGIC:='0';  --Reset-sequence has sucessfully been finished.
           RXUSERRDY                : out STD_LOGIC:='0';
           RUN_PHALIGNMENT          : out STD_LOGIC;
           PHALIGNMENT_DONE         : in  STD_LOGIC; 
           RESET_PHALIGNMENT        : out STD_LOGIC:='0';           
           RXDFEAGCHOLD             : out STD_LOGIC;
           RXDFELFHOLD              : out STD_LOGIC;
           RXLPMLFHOLD              : out STD_LOGIC;
           RXLPMHFHOLD              : out STD_LOGIC;
           RETRY_COUNTER            : out STD_LOGIC_VECTOR (RETRY_COUNTER_BITWIDTH-1 downto 0):=(others=>'0')-- Number of 
                                                            -- Retries it took to get the transceiver up and running
           );
end component;




component gtwizard_0_AUTO_PHASE_ALIGN     
    port ( STABLE_CLOCK             : in  STD_LOGIC;              --Stable Clock, either a stable clock from the PCB
                                                                  --or reference-clock present at startup.
           RUN_PHALIGNMENT          : in  STD_LOGIC;              --Signal from the main Reset-FSM to run the auto phase-alignment procedure
           PHASE_ALIGNMENT_DONE     : out STD_LOGIC;              -- Auto phase-alignment performed sucessfully
           PHALIGNDONE              : in  STD_LOGIC;              --\ Phase-alignment signals from and to the
           DLYSRESET                : out STD_LOGIC;              -- |transceiver.
           DLYSRESETDONE            : in  STD_LOGIC;              --/
           RECCLKSTABLE             : in  STD_LOGIC               --/on the RX-side.
           
           );
end component;


component gtwizard_0_TX_MANUAL_PHASE_ALIGN 
  Generic( NUMBER_OF_LANES          : integer range 1 to 32:= 4;  -- Number of lanes that are controlled using this FSM.
           MASTER_LANE_ID           : integer range 0 to 31:= 0   -- Number of the lane which is considered the master in manual phase-alignment
         );     

    Port ( STABLE_CLOCK             : in  STD_LOGIC;              --Stable Clock, either a stable clock from the PCB
                                                                  --or reference-clock present at startup.
           RESET_PHALIGNMENT        : in  STD_LOGIC;
           RUN_PHALIGNMENT          : in  STD_LOGIC;
           PHASE_ALIGNMENT_DONE     : out STD_LOGIC := '0';       -- Manual phase-alignment performed sucessfully  
           TXDLYSRESET              : out STD_LOGIC_VECTOR(NUMBER_OF_LANES-1 downto 0) := (others=> '0');
           TXDLYSRESETDONE          : in  STD_LOGIC_VECTOR(NUMBER_OF_LANES-1 downto 0);
           TXPHINIT                 : out STD_LOGIC_VECTOR(NUMBER_OF_LANES-1 downto 0) := (others=> '0');
           TXPHINITDONE             : in  STD_LOGIC_VECTOR(NUMBER_OF_LANES-1 downto 0);
           TXPHALIGN                : out STD_LOGIC_VECTOR(NUMBER_OF_LANES-1 downto 0) := (others=> '0');
           TXPHALIGNDONE            : in  STD_LOGIC_VECTOR(NUMBER_OF_LANES-1 downto 0);
           TXDLYEN                  : out STD_LOGIC_VECTOR(NUMBER_OF_LANES-1 downto 0) := (others=> '0')
           );
end component;

component gtwizard_0_RX_MANUAL_PHASE_ALIGN 
  Generic( NUMBER_OF_LANES          : integer range 1 to 32:= 4;  -- Number of lanes that are controlled using this FSM.
           MASTER_LANE_ID           : integer range 0 to 31:= 0   -- Number of the lane which is considered the master in manual phase-alignment
         );     

    Port ( STABLE_CLOCK             : in  STD_LOGIC;              --Stable Clock, either a stable clock from the PCB
                                                                  --or reference-clock present at startup.
           RESET_PHALIGNMENT        : in  STD_LOGIC;
           RUN_PHALIGNMENT          : in  STD_LOGIC;
           PHASE_ALIGNMENT_DONE     : out STD_LOGIC := '0';       -- Manual phase-alignment performed sucessfully    
           RXDLYSRESET              : out STD_LOGIC_VECTOR(NUMBER_OF_LANES-1 downto 0) := (others=> '0');
           RXDLYSRESETDONE          : in  STD_LOGIC_VECTOR(NUMBER_OF_LANES-1 downto 0);
           RXPHALIGN                : out STD_LOGIC_VECTOR(NUMBER_OF_LANES-1 downto 0) := (others=> '0');
           RXPHALIGNDONE            : in  STD_LOGIC_VECTOR(NUMBER_OF_LANES-1 downto 0);
           RXDLYEN                  : out STD_LOGIC_VECTOR(NUMBER_OF_LANES-1 downto 0) := (others=> '0')
           );
end component;

  function get_cdrlock_time(is_sim : in integer) return integer is
    variable lock_time: integer;
  begin
    if (is_sim = 1) then
      lock_time := 1000;
    else
      lock_time := 100000 / integer(5); --Typical CDR lock time is 50,000UI as per DS183
    end if;
    return lock_time;
  end function;


--***********************************Parameter Declarations********************

    constant DLY : time := 1 ns;
    constant RX_CDRLOCK_TIME      : integer := get_cdrlock_time(EXAMPLE_SIMULATION);       -- 200us
    constant WAIT_TIME_CDRLOCK    : integer := RX_CDRLOCK_TIME / STABLE_CLOCK_PERIOD;      -- 200 us time-out



    -------------------------- GT Wrapper Wires ------------------------------
    signal   gt0_txpmaresetdone_i            : std_logic;
    signal   gt0_rxpmaresetdone_i            : std_logic;
    signal   gt0_txresetdone_i               : std_logic;
    signal   gt0_rxresetdone_i               : std_logic;
    signal   gt0_txresetdone_ii              : std_logic;
    signal   gt0_rxresetdone_ii              : std_logic;
    signal   gt0_gttxreset_i                 : std_logic;
    signal   gt0_gttxreset_t                 : std_logic;
    signal   gt0_gtrxreset_i                 : std_logic;
    signal   gt0_gtrxreset_t                 : std_logic;
    signal   gt0_txuserrdy_i                 : std_logic;
    signal   gt0_txuserrdy_t                 : std_logic;
    signal   gt0_rxuserrdy_i                 : std_logic;
    signal   gt0_rxuserrdy_t                 : std_logic;

    signal   gt0_rxdfeagchold_i              : std_logic;
    signal   gt0_rxdfelfhold_i               : std_logic;
    signal   gt0_rxlpmlfhold_i               : std_logic;
    signal   gt0_rxlpmhfhold_i               : std_logic;


    signal   gt1_txpmaresetdone_i            : std_logic;
    signal   gt1_rxpmaresetdone_i            : std_logic;
    signal   gt1_txresetdone_i               : std_logic;
    signal   gt1_rxresetdone_i               : std_logic;
    signal   gt1_txresetdone_ii              : std_logic;
    signal   gt1_rxresetdone_ii              : std_logic;
    signal   gt1_gttxreset_i                 : std_logic;
    signal   gt1_gttxreset_t                 : std_logic;
    signal   gt1_gtrxreset_i                 : std_logic;
    signal   gt1_gtrxreset_t                 : std_logic;
    signal   gt1_txuserrdy_i                 : std_logic;
    signal   gt1_txuserrdy_t                 : std_logic;
    signal   gt1_rxuserrdy_i                 : std_logic;
    signal   gt1_rxuserrdy_t                 : std_logic;

    signal   gt1_rxdfeagchold_i              : std_logic;
    signal   gt1_rxdfelfhold_i               : std_logic;
    signal   gt1_rxlpmlfhold_i               : std_logic;
    signal   gt1_rxlpmhfhold_i               : std_logic;


    signal   gt2_txpmaresetdone_i            : std_logic;
    signal   gt2_rxpmaresetdone_i            : std_logic;
    signal   gt2_txresetdone_i               : std_logic;
    signal   gt2_rxresetdone_i               : std_logic;
    signal   gt2_txresetdone_ii              : std_logic;
    signal   gt2_rxresetdone_ii              : std_logic;
    signal   gt2_gttxreset_i                 : std_logic;
    signal   gt2_gttxreset_t                 : std_logic;
    signal   gt2_gtrxreset_i                 : std_logic;
    signal   gt2_gtrxreset_t                 : std_logic;
    signal   gt2_txuserrdy_i                 : std_logic;
    signal   gt2_txuserrdy_t                 : std_logic;
    signal   gt2_rxuserrdy_i                 : std_logic;
    signal   gt2_rxuserrdy_t                 : std_logic;

    signal   gt2_rxdfeagchold_i              : std_logic;
    signal   gt2_rxdfelfhold_i               : std_logic;
    signal   gt2_rxlpmlfhold_i               : std_logic;
    signal   gt2_rxlpmhfhold_i               : std_logic;


    signal   gt3_txpmaresetdone_i            : std_logic;
    signal   gt3_rxpmaresetdone_i            : std_logic;
    signal   gt3_txresetdone_i               : std_logic;
    signal   gt3_rxresetdone_i               : std_logic;
    signal   gt3_txresetdone_ii              : std_logic;
    signal   gt3_rxresetdone_ii              : std_logic;
    signal   gt3_gttxreset_i                 : std_logic;
    signal   gt3_gttxreset_t                 : std_logic;
    signal   gt3_gtrxreset_i                 : std_logic;
    signal   gt3_gtrxreset_t                 : std_logic;
    signal   gt3_txuserrdy_i                 : std_logic;
    signal   gt3_txuserrdy_t                 : std_logic;
    signal   gt3_rxuserrdy_i                 : std_logic;
    signal   gt3_rxuserrdy_t                 : std_logic;

    signal   gt3_rxdfeagchold_i              : std_logic;
    signal   gt3_rxdfelfhold_i               : std_logic;
    signal   gt3_rxlpmlfhold_i               : std_logic;
    signal   gt3_rxlpmhfhold_i               : std_logic;


    signal   gt4_txpmaresetdone_i            : std_logic;
    signal   gt4_rxpmaresetdone_i            : std_logic;
    signal   gt4_txresetdone_i               : std_logic;
    signal   gt4_rxresetdone_i               : std_logic;
    signal   gt4_txresetdone_ii              : std_logic;
    signal   gt4_rxresetdone_ii              : std_logic;
    signal   gt4_gttxreset_i                 : std_logic;
    signal   gt4_gttxreset_t                 : std_logic;
    signal   gt4_gtrxreset_i                 : std_logic;
    signal   gt4_gtrxreset_t                 : std_logic;
    signal   gt4_txuserrdy_i                 : std_logic;
    signal   gt4_txuserrdy_t                 : std_logic;
    signal   gt4_rxuserrdy_i                 : std_logic;
    signal   gt4_rxuserrdy_t                 : std_logic;

    signal   gt4_rxdfeagchold_i              : std_logic;
    signal   gt4_rxdfelfhold_i               : std_logic;
    signal   gt4_rxlpmlfhold_i               : std_logic;
    signal   gt4_rxlpmhfhold_i               : std_logic;


    signal   gt5_txpmaresetdone_i            : std_logic;
    signal   gt5_rxpmaresetdone_i            : std_logic;
    signal   gt5_txresetdone_i               : std_logic;
    signal   gt5_rxresetdone_i               : std_logic;
    signal   gt5_txresetdone_ii              : std_logic;
    signal   gt5_rxresetdone_ii              : std_logic;
    signal   gt5_gttxreset_i                 : std_logic;
    signal   gt5_gttxreset_t                 : std_logic;
    signal   gt5_gtrxreset_i                 : std_logic;
    signal   gt5_gtrxreset_t                 : std_logic;
    signal   gt5_txuserrdy_i                 : std_logic;
    signal   gt5_txuserrdy_t                 : std_logic;
    signal   gt5_rxuserrdy_i                 : std_logic;
    signal   gt5_rxuserrdy_t                 : std_logic;

    signal   gt5_rxdfeagchold_i              : std_logic;
    signal   gt5_rxdfelfhold_i               : std_logic;
    signal   gt5_rxlpmlfhold_i               : std_logic;
    signal   gt5_rxlpmhfhold_i               : std_logic;


    signal   gt6_txpmaresetdone_i            : std_logic;
    signal   gt6_rxpmaresetdone_i            : std_logic;
    signal   gt6_txresetdone_i               : std_logic;
    signal   gt6_rxresetdone_i               : std_logic;
    signal   gt6_txresetdone_ii              : std_logic;
    signal   gt6_rxresetdone_ii              : std_logic;
    signal   gt6_gttxreset_i                 : std_logic;
    signal   gt6_gttxreset_t                 : std_logic;
    signal   gt6_gtrxreset_i                 : std_logic;
    signal   gt6_gtrxreset_t                 : std_logic;
    signal   gt6_txuserrdy_i                 : std_logic;
    signal   gt6_txuserrdy_t                 : std_logic;
    signal   gt6_rxuserrdy_i                 : std_logic;
    signal   gt6_rxuserrdy_t                 : std_logic;

    signal   gt6_rxdfeagchold_i              : std_logic;
    signal   gt6_rxdfelfhold_i               : std_logic;
    signal   gt6_rxlpmlfhold_i               : std_logic;
    signal   gt6_rxlpmhfhold_i               : std_logic;


    signal   gt7_txpmaresetdone_i            : std_logic;
    signal   gt7_rxpmaresetdone_i            : std_logic;
    signal   gt7_txresetdone_i               : std_logic;
    signal   gt7_rxresetdone_i               : std_logic;
    signal   gt7_txresetdone_ii              : std_logic;
    signal   gt7_rxresetdone_ii              : std_logic;
    signal   gt7_gttxreset_i                 : std_logic;
    signal   gt7_gttxreset_t                 : std_logic;
    signal   gt7_gtrxreset_i                 : std_logic;
    signal   gt7_gtrxreset_t                 : std_logic;
    signal   gt7_txuserrdy_i                 : std_logic;
    signal   gt7_txuserrdy_t                 : std_logic;
    signal   gt7_rxuserrdy_i                 : std_logic;
    signal   gt7_rxuserrdy_t                 : std_logic;

    signal   gt7_rxdfeagchold_i              : std_logic;
    signal   gt7_rxdfelfhold_i               : std_logic;
    signal   gt7_rxlpmlfhold_i               : std_logic;
    signal   gt7_rxlpmhfhold_i               : std_logic;


    signal   gt8_txpmaresetdone_i            : std_logic;
    signal   gt8_rxpmaresetdone_i            : std_logic;
    signal   gt8_txresetdone_i               : std_logic;
    signal   gt8_rxresetdone_i               : std_logic;
    signal   gt8_txresetdone_ii              : std_logic;
    signal   gt8_rxresetdone_ii              : std_logic;
    signal   gt8_gttxreset_i                 : std_logic;
    signal   gt8_gttxreset_t                 : std_logic;
    signal   gt8_gtrxreset_i                 : std_logic;
    signal   gt8_gtrxreset_t                 : std_logic;
    signal   gt8_txuserrdy_i                 : std_logic;
    signal   gt8_txuserrdy_t                 : std_logic;
    signal   gt8_rxuserrdy_i                 : std_logic;
    signal   gt8_rxuserrdy_t                 : std_logic;

    signal   gt8_rxdfeagchold_i              : std_logic;
    signal   gt8_rxdfelfhold_i               : std_logic;
    signal   gt8_rxlpmlfhold_i               : std_logic;
    signal   gt8_rxlpmhfhold_i               : std_logic;


    signal   gt9_txpmaresetdone_i            : std_logic;
    signal   gt9_rxpmaresetdone_i            : std_logic;
    signal   gt9_txresetdone_i               : std_logic;
    signal   gt9_rxresetdone_i               : std_logic;
    signal   gt9_txresetdone_ii              : std_logic;
    signal   gt9_rxresetdone_ii              : std_logic;
    signal   gt9_gttxreset_i                 : std_logic;
    signal   gt9_gttxreset_t                 : std_logic;
    signal   gt9_gtrxreset_i                 : std_logic;
    signal   gt9_gtrxreset_t                 : std_logic;
    signal   gt9_txuserrdy_i                 : std_logic;
    signal   gt9_txuserrdy_t                 : std_logic;
    signal   gt9_rxuserrdy_i                 : std_logic;
    signal   gt9_rxuserrdy_t                 : std_logic;

    signal   gt9_rxdfeagchold_i              : std_logic;
    signal   gt9_rxdfelfhold_i               : std_logic;
    signal   gt9_rxlpmlfhold_i               : std_logic;
    signal   gt9_rxlpmhfhold_i               : std_logic;


    signal   gt10_txpmaresetdone_i           : std_logic;
    signal   gt10_rxpmaresetdone_i           : std_logic;
    signal   gt10_txresetdone_i              : std_logic;
    signal   gt10_rxresetdone_i              : std_logic;
    signal   gt10_txresetdone_ii             : std_logic;
    signal   gt10_rxresetdone_ii             : std_logic;
    signal   gt10_gttxreset_i                : std_logic;
    signal   gt10_gttxreset_t                : std_logic;
    signal   gt10_gtrxreset_i                : std_logic;
    signal   gt10_gtrxreset_t                : std_logic;
    signal   gt10_txuserrdy_i                : std_logic;
    signal   gt10_txuserrdy_t                : std_logic;
    signal   gt10_rxuserrdy_i                : std_logic;
    signal   gt10_rxuserrdy_t                : std_logic;

    signal   gt10_rxdfeagchold_i             : std_logic;
    signal   gt10_rxdfelfhold_i              : std_logic;
    signal   gt10_rxlpmlfhold_i              : std_logic;
    signal   gt10_rxlpmhfhold_i              : std_logic;


    signal   gt11_txpmaresetdone_i           : std_logic;
    signal   gt11_rxpmaresetdone_i           : std_logic;
    signal   gt11_txresetdone_i              : std_logic;
    signal   gt11_rxresetdone_i              : std_logic;
    signal   gt11_txresetdone_ii             : std_logic;
    signal   gt11_rxresetdone_ii             : std_logic;
    signal   gt11_gttxreset_i                : std_logic;
    signal   gt11_gttxreset_t                : std_logic;
    signal   gt11_gtrxreset_i                : std_logic;
    signal   gt11_gtrxreset_t                : std_logic;
    signal   gt11_txuserrdy_i                : std_logic;
    signal   gt11_txuserrdy_t                : std_logic;
    signal   gt11_rxuserrdy_i                : std_logic;
    signal   gt11_rxuserrdy_t                : std_logic;

    signal   gt11_rxdfeagchold_i             : std_logic;
    signal   gt11_rxdfelfhold_i              : std_logic;
    signal   gt11_rxlpmlfhold_i              : std_logic;
    signal   gt11_rxlpmhfhold_i              : std_logic;


    signal   gt12_txpmaresetdone_i           : std_logic;
    signal   gt12_rxpmaresetdone_i           : std_logic;
    signal   gt12_txresetdone_i              : std_logic;
    signal   gt12_rxresetdone_i              : std_logic;
    signal   gt12_txresetdone_ii             : std_logic;
    signal   gt12_rxresetdone_ii             : std_logic;
    signal   gt12_gttxreset_i                : std_logic;
    signal   gt12_gttxreset_t                : std_logic;
    signal   gt12_gtrxreset_i                : std_logic;
    signal   gt12_gtrxreset_t                : std_logic;
    signal   gt12_txuserrdy_i                : std_logic;
    signal   gt12_txuserrdy_t                : std_logic;
    signal   gt12_rxuserrdy_i                : std_logic;
    signal   gt12_rxuserrdy_t                : std_logic;

    signal   gt12_rxdfeagchold_i             : std_logic;
    signal   gt12_rxdfelfhold_i              : std_logic;
    signal   gt12_rxlpmlfhold_i              : std_logic;
    signal   gt12_rxlpmhfhold_i              : std_logic;


    signal   gt13_txpmaresetdone_i           : std_logic;
    signal   gt13_rxpmaresetdone_i           : std_logic;
    signal   gt13_txresetdone_i              : std_logic;
    signal   gt13_rxresetdone_i              : std_logic;
    signal   gt13_txresetdone_ii             : std_logic;
    signal   gt13_rxresetdone_ii             : std_logic;
    signal   gt13_gttxreset_i                : std_logic;
    signal   gt13_gttxreset_t                : std_logic;
    signal   gt13_gtrxreset_i                : std_logic;
    signal   gt13_gtrxreset_t                : std_logic;
    signal   gt13_txuserrdy_i                : std_logic;
    signal   gt13_txuserrdy_t                : std_logic;
    signal   gt13_rxuserrdy_i                : std_logic;
    signal   gt13_rxuserrdy_t                : std_logic;

    signal   gt13_rxdfeagchold_i             : std_logic;
    signal   gt13_rxdfelfhold_i              : std_logic;
    signal   gt13_rxlpmlfhold_i              : std_logic;
    signal   gt13_rxlpmhfhold_i              : std_logic;


    signal   gt14_txpmaresetdone_i           : std_logic;
    signal   gt14_rxpmaresetdone_i           : std_logic;
    signal   gt14_txresetdone_i              : std_logic;
    signal   gt14_rxresetdone_i              : std_logic;
    signal   gt14_txresetdone_ii             : std_logic;
    signal   gt14_rxresetdone_ii             : std_logic;
    signal   gt14_gttxreset_i                : std_logic;
    signal   gt14_gttxreset_t                : std_logic;
    signal   gt14_gtrxreset_i                : std_logic;
    signal   gt14_gtrxreset_t                : std_logic;
    signal   gt14_txuserrdy_i                : std_logic;
    signal   gt14_txuserrdy_t                : std_logic;
    signal   gt14_rxuserrdy_i                : std_logic;
    signal   gt14_rxuserrdy_t                : std_logic;

    signal   gt14_rxdfeagchold_i             : std_logic;
    signal   gt14_rxdfelfhold_i              : std_logic;
    signal   gt14_rxlpmlfhold_i              : std_logic;
    signal   gt14_rxlpmhfhold_i              : std_logic;


    signal   gt15_txpmaresetdone_i           : std_logic;
    signal   gt15_rxpmaresetdone_i           : std_logic;
    signal   gt15_txresetdone_i              : std_logic;
    signal   gt15_rxresetdone_i              : std_logic;
    signal   gt15_txresetdone_ii             : std_logic;
    signal   gt15_rxresetdone_ii             : std_logic;
    signal   gt15_gttxreset_i                : std_logic;
    signal   gt15_gttxreset_t                : std_logic;
    signal   gt15_gtrxreset_i                : std_logic;
    signal   gt15_gtrxreset_t                : std_logic;
    signal   gt15_txuserrdy_i                : std_logic;
    signal   gt15_txuserrdy_t                : std_logic;
    signal   gt15_rxuserrdy_i                : std_logic;
    signal   gt15_rxuserrdy_t                : std_logic;

    signal   gt15_rxdfeagchold_i             : std_logic;
    signal   gt15_rxdfelfhold_i              : std_logic;
    signal   gt15_rxlpmlfhold_i              : std_logic;
    signal   gt15_rxlpmhfhold_i              : std_logic;


    signal   gt16_txpmaresetdone_i           : std_logic;
    signal   gt16_rxpmaresetdone_i           : std_logic;
    signal   gt16_txresetdone_i              : std_logic;
    signal   gt16_rxresetdone_i              : std_logic;
    signal   gt16_txresetdone_ii             : std_logic;
    signal   gt16_rxresetdone_ii             : std_logic;
    signal   gt16_gttxreset_i                : std_logic;
    signal   gt16_gttxreset_t                : std_logic;
    signal   gt16_gtrxreset_i                : std_logic;
    signal   gt16_gtrxreset_t                : std_logic;
    signal   gt16_txuserrdy_i                : std_logic;
    signal   gt16_txuserrdy_t                : std_logic;
    signal   gt16_rxuserrdy_i                : std_logic;
    signal   gt16_rxuserrdy_t                : std_logic;

    signal   gt16_rxdfeagchold_i             : std_logic;
    signal   gt16_rxdfelfhold_i              : std_logic;
    signal   gt16_rxlpmlfhold_i              : std_logic;
    signal   gt16_rxlpmhfhold_i              : std_logic;


    signal   gt17_txpmaresetdone_i           : std_logic;
    signal   gt17_rxpmaresetdone_i           : std_logic;
    signal   gt17_txresetdone_i              : std_logic;
    signal   gt17_rxresetdone_i              : std_logic;
    signal   gt17_txresetdone_ii             : std_logic;
    signal   gt17_rxresetdone_ii             : std_logic;
    signal   gt17_gttxreset_i                : std_logic;
    signal   gt17_gttxreset_t                : std_logic;
    signal   gt17_gtrxreset_i                : std_logic;
    signal   gt17_gtrxreset_t                : std_logic;
    signal   gt17_txuserrdy_i                : std_logic;
    signal   gt17_txuserrdy_t                : std_logic;
    signal   gt17_rxuserrdy_i                : std_logic;
    signal   gt17_rxuserrdy_t                : std_logic;

    signal   gt17_rxdfeagchold_i             : std_logic;
    signal   gt17_rxdfelfhold_i              : std_logic;
    signal   gt17_rxlpmlfhold_i              : std_logic;
    signal   gt17_rxlpmhfhold_i              : std_logic;


    signal   gt18_txpmaresetdone_i           : std_logic;
    signal   gt18_rxpmaresetdone_i           : std_logic;
    signal   gt18_txresetdone_i              : std_logic;
    signal   gt18_rxresetdone_i              : std_logic;
    signal   gt18_txresetdone_ii             : std_logic;
    signal   gt18_rxresetdone_ii             : std_logic;
    signal   gt18_gttxreset_i                : std_logic;
    signal   gt18_gttxreset_t                : std_logic;
    signal   gt18_gtrxreset_i                : std_logic;
    signal   gt18_gtrxreset_t                : std_logic;
    signal   gt18_txuserrdy_i                : std_logic;
    signal   gt18_txuserrdy_t                : std_logic;
    signal   gt18_rxuserrdy_i                : std_logic;
    signal   gt18_rxuserrdy_t                : std_logic;

    signal   gt18_rxdfeagchold_i             : std_logic;
    signal   gt18_rxdfelfhold_i              : std_logic;
    signal   gt18_rxlpmlfhold_i              : std_logic;
    signal   gt18_rxlpmhfhold_i              : std_logic;


    signal   gt19_txpmaresetdone_i           : std_logic;
    signal   gt19_rxpmaresetdone_i           : std_logic;
    signal   gt19_txresetdone_i              : std_logic;
    signal   gt19_rxresetdone_i              : std_logic;
    signal   gt19_txresetdone_ii             : std_logic;
    signal   gt19_rxresetdone_ii             : std_logic;
    signal   gt19_gttxreset_i                : std_logic;
    signal   gt19_gttxreset_t                : std_logic;
    signal   gt19_gtrxreset_i                : std_logic;
    signal   gt19_gtrxreset_t                : std_logic;
    signal   gt19_txuserrdy_i                : std_logic;
    signal   gt19_txuserrdy_t                : std_logic;
    signal   gt19_rxuserrdy_i                : std_logic;
    signal   gt19_rxuserrdy_t                : std_logic;

    signal   gt19_rxdfeagchold_i             : std_logic;
    signal   gt19_rxdfelfhold_i              : std_logic;
    signal   gt19_rxlpmlfhold_i              : std_logic;
    signal   gt19_rxlpmhfhold_i              : std_logic;


    signal   gt20_txpmaresetdone_i           : std_logic;
    signal   gt20_rxpmaresetdone_i           : std_logic;
    signal   gt20_txresetdone_i              : std_logic;
    signal   gt20_rxresetdone_i              : std_logic;
    signal   gt20_txresetdone_ii             : std_logic;
    signal   gt20_rxresetdone_ii             : std_logic;
    signal   gt20_gttxreset_i                : std_logic;
    signal   gt20_gttxreset_t                : std_logic;
    signal   gt20_gtrxreset_i                : std_logic;
    signal   gt20_gtrxreset_t                : std_logic;
    signal   gt20_txuserrdy_i                : std_logic;
    signal   gt20_txuserrdy_t                : std_logic;
    signal   gt20_rxuserrdy_i                : std_logic;
    signal   gt20_rxuserrdy_t                : std_logic;

    signal   gt20_rxdfeagchold_i             : std_logic;
    signal   gt20_rxdfelfhold_i              : std_logic;
    signal   gt20_rxlpmlfhold_i              : std_logic;
    signal   gt20_rxlpmhfhold_i              : std_logic;


    signal   gt21_txpmaresetdone_i           : std_logic;
    signal   gt21_rxpmaresetdone_i           : std_logic;
    signal   gt21_txresetdone_i              : std_logic;
    signal   gt21_rxresetdone_i              : std_logic;
    signal   gt21_txresetdone_ii             : std_logic;
    signal   gt21_rxresetdone_ii             : std_logic;
    signal   gt21_gttxreset_i                : std_logic;
    signal   gt21_gttxreset_t                : std_logic;
    signal   gt21_gtrxreset_i                : std_logic;
    signal   gt21_gtrxreset_t                : std_logic;
    signal   gt21_txuserrdy_i                : std_logic;
    signal   gt21_txuserrdy_t                : std_logic;
    signal   gt21_rxuserrdy_i                : std_logic;
    signal   gt21_rxuserrdy_t                : std_logic;

    signal   gt21_rxdfeagchold_i             : std_logic;
    signal   gt21_rxdfelfhold_i              : std_logic;
    signal   gt21_rxlpmlfhold_i              : std_logic;
    signal   gt21_rxlpmhfhold_i              : std_logic;


    signal   gt22_txpmaresetdone_i           : std_logic;
    signal   gt22_rxpmaresetdone_i           : std_logic;
    signal   gt22_txresetdone_i              : std_logic;
    signal   gt22_rxresetdone_i              : std_logic;
    signal   gt22_txresetdone_ii             : std_logic;
    signal   gt22_rxresetdone_ii             : std_logic;
    signal   gt22_gttxreset_i                : std_logic;
    signal   gt22_gttxreset_t                : std_logic;
    signal   gt22_gtrxreset_i                : std_logic;
    signal   gt22_gtrxreset_t                : std_logic;
    signal   gt22_txuserrdy_i                : std_logic;
    signal   gt22_txuserrdy_t                : std_logic;
    signal   gt22_rxuserrdy_i                : std_logic;
    signal   gt22_rxuserrdy_t                : std_logic;

    signal   gt22_rxdfeagchold_i             : std_logic;
    signal   gt22_rxdfelfhold_i              : std_logic;
    signal   gt22_rxlpmlfhold_i              : std_logic;
    signal   gt22_rxlpmhfhold_i              : std_logic;


    signal   gt23_txpmaresetdone_i           : std_logic;
    signal   gt23_rxpmaresetdone_i           : std_logic;
    signal   gt23_txresetdone_i              : std_logic;
    signal   gt23_rxresetdone_i              : std_logic;
    signal   gt23_txresetdone_ii             : std_logic;
    signal   gt23_rxresetdone_ii             : std_logic;
    signal   gt23_gttxreset_i                : std_logic;
    signal   gt23_gttxreset_t                : std_logic;
    signal   gt23_gtrxreset_i                : std_logic;
    signal   gt23_gtrxreset_t                : std_logic;
    signal   gt23_txuserrdy_i                : std_logic;
    signal   gt23_txuserrdy_t                : std_logic;
    signal   gt23_rxuserrdy_i                : std_logic;
    signal   gt23_rxuserrdy_t                : std_logic;

    signal   gt23_rxdfeagchold_i             : std_logic;
    signal   gt23_rxdfelfhold_i              : std_logic;
    signal   gt23_rxlpmlfhold_i              : std_logic;
    signal   gt23_rxlpmhfhold_i              : std_logic;


    signal   gt24_txpmaresetdone_i           : std_logic;
    signal   gt24_rxpmaresetdone_i           : std_logic;
    signal   gt24_txresetdone_i              : std_logic;
    signal   gt24_rxresetdone_i              : std_logic;
    signal   gt24_txresetdone_ii             : std_logic;
    signal   gt24_rxresetdone_ii             : std_logic;
    signal   gt24_gttxreset_i                : std_logic;
    signal   gt24_gttxreset_t                : std_logic;
    signal   gt24_gtrxreset_i                : std_logic;
    signal   gt24_gtrxreset_t                : std_logic;
    signal   gt24_txuserrdy_i                : std_logic;
    signal   gt24_txuserrdy_t                : std_logic;
    signal   gt24_rxuserrdy_i                : std_logic;
    signal   gt24_rxuserrdy_t                : std_logic;

    signal   gt24_rxdfeagchold_i             : std_logic;
    signal   gt24_rxdfelfhold_i              : std_logic;
    signal   gt24_rxlpmlfhold_i              : std_logic;
    signal   gt24_rxlpmhfhold_i              : std_logic;


    signal   gt25_txpmaresetdone_i           : std_logic;
    signal   gt25_rxpmaresetdone_i           : std_logic;
    signal   gt25_txresetdone_i              : std_logic;
    signal   gt25_rxresetdone_i              : std_logic;
    signal   gt25_txresetdone_ii             : std_logic;
    signal   gt25_rxresetdone_ii             : std_logic;
    signal   gt25_gttxreset_i                : std_logic;
    signal   gt25_gttxreset_t                : std_logic;
    signal   gt25_gtrxreset_i                : std_logic;
    signal   gt25_gtrxreset_t                : std_logic;
    signal   gt25_txuserrdy_i                : std_logic;
    signal   gt25_txuserrdy_t                : std_logic;
    signal   gt25_rxuserrdy_i                : std_logic;
    signal   gt25_rxuserrdy_t                : std_logic;

    signal   gt25_rxdfeagchold_i             : std_logic;
    signal   gt25_rxdfelfhold_i              : std_logic;
    signal   gt25_rxlpmlfhold_i              : std_logic;
    signal   gt25_rxlpmhfhold_i              : std_logic;


    signal   gt26_txpmaresetdone_i           : std_logic;
    signal   gt26_rxpmaresetdone_i           : std_logic;
    signal   gt26_txresetdone_i              : std_logic;
    signal   gt26_rxresetdone_i              : std_logic;
    signal   gt26_txresetdone_ii             : std_logic;
    signal   gt26_rxresetdone_ii             : std_logic;
    signal   gt26_gttxreset_i                : std_logic;
    signal   gt26_gttxreset_t                : std_logic;
    signal   gt26_gtrxreset_i                : std_logic;
    signal   gt26_gtrxreset_t                : std_logic;
    signal   gt26_txuserrdy_i                : std_logic;
    signal   gt26_txuserrdy_t                : std_logic;
    signal   gt26_rxuserrdy_i                : std_logic;
    signal   gt26_rxuserrdy_t                : std_logic;

    signal   gt26_rxdfeagchold_i             : std_logic;
    signal   gt26_rxdfelfhold_i              : std_logic;
    signal   gt26_rxlpmlfhold_i              : std_logic;
    signal   gt26_rxlpmhfhold_i              : std_logic;


    signal   gt27_txpmaresetdone_i           : std_logic;
    signal   gt27_rxpmaresetdone_i           : std_logic;
    signal   gt27_txresetdone_i              : std_logic;
    signal   gt27_rxresetdone_i              : std_logic;
    signal   gt27_txresetdone_ii             : std_logic;
    signal   gt27_rxresetdone_ii             : std_logic;
    signal   gt27_gttxreset_i                : std_logic;
    signal   gt27_gttxreset_t                : std_logic;
    signal   gt27_gtrxreset_i                : std_logic;
    signal   gt27_gtrxreset_t                : std_logic;
    signal   gt27_txuserrdy_i                : std_logic;
    signal   gt27_txuserrdy_t                : std_logic;
    signal   gt27_rxuserrdy_i                : std_logic;
    signal   gt27_rxuserrdy_t                : std_logic;

    signal   gt27_rxdfeagchold_i             : std_logic;
    signal   gt27_rxdfelfhold_i              : std_logic;
    signal   gt27_rxlpmlfhold_i              : std_logic;
    signal   gt27_rxlpmhfhold_i              : std_logic;


    signal   gt28_txpmaresetdone_i           : std_logic;
    signal   gt28_rxpmaresetdone_i           : std_logic;
    signal   gt28_txresetdone_i              : std_logic;
    signal   gt28_rxresetdone_i              : std_logic;
    signal   gt28_txresetdone_ii             : std_logic;
    signal   gt28_rxresetdone_ii             : std_logic;
    signal   gt28_gttxreset_i                : std_logic;
    signal   gt28_gttxreset_t                : std_logic;
    signal   gt28_gtrxreset_i                : std_logic;
    signal   gt28_gtrxreset_t                : std_logic;
    signal   gt28_txuserrdy_i                : std_logic;
    signal   gt28_txuserrdy_t                : std_logic;
    signal   gt28_rxuserrdy_i                : std_logic;
    signal   gt28_rxuserrdy_t                : std_logic;

    signal   gt28_rxdfeagchold_i             : std_logic;
    signal   gt28_rxdfelfhold_i              : std_logic;
    signal   gt28_rxlpmlfhold_i              : std_logic;
    signal   gt28_rxlpmhfhold_i              : std_logic;


    signal   gt29_txpmaresetdone_i           : std_logic;
    signal   gt29_rxpmaresetdone_i           : std_logic;
    signal   gt29_txresetdone_i              : std_logic;
    signal   gt29_rxresetdone_i              : std_logic;
    signal   gt29_txresetdone_ii             : std_logic;
    signal   gt29_rxresetdone_ii             : std_logic;
    signal   gt29_gttxreset_i                : std_logic;
    signal   gt29_gttxreset_t                : std_logic;
    signal   gt29_gtrxreset_i                : std_logic;
    signal   gt29_gtrxreset_t                : std_logic;
    signal   gt29_txuserrdy_i                : std_logic;
    signal   gt29_txuserrdy_t                : std_logic;
    signal   gt29_rxuserrdy_i                : std_logic;
    signal   gt29_rxuserrdy_t                : std_logic;

    signal   gt29_rxdfeagchold_i             : std_logic;
    signal   gt29_rxdfelfhold_i              : std_logic;
    signal   gt29_rxlpmlfhold_i              : std_logic;
    signal   gt29_rxlpmhfhold_i              : std_logic;


    signal   gt30_txpmaresetdone_i           : std_logic;
    signal   gt30_rxpmaresetdone_i           : std_logic;
    signal   gt30_txresetdone_i              : std_logic;
    signal   gt30_rxresetdone_i              : std_logic;
    signal   gt30_txresetdone_ii             : std_logic;
    signal   gt30_rxresetdone_ii             : std_logic;
    signal   gt30_gttxreset_i                : std_logic;
    signal   gt30_gttxreset_t                : std_logic;
    signal   gt30_gtrxreset_i                : std_logic;
    signal   gt30_gtrxreset_t                : std_logic;
    signal   gt30_txuserrdy_i                : std_logic;
    signal   gt30_txuserrdy_t                : std_logic;
    signal   gt30_rxuserrdy_i                : std_logic;
    signal   gt30_rxuserrdy_t                : std_logic;

    signal   gt30_rxdfeagchold_i             : std_logic;
    signal   gt30_rxdfelfhold_i              : std_logic;
    signal   gt30_rxlpmlfhold_i              : std_logic;
    signal   gt30_rxlpmhfhold_i              : std_logic;


    signal   gt31_txpmaresetdone_i           : std_logic;
    signal   gt31_rxpmaresetdone_i           : std_logic;
    signal   gt31_txresetdone_i              : std_logic;
    signal   gt31_rxresetdone_i              : std_logic;
    signal   gt31_txresetdone_ii             : std_logic;
    signal   gt31_rxresetdone_ii             : std_logic;
    signal   gt31_gttxreset_i                : std_logic;
    signal   gt31_gttxreset_t                : std_logic;
    signal   gt31_gtrxreset_i                : std_logic;
    signal   gt31_gtrxreset_t                : std_logic;
    signal   gt31_txuserrdy_i                : std_logic;
    signal   gt31_txuserrdy_t                : std_logic;
    signal   gt31_rxuserrdy_i                : std_logic;
    signal   gt31_rxuserrdy_t                : std_logic;

    signal   gt31_rxdfeagchold_i             : std_logic;
    signal   gt31_rxdfelfhold_i              : std_logic;
    signal   gt31_rxlpmlfhold_i              : std_logic;
    signal   gt31_rxlpmhfhold_i              : std_logic;



    signal   gt0_qpllreset_i                 : std_logic;
    signal   gt0_qpllreset_t                 : std_logic;
    signal   gt0_qpllrefclklost_i            : std_logic;
    signal   gt0_qplllock_i                  : std_logic;
    signal   gt1_qpllreset_i                 : std_logic;
    signal   gt1_qpllreset_t                 : std_logic;
    signal   gt1_qpllrefclklost_i            : std_logic;
    signal   gt1_qplllock_i                  : std_logic;
    signal   gt2_qpllreset_i                 : std_logic;
    signal   gt2_qpllreset_t                 : std_logic;
    signal   gt2_qpllrefclklost_i            : std_logic;
    signal   gt2_qplllock_i                  : std_logic;
    signal   gt3_qpllreset_i                 : std_logic;
    signal   gt3_qpllreset_t                 : std_logic;
    signal   gt3_qpllrefclklost_i            : std_logic;
    signal   gt3_qplllock_i                  : std_logic;
    signal   gt4_qpllreset_i                 : std_logic;
    signal   gt4_qpllreset_t                 : std_logic;
    signal   gt4_qpllrefclklost_i            : std_logic;
    signal   gt4_qplllock_i                  : std_logic;
    signal   gt5_qpllreset_i                 : std_logic;
    signal   gt5_qpllreset_t                 : std_logic;
    signal   gt5_qpllrefclklost_i            : std_logic;
    signal   gt5_qplllock_i                  : std_logic;
    signal   gt6_qpllreset_i                 : std_logic;
    signal   gt6_qpllreset_t                 : std_logic;
    signal   gt6_qpllrefclklost_i            : std_logic;
    signal   gt6_qplllock_i                  : std_logic;
    signal   gt7_qpllreset_i                 : std_logic;
    signal   gt7_qpllreset_t                 : std_logic;
    signal   gt7_qpllrefclklost_i            : std_logic;
    signal   gt7_qplllock_i                  : std_logic;


    ------------------------------- Global Signals -----------------------------
    signal  tied_to_ground_i                : std_logic;
    signal  tied_to_vcc_i                   : std_logic;
    signal   gt0_txphaligndone_i             : std_logic;
    signal   gt0_txdlysreset_i               : std_logic;
    signal   gt0_txdlysresetdone_i           : std_logic;
    signal   gt0_txphdlyreset_i              : std_logic;
    signal   gt0_txphalignen_i               : std_logic;
    signal   gt0_txdlyen_i                   : std_logic;
    signal   gt0_txphalign_i                 : std_logic;
    signal   gt0_txphinit_i                  : std_logic;
    signal   gt0_txphinitdone_i              : std_logic;
    signal   gt0_run_tx_phalignment_i        : std_logic;
    signal   gt0_rst_tx_phalignment_i        : std_logic;
    signal   gt0_tx_phalignment_done_i       : std_logic;
    signal   gt0_txsyncallin_i               : std_logic;
    signal   gt0_txsyncin_i                  : std_logic;
    signal   gt0_txsyncmode_i                : std_logic;
    signal   gt0_txsyncout_i                 : std_logic;
    signal   gt0_txsyncdone_i                : std_logic;

    signal   gt0_txoutclk_i                  : std_logic;
    signal   gt0_rxoutclk_i                  : std_logic;
    signal   gt0_rxoutclk_i2                 : std_logic;
    signal   gt0_txoutclk_i2                 : std_logic;
    signal   gt0_recclk_stable_i             : std_logic;
    signal   gt0_rx_cdrlocked                : std_logic;
    signal   gt0_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt0_rxphaligndone_i             : std_logic;
    signal   gt0_rxdlysreset_i               : std_logic;
    signal   gt0_rxdlysresetdone_i           : std_logic;
    signal   gt0_rxphdlyreset_i              : std_logic;
    signal   gt0_rxphalignen_i               : std_logic;
    signal   gt0_rxdlyen_i                   : std_logic;
    signal   gt0_rxphalign_i                 : std_logic;
    signal   gt0_run_rx_phalignment_i        : std_logic;
    signal   gt0_rst_rx_phalignment_i        : std_logic;
    signal   gt0_rx_phalignment_done_i       : std_logic;
    signal   gt0_rxsyncallin_i               : std_logic;
    signal   gt0_rxsyncin_i                  : std_logic;
    signal   gt0_rxsyncmode_i                : std_logic;
    signal   gt0_rxsyncout_i                 : std_logic;
    signal   gt0_rxsyncdone_i                : std_logic;
    signal   gt1_txphaligndone_i             : std_logic;
    signal   gt1_txdlysreset_i               : std_logic;
    signal   gt1_txdlysresetdone_i           : std_logic;
    signal   gt1_txphdlyreset_i              : std_logic;
    signal   gt1_txphalignen_i               : std_logic;
    signal   gt1_txdlyen_i                   : std_logic;
    signal   gt1_txphalign_i                 : std_logic;
    signal   gt1_txphinit_i                  : std_logic;
    signal   gt1_txphinitdone_i              : std_logic;
    signal   gt1_run_tx_phalignment_i        : std_logic;
    signal   gt1_rst_tx_phalignment_i        : std_logic;
    signal   gt1_tx_phalignment_done_i       : std_logic;
    signal   gt1_txsyncallin_i               : std_logic;
    signal   gt1_txsyncin_i                  : std_logic;
    signal   gt1_txsyncmode_i                : std_logic;
    signal   gt1_txsyncout_i                 : std_logic;
    signal   gt1_txsyncdone_i                : std_logic;

    signal   gt1_txoutclk_i                  : std_logic;
    signal   gt1_rxoutclk_i                  : std_logic;
    signal   gt1_rxoutclk_i2                 : std_logic;
    signal   gt1_txoutclk_i2                 : std_logic;
    signal   gt1_recclk_stable_i             : std_logic;
    signal   gt1_rx_cdrlocked                : std_logic;
    signal   gt1_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt1_rxphaligndone_i             : std_logic;
    signal   gt1_rxdlysreset_i               : std_logic;
    signal   gt1_rxdlysresetdone_i           : std_logic;
    signal   gt1_rxphdlyreset_i              : std_logic;
    signal   gt1_rxphalignen_i               : std_logic;
    signal   gt1_rxdlyen_i                   : std_logic;
    signal   gt1_rxphalign_i                 : std_logic;
    signal   gt1_run_rx_phalignment_i        : std_logic;
    signal   gt1_rst_rx_phalignment_i        : std_logic;
    signal   gt1_rx_phalignment_done_i       : std_logic;
    signal   gt1_rxsyncallin_i               : std_logic;
    signal   gt1_rxsyncin_i                  : std_logic;
    signal   gt1_rxsyncmode_i                : std_logic;
    signal   gt1_rxsyncout_i                 : std_logic;
    signal   gt1_rxsyncdone_i                : std_logic;
    signal   gt2_txphaligndone_i             : std_logic;
    signal   gt2_txdlysreset_i               : std_logic;
    signal   gt2_txdlysresetdone_i           : std_logic;
    signal   gt2_txphdlyreset_i              : std_logic;
    signal   gt2_txphalignen_i               : std_logic;
    signal   gt2_txdlyen_i                   : std_logic;
    signal   gt2_txphalign_i                 : std_logic;
    signal   gt2_txphinit_i                  : std_logic;
    signal   gt2_txphinitdone_i              : std_logic;
    signal   gt2_run_tx_phalignment_i        : std_logic;
    signal   gt2_rst_tx_phalignment_i        : std_logic;
    signal   gt2_tx_phalignment_done_i       : std_logic;
    signal   gt2_txsyncallin_i               : std_logic;
    signal   gt2_txsyncin_i                  : std_logic;
    signal   gt2_txsyncmode_i                : std_logic;
    signal   gt2_txsyncout_i                 : std_logic;
    signal   gt2_txsyncdone_i                : std_logic;

    signal   gt2_txoutclk_i                  : std_logic;
    signal   gt2_rxoutclk_i                  : std_logic;
    signal   gt2_rxoutclk_i2                 : std_logic;
    signal   gt2_txoutclk_i2                 : std_logic;
    signal   gt2_recclk_stable_i             : std_logic;
    signal   gt2_rx_cdrlocked                : std_logic;
    signal   gt2_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt2_rxphaligndone_i             : std_logic;
    signal   gt2_rxdlysreset_i               : std_logic;
    signal   gt2_rxdlysresetdone_i           : std_logic;
    signal   gt2_rxphdlyreset_i              : std_logic;
    signal   gt2_rxphalignen_i               : std_logic;
    signal   gt2_rxdlyen_i                   : std_logic;
    signal   gt2_rxphalign_i                 : std_logic;
    signal   gt2_run_rx_phalignment_i        : std_logic;
    signal   gt2_rst_rx_phalignment_i        : std_logic;
    signal   gt2_rx_phalignment_done_i       : std_logic;
    signal   gt2_rxsyncallin_i               : std_logic;
    signal   gt2_rxsyncin_i                  : std_logic;
    signal   gt2_rxsyncmode_i                : std_logic;
    signal   gt2_rxsyncout_i                 : std_logic;
    signal   gt2_rxsyncdone_i                : std_logic;
    signal   gt3_txphaligndone_i             : std_logic;
    signal   gt3_txdlysreset_i               : std_logic;
    signal   gt3_txdlysresetdone_i           : std_logic;
    signal   gt3_txphdlyreset_i              : std_logic;
    signal   gt3_txphalignen_i               : std_logic;
    signal   gt3_txdlyen_i                   : std_logic;
    signal   gt3_txphalign_i                 : std_logic;
    signal   gt3_txphinit_i                  : std_logic;
    signal   gt3_txphinitdone_i              : std_logic;
    signal   gt3_run_tx_phalignment_i        : std_logic;
    signal   gt3_rst_tx_phalignment_i        : std_logic;
    signal   gt3_tx_phalignment_done_i       : std_logic;
    signal   gt3_txsyncallin_i               : std_logic;
    signal   gt3_txsyncin_i                  : std_logic;
    signal   gt3_txsyncmode_i                : std_logic;
    signal   gt3_txsyncout_i                 : std_logic;
    signal   gt3_txsyncdone_i                : std_logic;

    signal   gt3_txoutclk_i                  : std_logic;
    signal   gt3_rxoutclk_i                  : std_logic;
    signal   gt3_rxoutclk_i2                 : std_logic;
    signal   gt3_txoutclk_i2                 : std_logic;
    signal   gt3_recclk_stable_i             : std_logic;
    signal   gt3_rx_cdrlocked                : std_logic;
    signal   gt3_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt3_rxphaligndone_i             : std_logic;
    signal   gt3_rxdlysreset_i               : std_logic;
    signal   gt3_rxdlysresetdone_i           : std_logic;
    signal   gt3_rxphdlyreset_i              : std_logic;
    signal   gt3_rxphalignen_i               : std_logic;
    signal   gt3_rxdlyen_i                   : std_logic;
    signal   gt3_rxphalign_i                 : std_logic;
    signal   gt3_run_rx_phalignment_i        : std_logic;
    signal   gt3_rst_rx_phalignment_i        : std_logic;
    signal   gt3_rx_phalignment_done_i       : std_logic;
    signal   gt3_rxsyncallin_i               : std_logic;
    signal   gt3_rxsyncin_i                  : std_logic;
    signal   gt3_rxsyncmode_i                : std_logic;
    signal   gt3_rxsyncout_i                 : std_logic;
    signal   gt3_rxsyncdone_i                : std_logic;
    signal   gt4_txphaligndone_i             : std_logic;
    signal   gt4_txdlysreset_i               : std_logic;
    signal   gt4_txdlysresetdone_i           : std_logic;
    signal   gt4_txphdlyreset_i              : std_logic;
    signal   gt4_txphalignen_i               : std_logic;
    signal   gt4_txdlyen_i                   : std_logic;
    signal   gt4_txphalign_i                 : std_logic;
    signal   gt4_txphinit_i                  : std_logic;
    signal   gt4_txphinitdone_i              : std_logic;
    signal   gt4_run_tx_phalignment_i        : std_logic;
    signal   gt4_rst_tx_phalignment_i        : std_logic;
    signal   gt4_tx_phalignment_done_i       : std_logic;
    signal   gt4_txsyncallin_i               : std_logic;
    signal   gt4_txsyncin_i                  : std_logic;
    signal   gt4_txsyncmode_i                : std_logic;
    signal   gt4_txsyncout_i                 : std_logic;
    signal   gt4_txsyncdone_i                : std_logic;

    signal   gt4_txoutclk_i                  : std_logic;
    signal   gt4_rxoutclk_i                  : std_logic;
    signal   gt4_rxoutclk_i2                 : std_logic;
    signal   gt4_txoutclk_i2                 : std_logic;
    signal   gt4_recclk_stable_i             : std_logic;
    signal   gt4_rx_cdrlocked                : std_logic;
    signal   gt4_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt4_rxphaligndone_i             : std_logic;
    signal   gt4_rxdlysreset_i               : std_logic;
    signal   gt4_rxdlysresetdone_i           : std_logic;
    signal   gt4_rxphdlyreset_i              : std_logic;
    signal   gt4_rxphalignen_i               : std_logic;
    signal   gt4_rxdlyen_i                   : std_logic;
    signal   gt4_rxphalign_i                 : std_logic;
    signal   gt4_run_rx_phalignment_i        : std_logic;
    signal   gt4_rst_rx_phalignment_i        : std_logic;
    signal   gt4_rx_phalignment_done_i       : std_logic;
    signal   gt4_rxsyncallin_i               : std_logic;
    signal   gt4_rxsyncin_i                  : std_logic;
    signal   gt4_rxsyncmode_i                : std_logic;
    signal   gt4_rxsyncout_i                 : std_logic;
    signal   gt4_rxsyncdone_i                : std_logic;
    signal   gt5_txphaligndone_i             : std_logic;
    signal   gt5_txdlysreset_i               : std_logic;
    signal   gt5_txdlysresetdone_i           : std_logic;
    signal   gt5_txphdlyreset_i              : std_logic;
    signal   gt5_txphalignen_i               : std_logic;
    signal   gt5_txdlyen_i                   : std_logic;
    signal   gt5_txphalign_i                 : std_logic;
    signal   gt5_txphinit_i                  : std_logic;
    signal   gt5_txphinitdone_i              : std_logic;
    signal   gt5_run_tx_phalignment_i        : std_logic;
    signal   gt5_rst_tx_phalignment_i        : std_logic;
    signal   gt5_tx_phalignment_done_i       : std_logic;
    signal   gt5_txsyncallin_i               : std_logic;
    signal   gt5_txsyncin_i                  : std_logic;
    signal   gt5_txsyncmode_i                : std_logic;
    signal   gt5_txsyncout_i                 : std_logic;
    signal   gt5_txsyncdone_i                : std_logic;

    signal   gt5_txoutclk_i                  : std_logic;
    signal   gt5_rxoutclk_i                  : std_logic;
    signal   gt5_rxoutclk_i2                 : std_logic;
    signal   gt5_txoutclk_i2                 : std_logic;
    signal   gt5_recclk_stable_i             : std_logic;
    signal   gt5_rx_cdrlocked                : std_logic;
    signal   gt5_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt5_rxphaligndone_i             : std_logic;
    signal   gt5_rxdlysreset_i               : std_logic;
    signal   gt5_rxdlysresetdone_i           : std_logic;
    signal   gt5_rxphdlyreset_i              : std_logic;
    signal   gt5_rxphalignen_i               : std_logic;
    signal   gt5_rxdlyen_i                   : std_logic;
    signal   gt5_rxphalign_i                 : std_logic;
    signal   gt5_run_rx_phalignment_i        : std_logic;
    signal   gt5_rst_rx_phalignment_i        : std_logic;
    signal   gt5_rx_phalignment_done_i       : std_logic;
    signal   gt5_rxsyncallin_i               : std_logic;
    signal   gt5_rxsyncin_i                  : std_logic;
    signal   gt5_rxsyncmode_i                : std_logic;
    signal   gt5_rxsyncout_i                 : std_logic;
    signal   gt5_rxsyncdone_i                : std_logic;
    signal   gt6_txphaligndone_i             : std_logic;
    signal   gt6_txdlysreset_i               : std_logic;
    signal   gt6_txdlysresetdone_i           : std_logic;
    signal   gt6_txphdlyreset_i              : std_logic;
    signal   gt6_txphalignen_i               : std_logic;
    signal   gt6_txdlyen_i                   : std_logic;
    signal   gt6_txphalign_i                 : std_logic;
    signal   gt6_txphinit_i                  : std_logic;
    signal   gt6_txphinitdone_i              : std_logic;
    signal   gt6_run_tx_phalignment_i        : std_logic;
    signal   gt6_rst_tx_phalignment_i        : std_logic;
    signal   gt6_tx_phalignment_done_i       : std_logic;
    signal   gt6_txsyncallin_i               : std_logic;
    signal   gt6_txsyncin_i                  : std_logic;
    signal   gt6_txsyncmode_i                : std_logic;
    signal   gt6_txsyncout_i                 : std_logic;
    signal   gt6_txsyncdone_i                : std_logic;

    signal   gt6_txoutclk_i                  : std_logic;
    signal   gt6_rxoutclk_i                  : std_logic;
    signal   gt6_rxoutclk_i2                 : std_logic;
    signal   gt6_txoutclk_i2                 : std_logic;
    signal   gt6_recclk_stable_i             : std_logic;
    signal   gt6_rx_cdrlocked                : std_logic;
    signal   gt6_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt6_rxphaligndone_i             : std_logic;
    signal   gt6_rxdlysreset_i               : std_logic;
    signal   gt6_rxdlysresetdone_i           : std_logic;
    signal   gt6_rxphdlyreset_i              : std_logic;
    signal   gt6_rxphalignen_i               : std_logic;
    signal   gt6_rxdlyen_i                   : std_logic;
    signal   gt6_rxphalign_i                 : std_logic;
    signal   gt6_run_rx_phalignment_i        : std_logic;
    signal   gt6_rst_rx_phalignment_i        : std_logic;
    signal   gt6_rx_phalignment_done_i       : std_logic;
    signal   gt6_rxsyncallin_i               : std_logic;
    signal   gt6_rxsyncin_i                  : std_logic;
    signal   gt6_rxsyncmode_i                : std_logic;
    signal   gt6_rxsyncout_i                 : std_logic;
    signal   gt6_rxsyncdone_i                : std_logic;
    signal   gt7_txphaligndone_i             : std_logic;
    signal   gt7_txdlysreset_i               : std_logic;
    signal   gt7_txdlysresetdone_i           : std_logic;
    signal   gt7_txphdlyreset_i              : std_logic;
    signal   gt7_txphalignen_i               : std_logic;
    signal   gt7_txdlyen_i                   : std_logic;
    signal   gt7_txphalign_i                 : std_logic;
    signal   gt7_txphinit_i                  : std_logic;
    signal   gt7_txphinitdone_i              : std_logic;
    signal   gt7_run_tx_phalignment_i        : std_logic;
    signal   gt7_rst_tx_phalignment_i        : std_logic;
    signal   gt7_tx_phalignment_done_i       : std_logic;
    signal   gt7_txsyncallin_i               : std_logic;
    signal   gt7_txsyncin_i                  : std_logic;
    signal   gt7_txsyncmode_i                : std_logic;
    signal   gt7_txsyncout_i                 : std_logic;
    signal   gt7_txsyncdone_i                : std_logic;

    signal   gt7_txoutclk_i                  : std_logic;
    signal   gt7_rxoutclk_i                  : std_logic;
    signal   gt7_rxoutclk_i2                 : std_logic;
    signal   gt7_txoutclk_i2                 : std_logic;
    signal   gt7_recclk_stable_i             : std_logic;
    signal   gt7_rx_cdrlocked                : std_logic;
    signal   gt7_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt7_rxphaligndone_i             : std_logic;
    signal   gt7_rxdlysreset_i               : std_logic;
    signal   gt7_rxdlysresetdone_i           : std_logic;
    signal   gt7_rxphdlyreset_i              : std_logic;
    signal   gt7_rxphalignen_i               : std_logic;
    signal   gt7_rxdlyen_i                   : std_logic;
    signal   gt7_rxphalign_i                 : std_logic;
    signal   gt7_run_rx_phalignment_i        : std_logic;
    signal   gt7_rst_rx_phalignment_i        : std_logic;
    signal   gt7_rx_phalignment_done_i       : std_logic;
    signal   gt7_rxsyncallin_i               : std_logic;
    signal   gt7_rxsyncin_i                  : std_logic;
    signal   gt7_rxsyncmode_i                : std_logic;
    signal   gt7_rxsyncout_i                 : std_logic;
    signal   gt7_rxsyncdone_i                : std_logic;
    signal   gt8_txphaligndone_i             : std_logic;
    signal   gt8_txdlysreset_i               : std_logic;
    signal   gt8_txdlysresetdone_i           : std_logic;
    signal   gt8_txphdlyreset_i              : std_logic;
    signal   gt8_txphalignen_i               : std_logic;
    signal   gt8_txdlyen_i                   : std_logic;
    signal   gt8_txphalign_i                 : std_logic;
    signal   gt8_txphinit_i                  : std_logic;
    signal   gt8_txphinitdone_i              : std_logic;
    signal   gt8_run_tx_phalignment_i        : std_logic;
    signal   gt8_rst_tx_phalignment_i        : std_logic;
    signal   gt8_tx_phalignment_done_i       : std_logic;
    signal   gt8_txsyncallin_i               : std_logic;
    signal   gt8_txsyncin_i                  : std_logic;
    signal   gt8_txsyncmode_i                : std_logic;
    signal   gt8_txsyncout_i                 : std_logic;
    signal   gt8_txsyncdone_i                : std_logic;

    signal   gt8_txoutclk_i                  : std_logic;
    signal   gt8_rxoutclk_i                  : std_logic;
    signal   gt8_rxoutclk_i2                 : std_logic;
    signal   gt8_txoutclk_i2                 : std_logic;
    signal   gt8_recclk_stable_i             : std_logic;
    signal   gt8_rx_cdrlocked                : std_logic;
    signal   gt8_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt8_rxphaligndone_i             : std_logic;
    signal   gt8_rxdlysreset_i               : std_logic;
    signal   gt8_rxdlysresetdone_i           : std_logic;
    signal   gt8_rxphdlyreset_i              : std_logic;
    signal   gt8_rxphalignen_i               : std_logic;
    signal   gt8_rxdlyen_i                   : std_logic;
    signal   gt8_rxphalign_i                 : std_logic;
    signal   gt8_run_rx_phalignment_i        : std_logic;
    signal   gt8_rst_rx_phalignment_i        : std_logic;
    signal   gt8_rx_phalignment_done_i       : std_logic;
    signal   gt8_rxsyncallin_i               : std_logic;
    signal   gt8_rxsyncin_i                  : std_logic;
    signal   gt8_rxsyncmode_i                : std_logic;
    signal   gt8_rxsyncout_i                 : std_logic;
    signal   gt8_rxsyncdone_i                : std_logic;
    signal   gt9_txphaligndone_i             : std_logic;
    signal   gt9_txdlysreset_i               : std_logic;
    signal   gt9_txdlysresetdone_i           : std_logic;
    signal   gt9_txphdlyreset_i              : std_logic;
    signal   gt9_txphalignen_i               : std_logic;
    signal   gt9_txdlyen_i                   : std_logic;
    signal   gt9_txphalign_i                 : std_logic;
    signal   gt9_txphinit_i                  : std_logic;
    signal   gt9_txphinitdone_i              : std_logic;
    signal   gt9_run_tx_phalignment_i        : std_logic;
    signal   gt9_rst_tx_phalignment_i        : std_logic;
    signal   gt9_tx_phalignment_done_i       : std_logic;
    signal   gt9_txsyncallin_i               : std_logic;
    signal   gt9_txsyncin_i                  : std_logic;
    signal   gt9_txsyncmode_i                : std_logic;
    signal   gt9_txsyncout_i                 : std_logic;
    signal   gt9_txsyncdone_i                : std_logic;

    signal   gt9_txoutclk_i                  : std_logic;
    signal   gt9_rxoutclk_i                  : std_logic;
    signal   gt9_rxoutclk_i2                 : std_logic;
    signal   gt9_txoutclk_i2                 : std_logic;
    signal   gt9_recclk_stable_i             : std_logic;
    signal   gt9_rx_cdrlocked                : std_logic;
    signal   gt9_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt9_rxphaligndone_i             : std_logic;
    signal   gt9_rxdlysreset_i               : std_logic;
    signal   gt9_rxdlysresetdone_i           : std_logic;
    signal   gt9_rxphdlyreset_i              : std_logic;
    signal   gt9_rxphalignen_i               : std_logic;
    signal   gt9_rxdlyen_i                   : std_logic;
    signal   gt9_rxphalign_i                 : std_logic;
    signal   gt9_run_rx_phalignment_i        : std_logic;
    signal   gt9_rst_rx_phalignment_i        : std_logic;
    signal   gt9_rx_phalignment_done_i       : std_logic;
    signal   gt9_rxsyncallin_i               : std_logic;
    signal   gt9_rxsyncin_i                  : std_logic;
    signal   gt9_rxsyncmode_i                : std_logic;
    signal   gt9_rxsyncout_i                 : std_logic;
    signal   gt9_rxsyncdone_i                : std_logic;
    signal   gt10_txphaligndone_i            : std_logic;
    signal   gt10_txdlysreset_i              : std_logic;
    signal   gt10_txdlysresetdone_i          : std_logic;
    signal   gt10_txphdlyreset_i             : std_logic;
    signal   gt10_txphalignen_i              : std_logic;
    signal   gt10_txdlyen_i                  : std_logic;
    signal   gt10_txphalign_i                : std_logic;
    signal   gt10_txphinit_i                 : std_logic;
    signal   gt10_txphinitdone_i             : std_logic;
    signal   gt10_run_tx_phalignment_i       : std_logic;
    signal   gt10_rst_tx_phalignment_i       : std_logic;
    signal   gt10_tx_phalignment_done_i      : std_logic;
    signal   gt10_txsyncallin_i              : std_logic;
    signal   gt10_txsyncin_i                 : std_logic;
    signal   gt10_txsyncmode_i               : std_logic;
    signal   gt10_txsyncout_i                : std_logic;
    signal   gt10_txsyncdone_i               : std_logic;

    signal   gt10_txoutclk_i                 : std_logic;
    signal   gt10_rxoutclk_i                 : std_logic;
    signal   gt10_rxoutclk_i2                : std_logic;
    signal   gt10_txoutclk_i2                : std_logic;
    signal   gt10_recclk_stable_i            : std_logic;
    signal   gt10_rx_cdrlocked               : std_logic;
    signal   gt10_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt10_rxphaligndone_i            : std_logic;
    signal   gt10_rxdlysreset_i              : std_logic;
    signal   gt10_rxdlysresetdone_i          : std_logic;
    signal   gt10_rxphdlyreset_i             : std_logic;
    signal   gt10_rxphalignen_i              : std_logic;
    signal   gt10_rxdlyen_i                  : std_logic;
    signal   gt10_rxphalign_i                : std_logic;
    signal   gt10_run_rx_phalignment_i       : std_logic;
    signal   gt10_rst_rx_phalignment_i       : std_logic;
    signal   gt10_rx_phalignment_done_i      : std_logic;
    signal   gt10_rxsyncallin_i              : std_logic;
    signal   gt10_rxsyncin_i                 : std_logic;
    signal   gt10_rxsyncmode_i               : std_logic;
    signal   gt10_rxsyncout_i                : std_logic;
    signal   gt10_rxsyncdone_i               : std_logic;
    signal   gt11_txphaligndone_i            : std_logic;
    signal   gt11_txdlysreset_i              : std_logic;
    signal   gt11_txdlysresetdone_i          : std_logic;
    signal   gt11_txphdlyreset_i             : std_logic;
    signal   gt11_txphalignen_i              : std_logic;
    signal   gt11_txdlyen_i                  : std_logic;
    signal   gt11_txphalign_i                : std_logic;
    signal   gt11_txphinit_i                 : std_logic;
    signal   gt11_txphinitdone_i             : std_logic;
    signal   gt11_run_tx_phalignment_i       : std_logic;
    signal   gt11_rst_tx_phalignment_i       : std_logic;
    signal   gt11_tx_phalignment_done_i      : std_logic;
    signal   gt11_txsyncallin_i              : std_logic;
    signal   gt11_txsyncin_i                 : std_logic;
    signal   gt11_txsyncmode_i               : std_logic;
    signal   gt11_txsyncout_i                : std_logic;
    signal   gt11_txsyncdone_i               : std_logic;

    signal   gt11_txoutclk_i                 : std_logic;
    signal   gt11_rxoutclk_i                 : std_logic;
    signal   gt11_rxoutclk_i2                : std_logic;
    signal   gt11_txoutclk_i2                : std_logic;
    signal   gt11_recclk_stable_i            : std_logic;
    signal   gt11_rx_cdrlocked               : std_logic;
    signal   gt11_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt11_rxphaligndone_i            : std_logic;
    signal   gt11_rxdlysreset_i              : std_logic;
    signal   gt11_rxdlysresetdone_i          : std_logic;
    signal   gt11_rxphdlyreset_i             : std_logic;
    signal   gt11_rxphalignen_i              : std_logic;
    signal   gt11_rxdlyen_i                  : std_logic;
    signal   gt11_rxphalign_i                : std_logic;
    signal   gt11_run_rx_phalignment_i       : std_logic;
    signal   gt11_rst_rx_phalignment_i       : std_logic;
    signal   gt11_rx_phalignment_done_i      : std_logic;
    signal   gt11_rxsyncallin_i              : std_logic;
    signal   gt11_rxsyncin_i                 : std_logic;
    signal   gt11_rxsyncmode_i               : std_logic;
    signal   gt11_rxsyncout_i                : std_logic;
    signal   gt11_rxsyncdone_i               : std_logic;
    signal   gt12_txphaligndone_i            : std_logic;
    signal   gt12_txdlysreset_i              : std_logic;
    signal   gt12_txdlysresetdone_i          : std_logic;
    signal   gt12_txphdlyreset_i             : std_logic;
    signal   gt12_txphalignen_i              : std_logic;
    signal   gt12_txdlyen_i                  : std_logic;
    signal   gt12_txphalign_i                : std_logic;
    signal   gt12_txphinit_i                 : std_logic;
    signal   gt12_txphinitdone_i             : std_logic;
    signal   gt12_run_tx_phalignment_i       : std_logic;
    signal   gt12_rst_tx_phalignment_i       : std_logic;
    signal   gt12_tx_phalignment_done_i      : std_logic;
    signal   gt12_txsyncallin_i              : std_logic;
    signal   gt12_txsyncin_i                 : std_logic;
    signal   gt12_txsyncmode_i               : std_logic;
    signal   gt12_txsyncout_i                : std_logic;
    signal   gt12_txsyncdone_i               : std_logic;

    signal   gt12_txoutclk_i                 : std_logic;
    signal   gt12_rxoutclk_i                 : std_logic;
    signal   gt12_rxoutclk_i2                : std_logic;
    signal   gt12_txoutclk_i2                : std_logic;
    signal   gt12_recclk_stable_i            : std_logic;
    signal   gt12_rx_cdrlocked               : std_logic;
    signal   gt12_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt12_rxphaligndone_i            : std_logic;
    signal   gt12_rxdlysreset_i              : std_logic;
    signal   gt12_rxdlysresetdone_i          : std_logic;
    signal   gt12_rxphdlyreset_i             : std_logic;
    signal   gt12_rxphalignen_i              : std_logic;
    signal   gt12_rxdlyen_i                  : std_logic;
    signal   gt12_rxphalign_i                : std_logic;
    signal   gt12_run_rx_phalignment_i       : std_logic;
    signal   gt12_rst_rx_phalignment_i       : std_logic;
    signal   gt12_rx_phalignment_done_i      : std_logic;
    signal   gt12_rxsyncallin_i              : std_logic;
    signal   gt12_rxsyncin_i                 : std_logic;
    signal   gt12_rxsyncmode_i               : std_logic;
    signal   gt12_rxsyncout_i                : std_logic;
    signal   gt12_rxsyncdone_i               : std_logic;
    signal   gt13_txphaligndone_i            : std_logic;
    signal   gt13_txdlysreset_i              : std_logic;
    signal   gt13_txdlysresetdone_i          : std_logic;
    signal   gt13_txphdlyreset_i             : std_logic;
    signal   gt13_txphalignen_i              : std_logic;
    signal   gt13_txdlyen_i                  : std_logic;
    signal   gt13_txphalign_i                : std_logic;
    signal   gt13_txphinit_i                 : std_logic;
    signal   gt13_txphinitdone_i             : std_logic;
    signal   gt13_run_tx_phalignment_i       : std_logic;
    signal   gt13_rst_tx_phalignment_i       : std_logic;
    signal   gt13_tx_phalignment_done_i      : std_logic;
    signal   gt13_txsyncallin_i              : std_logic;
    signal   gt13_txsyncin_i                 : std_logic;
    signal   gt13_txsyncmode_i               : std_logic;
    signal   gt13_txsyncout_i                : std_logic;
    signal   gt13_txsyncdone_i               : std_logic;

    signal   gt13_txoutclk_i                 : std_logic;
    signal   gt13_rxoutclk_i                 : std_logic;
    signal   gt13_rxoutclk_i2                : std_logic;
    signal   gt13_txoutclk_i2                : std_logic;
    signal   gt13_recclk_stable_i            : std_logic;
    signal   gt13_rx_cdrlocked               : std_logic;
    signal   gt13_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt13_rxphaligndone_i            : std_logic;
    signal   gt13_rxdlysreset_i              : std_logic;
    signal   gt13_rxdlysresetdone_i          : std_logic;
    signal   gt13_rxphdlyreset_i             : std_logic;
    signal   gt13_rxphalignen_i              : std_logic;
    signal   gt13_rxdlyen_i                  : std_logic;
    signal   gt13_rxphalign_i                : std_logic;
    signal   gt13_run_rx_phalignment_i       : std_logic;
    signal   gt13_rst_rx_phalignment_i       : std_logic;
    signal   gt13_rx_phalignment_done_i      : std_logic;
    signal   gt13_rxsyncallin_i              : std_logic;
    signal   gt13_rxsyncin_i                 : std_logic;
    signal   gt13_rxsyncmode_i               : std_logic;
    signal   gt13_rxsyncout_i                : std_logic;
    signal   gt13_rxsyncdone_i               : std_logic;
    signal   gt14_txphaligndone_i            : std_logic;
    signal   gt14_txdlysreset_i              : std_logic;
    signal   gt14_txdlysresetdone_i          : std_logic;
    signal   gt14_txphdlyreset_i             : std_logic;
    signal   gt14_txphalignen_i              : std_logic;
    signal   gt14_txdlyen_i                  : std_logic;
    signal   gt14_txphalign_i                : std_logic;
    signal   gt14_txphinit_i                 : std_logic;
    signal   gt14_txphinitdone_i             : std_logic;
    signal   gt14_run_tx_phalignment_i       : std_logic;
    signal   gt14_rst_tx_phalignment_i       : std_logic;
    signal   gt14_tx_phalignment_done_i      : std_logic;
    signal   gt14_txsyncallin_i              : std_logic;
    signal   gt14_txsyncin_i                 : std_logic;
    signal   gt14_txsyncmode_i               : std_logic;
    signal   gt14_txsyncout_i                : std_logic;
    signal   gt14_txsyncdone_i               : std_logic;

    signal   gt14_txoutclk_i                 : std_logic;
    signal   gt14_rxoutclk_i                 : std_logic;
    signal   gt14_rxoutclk_i2                : std_logic;
    signal   gt14_txoutclk_i2                : std_logic;
    signal   gt14_recclk_stable_i            : std_logic;
    signal   gt14_rx_cdrlocked               : std_logic;
    signal   gt14_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt14_rxphaligndone_i            : std_logic;
    signal   gt14_rxdlysreset_i              : std_logic;
    signal   gt14_rxdlysresetdone_i          : std_logic;
    signal   gt14_rxphdlyreset_i             : std_logic;
    signal   gt14_rxphalignen_i              : std_logic;
    signal   gt14_rxdlyen_i                  : std_logic;
    signal   gt14_rxphalign_i                : std_logic;
    signal   gt14_run_rx_phalignment_i       : std_logic;
    signal   gt14_rst_rx_phalignment_i       : std_logic;
    signal   gt14_rx_phalignment_done_i      : std_logic;
    signal   gt14_rxsyncallin_i              : std_logic;
    signal   gt14_rxsyncin_i                 : std_logic;
    signal   gt14_rxsyncmode_i               : std_logic;
    signal   gt14_rxsyncout_i                : std_logic;
    signal   gt14_rxsyncdone_i               : std_logic;
    signal   gt15_txphaligndone_i            : std_logic;
    signal   gt15_txdlysreset_i              : std_logic;
    signal   gt15_txdlysresetdone_i          : std_logic;
    signal   gt15_txphdlyreset_i             : std_logic;
    signal   gt15_txphalignen_i              : std_logic;
    signal   gt15_txdlyen_i                  : std_logic;
    signal   gt15_txphalign_i                : std_logic;
    signal   gt15_txphinit_i                 : std_logic;
    signal   gt15_txphinitdone_i             : std_logic;
    signal   gt15_run_tx_phalignment_i       : std_logic;
    signal   gt15_rst_tx_phalignment_i       : std_logic;
    signal   gt15_tx_phalignment_done_i      : std_logic;
    signal   gt15_txsyncallin_i              : std_logic;
    signal   gt15_txsyncin_i                 : std_logic;
    signal   gt15_txsyncmode_i               : std_logic;
    signal   gt15_txsyncout_i                : std_logic;
    signal   gt15_txsyncdone_i               : std_logic;

    signal   gt15_txoutclk_i                 : std_logic;
    signal   gt15_rxoutclk_i                 : std_logic;
    signal   gt15_rxoutclk_i2                : std_logic;
    signal   gt15_txoutclk_i2                : std_logic;
    signal   gt15_recclk_stable_i            : std_logic;
    signal   gt15_rx_cdrlocked               : std_logic;
    signal   gt15_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt15_rxphaligndone_i            : std_logic;
    signal   gt15_rxdlysreset_i              : std_logic;
    signal   gt15_rxdlysresetdone_i          : std_logic;
    signal   gt15_rxphdlyreset_i             : std_logic;
    signal   gt15_rxphalignen_i              : std_logic;
    signal   gt15_rxdlyen_i                  : std_logic;
    signal   gt15_rxphalign_i                : std_logic;
    signal   gt15_run_rx_phalignment_i       : std_logic;
    signal   gt15_rst_rx_phalignment_i       : std_logic;
    signal   gt15_rx_phalignment_done_i      : std_logic;
    signal   gt15_rxsyncallin_i              : std_logic;
    signal   gt15_rxsyncin_i                 : std_logic;
    signal   gt15_rxsyncmode_i               : std_logic;
    signal   gt15_rxsyncout_i                : std_logic;
    signal   gt15_rxsyncdone_i               : std_logic;
    signal   gt16_txphaligndone_i            : std_logic;
    signal   gt16_txdlysreset_i              : std_logic;
    signal   gt16_txdlysresetdone_i          : std_logic;
    signal   gt16_txphdlyreset_i             : std_logic;
    signal   gt16_txphalignen_i              : std_logic;
    signal   gt16_txdlyen_i                  : std_logic;
    signal   gt16_txphalign_i                : std_logic;
    signal   gt16_txphinit_i                 : std_logic;
    signal   gt16_txphinitdone_i             : std_logic;
    signal   gt16_run_tx_phalignment_i       : std_logic;
    signal   gt16_rst_tx_phalignment_i       : std_logic;
    signal   gt16_tx_phalignment_done_i      : std_logic;
    signal   gt16_txsyncallin_i              : std_logic;
    signal   gt16_txsyncin_i                 : std_logic;
    signal   gt16_txsyncmode_i               : std_logic;
    signal   gt16_txsyncout_i                : std_logic;
    signal   gt16_txsyncdone_i               : std_logic;

    signal   gt16_txoutclk_i                 : std_logic;
    signal   gt16_rxoutclk_i                 : std_logic;
    signal   gt16_rxoutclk_i2                : std_logic;
    signal   gt16_txoutclk_i2                : std_logic;
    signal   gt16_recclk_stable_i            : std_logic;
    signal   gt16_rx_cdrlocked               : std_logic;
    signal   gt16_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt16_rxphaligndone_i            : std_logic;
    signal   gt16_rxdlysreset_i              : std_logic;
    signal   gt16_rxdlysresetdone_i          : std_logic;
    signal   gt16_rxphdlyreset_i             : std_logic;
    signal   gt16_rxphalignen_i              : std_logic;
    signal   gt16_rxdlyen_i                  : std_logic;
    signal   gt16_rxphalign_i                : std_logic;
    signal   gt16_run_rx_phalignment_i       : std_logic;
    signal   gt16_rst_rx_phalignment_i       : std_logic;
    signal   gt16_rx_phalignment_done_i      : std_logic;
    signal   gt16_rxsyncallin_i              : std_logic;
    signal   gt16_rxsyncin_i                 : std_logic;
    signal   gt16_rxsyncmode_i               : std_logic;
    signal   gt16_rxsyncout_i                : std_logic;
    signal   gt16_rxsyncdone_i               : std_logic;
    signal   gt17_txphaligndone_i            : std_logic;
    signal   gt17_txdlysreset_i              : std_logic;
    signal   gt17_txdlysresetdone_i          : std_logic;
    signal   gt17_txphdlyreset_i             : std_logic;
    signal   gt17_txphalignen_i              : std_logic;
    signal   gt17_txdlyen_i                  : std_logic;
    signal   gt17_txphalign_i                : std_logic;
    signal   gt17_txphinit_i                 : std_logic;
    signal   gt17_txphinitdone_i             : std_logic;
    signal   gt17_run_tx_phalignment_i       : std_logic;
    signal   gt17_rst_tx_phalignment_i       : std_logic;
    signal   gt17_tx_phalignment_done_i      : std_logic;
    signal   gt17_txsyncallin_i              : std_logic;
    signal   gt17_txsyncin_i                 : std_logic;
    signal   gt17_txsyncmode_i               : std_logic;
    signal   gt17_txsyncout_i                : std_logic;
    signal   gt17_txsyncdone_i               : std_logic;

    signal   gt17_txoutclk_i                 : std_logic;
    signal   gt17_rxoutclk_i                 : std_logic;
    signal   gt17_rxoutclk_i2                : std_logic;
    signal   gt17_txoutclk_i2                : std_logic;
    signal   gt17_recclk_stable_i            : std_logic;
    signal   gt17_rx_cdrlocked               : std_logic;
    signal   gt17_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt17_rxphaligndone_i            : std_logic;
    signal   gt17_rxdlysreset_i              : std_logic;
    signal   gt17_rxdlysresetdone_i          : std_logic;
    signal   gt17_rxphdlyreset_i             : std_logic;
    signal   gt17_rxphalignen_i              : std_logic;
    signal   gt17_rxdlyen_i                  : std_logic;
    signal   gt17_rxphalign_i                : std_logic;
    signal   gt17_run_rx_phalignment_i       : std_logic;
    signal   gt17_rst_rx_phalignment_i       : std_logic;
    signal   gt17_rx_phalignment_done_i      : std_logic;
    signal   gt17_rxsyncallin_i              : std_logic;
    signal   gt17_rxsyncin_i                 : std_logic;
    signal   gt17_rxsyncmode_i               : std_logic;
    signal   gt17_rxsyncout_i                : std_logic;
    signal   gt17_rxsyncdone_i               : std_logic;
    signal   gt18_txphaligndone_i            : std_logic;
    signal   gt18_txdlysreset_i              : std_logic;
    signal   gt18_txdlysresetdone_i          : std_logic;
    signal   gt18_txphdlyreset_i             : std_logic;
    signal   gt18_txphalignen_i              : std_logic;
    signal   gt18_txdlyen_i                  : std_logic;
    signal   gt18_txphalign_i                : std_logic;
    signal   gt18_txphinit_i                 : std_logic;
    signal   gt18_txphinitdone_i             : std_logic;
    signal   gt18_run_tx_phalignment_i       : std_logic;
    signal   gt18_rst_tx_phalignment_i       : std_logic;
    signal   gt18_tx_phalignment_done_i      : std_logic;
    signal   gt18_txsyncallin_i              : std_logic;
    signal   gt18_txsyncin_i                 : std_logic;
    signal   gt18_txsyncmode_i               : std_logic;
    signal   gt18_txsyncout_i                : std_logic;
    signal   gt18_txsyncdone_i               : std_logic;

    signal   gt18_txoutclk_i                 : std_logic;
    signal   gt18_rxoutclk_i                 : std_logic;
    signal   gt18_rxoutclk_i2                : std_logic;
    signal   gt18_txoutclk_i2                : std_logic;
    signal   gt18_recclk_stable_i            : std_logic;
    signal   gt18_rx_cdrlocked               : std_logic;
    signal   gt18_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt18_rxphaligndone_i            : std_logic;
    signal   gt18_rxdlysreset_i              : std_logic;
    signal   gt18_rxdlysresetdone_i          : std_logic;
    signal   gt18_rxphdlyreset_i             : std_logic;
    signal   gt18_rxphalignen_i              : std_logic;
    signal   gt18_rxdlyen_i                  : std_logic;
    signal   gt18_rxphalign_i                : std_logic;
    signal   gt18_run_rx_phalignment_i       : std_logic;
    signal   gt18_rst_rx_phalignment_i       : std_logic;
    signal   gt18_rx_phalignment_done_i      : std_logic;
    signal   gt18_rxsyncallin_i              : std_logic;
    signal   gt18_rxsyncin_i                 : std_logic;
    signal   gt18_rxsyncmode_i               : std_logic;
    signal   gt18_rxsyncout_i                : std_logic;
    signal   gt18_rxsyncdone_i               : std_logic;
    signal   gt19_txphaligndone_i            : std_logic;
    signal   gt19_txdlysreset_i              : std_logic;
    signal   gt19_txdlysresetdone_i          : std_logic;
    signal   gt19_txphdlyreset_i             : std_logic;
    signal   gt19_txphalignen_i              : std_logic;
    signal   gt19_txdlyen_i                  : std_logic;
    signal   gt19_txphalign_i                : std_logic;
    signal   gt19_txphinit_i                 : std_logic;
    signal   gt19_txphinitdone_i             : std_logic;
    signal   gt19_run_tx_phalignment_i       : std_logic;
    signal   gt19_rst_tx_phalignment_i       : std_logic;
    signal   gt19_tx_phalignment_done_i      : std_logic;
    signal   gt19_txsyncallin_i              : std_logic;
    signal   gt19_txsyncin_i                 : std_logic;
    signal   gt19_txsyncmode_i               : std_logic;
    signal   gt19_txsyncout_i                : std_logic;
    signal   gt19_txsyncdone_i               : std_logic;

    signal   gt19_txoutclk_i                 : std_logic;
    signal   gt19_rxoutclk_i                 : std_logic;
    signal   gt19_rxoutclk_i2                : std_logic;
    signal   gt19_txoutclk_i2                : std_logic;
    signal   gt19_recclk_stable_i            : std_logic;
    signal   gt19_rx_cdrlocked               : std_logic;
    signal   gt19_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt19_rxphaligndone_i            : std_logic;
    signal   gt19_rxdlysreset_i              : std_logic;
    signal   gt19_rxdlysresetdone_i          : std_logic;
    signal   gt19_rxphdlyreset_i             : std_logic;
    signal   gt19_rxphalignen_i              : std_logic;
    signal   gt19_rxdlyen_i                  : std_logic;
    signal   gt19_rxphalign_i                : std_logic;
    signal   gt19_run_rx_phalignment_i       : std_logic;
    signal   gt19_rst_rx_phalignment_i       : std_logic;
    signal   gt19_rx_phalignment_done_i      : std_logic;
    signal   gt19_rxsyncallin_i              : std_logic;
    signal   gt19_rxsyncin_i                 : std_logic;
    signal   gt19_rxsyncmode_i               : std_logic;
    signal   gt19_rxsyncout_i                : std_logic;
    signal   gt19_rxsyncdone_i               : std_logic;
    signal   gt20_txphaligndone_i            : std_logic;
    signal   gt20_txdlysreset_i              : std_logic;
    signal   gt20_txdlysresetdone_i          : std_logic;
    signal   gt20_txphdlyreset_i             : std_logic;
    signal   gt20_txphalignen_i              : std_logic;
    signal   gt20_txdlyen_i                  : std_logic;
    signal   gt20_txphalign_i                : std_logic;
    signal   gt20_txphinit_i                 : std_logic;
    signal   gt20_txphinitdone_i             : std_logic;
    signal   gt20_run_tx_phalignment_i       : std_logic;
    signal   gt20_rst_tx_phalignment_i       : std_logic;
    signal   gt20_tx_phalignment_done_i      : std_logic;
    signal   gt20_txsyncallin_i              : std_logic;
    signal   gt20_txsyncin_i                 : std_logic;
    signal   gt20_txsyncmode_i               : std_logic;
    signal   gt20_txsyncout_i                : std_logic;
    signal   gt20_txsyncdone_i               : std_logic;

    signal   gt20_txoutclk_i                 : std_logic;
    signal   gt20_rxoutclk_i                 : std_logic;
    signal   gt20_rxoutclk_i2                : std_logic;
    signal   gt20_txoutclk_i2                : std_logic;
    signal   gt20_recclk_stable_i            : std_logic;
    signal   gt20_rx_cdrlocked               : std_logic;
    signal   gt20_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt20_rxphaligndone_i            : std_logic;
    signal   gt20_rxdlysreset_i              : std_logic;
    signal   gt20_rxdlysresetdone_i          : std_logic;
    signal   gt20_rxphdlyreset_i             : std_logic;
    signal   gt20_rxphalignen_i              : std_logic;
    signal   gt20_rxdlyen_i                  : std_logic;
    signal   gt20_rxphalign_i                : std_logic;
    signal   gt20_run_rx_phalignment_i       : std_logic;
    signal   gt20_rst_rx_phalignment_i       : std_logic;
    signal   gt20_rx_phalignment_done_i      : std_logic;
    signal   gt20_rxsyncallin_i              : std_logic;
    signal   gt20_rxsyncin_i                 : std_logic;
    signal   gt20_rxsyncmode_i               : std_logic;
    signal   gt20_rxsyncout_i                : std_logic;
    signal   gt20_rxsyncdone_i               : std_logic;
    signal   gt21_txphaligndone_i            : std_logic;
    signal   gt21_txdlysreset_i              : std_logic;
    signal   gt21_txdlysresetdone_i          : std_logic;
    signal   gt21_txphdlyreset_i             : std_logic;
    signal   gt21_txphalignen_i              : std_logic;
    signal   gt21_txdlyen_i                  : std_logic;
    signal   gt21_txphalign_i                : std_logic;
    signal   gt21_txphinit_i                 : std_logic;
    signal   gt21_txphinitdone_i             : std_logic;
    signal   gt21_run_tx_phalignment_i       : std_logic;
    signal   gt21_rst_tx_phalignment_i       : std_logic;
    signal   gt21_tx_phalignment_done_i      : std_logic;
    signal   gt21_txsyncallin_i              : std_logic;
    signal   gt21_txsyncin_i                 : std_logic;
    signal   gt21_txsyncmode_i               : std_logic;
    signal   gt21_txsyncout_i                : std_logic;
    signal   gt21_txsyncdone_i               : std_logic;

    signal   gt21_txoutclk_i                 : std_logic;
    signal   gt21_rxoutclk_i                 : std_logic;
    signal   gt21_rxoutclk_i2                : std_logic;
    signal   gt21_txoutclk_i2                : std_logic;
    signal   gt21_recclk_stable_i            : std_logic;
    signal   gt21_rx_cdrlocked               : std_logic;
    signal   gt21_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt21_rxphaligndone_i            : std_logic;
    signal   gt21_rxdlysreset_i              : std_logic;
    signal   gt21_rxdlysresetdone_i          : std_logic;
    signal   gt21_rxphdlyreset_i             : std_logic;
    signal   gt21_rxphalignen_i              : std_logic;
    signal   gt21_rxdlyen_i                  : std_logic;
    signal   gt21_rxphalign_i                : std_logic;
    signal   gt21_run_rx_phalignment_i       : std_logic;
    signal   gt21_rst_rx_phalignment_i       : std_logic;
    signal   gt21_rx_phalignment_done_i      : std_logic;
    signal   gt21_rxsyncallin_i              : std_logic;
    signal   gt21_rxsyncin_i                 : std_logic;
    signal   gt21_rxsyncmode_i               : std_logic;
    signal   gt21_rxsyncout_i                : std_logic;
    signal   gt21_rxsyncdone_i               : std_logic;
    signal   gt22_txphaligndone_i            : std_logic;
    signal   gt22_txdlysreset_i              : std_logic;
    signal   gt22_txdlysresetdone_i          : std_logic;
    signal   gt22_txphdlyreset_i             : std_logic;
    signal   gt22_txphalignen_i              : std_logic;
    signal   gt22_txdlyen_i                  : std_logic;
    signal   gt22_txphalign_i                : std_logic;
    signal   gt22_txphinit_i                 : std_logic;
    signal   gt22_txphinitdone_i             : std_logic;
    signal   gt22_run_tx_phalignment_i       : std_logic;
    signal   gt22_rst_tx_phalignment_i       : std_logic;
    signal   gt22_tx_phalignment_done_i      : std_logic;
    signal   gt22_txsyncallin_i              : std_logic;
    signal   gt22_txsyncin_i                 : std_logic;
    signal   gt22_txsyncmode_i               : std_logic;
    signal   gt22_txsyncout_i                : std_logic;
    signal   gt22_txsyncdone_i               : std_logic;

    signal   gt22_txoutclk_i                 : std_logic;
    signal   gt22_rxoutclk_i                 : std_logic;
    signal   gt22_rxoutclk_i2                : std_logic;
    signal   gt22_txoutclk_i2                : std_logic;
    signal   gt22_recclk_stable_i            : std_logic;
    signal   gt22_rx_cdrlocked               : std_logic;
    signal   gt22_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt22_rxphaligndone_i            : std_logic;
    signal   gt22_rxdlysreset_i              : std_logic;
    signal   gt22_rxdlysresetdone_i          : std_logic;
    signal   gt22_rxphdlyreset_i             : std_logic;
    signal   gt22_rxphalignen_i              : std_logic;
    signal   gt22_rxdlyen_i                  : std_logic;
    signal   gt22_rxphalign_i                : std_logic;
    signal   gt22_run_rx_phalignment_i       : std_logic;
    signal   gt22_rst_rx_phalignment_i       : std_logic;
    signal   gt22_rx_phalignment_done_i      : std_logic;
    signal   gt22_rxsyncallin_i              : std_logic;
    signal   gt22_rxsyncin_i                 : std_logic;
    signal   gt22_rxsyncmode_i               : std_logic;
    signal   gt22_rxsyncout_i                : std_logic;
    signal   gt22_rxsyncdone_i               : std_logic;
    signal   gt23_txphaligndone_i            : std_logic;
    signal   gt23_txdlysreset_i              : std_logic;
    signal   gt23_txdlysresetdone_i          : std_logic;
    signal   gt23_txphdlyreset_i             : std_logic;
    signal   gt23_txphalignen_i              : std_logic;
    signal   gt23_txdlyen_i                  : std_logic;
    signal   gt23_txphalign_i                : std_logic;
    signal   gt23_txphinit_i                 : std_logic;
    signal   gt23_txphinitdone_i             : std_logic;
    signal   gt23_run_tx_phalignment_i       : std_logic;
    signal   gt23_rst_tx_phalignment_i       : std_logic;
    signal   gt23_tx_phalignment_done_i      : std_logic;
    signal   gt23_txsyncallin_i              : std_logic;
    signal   gt23_txsyncin_i                 : std_logic;
    signal   gt23_txsyncmode_i               : std_logic;
    signal   gt23_txsyncout_i                : std_logic;
    signal   gt23_txsyncdone_i               : std_logic;

    signal   gt23_txoutclk_i                 : std_logic;
    signal   gt23_rxoutclk_i                 : std_logic;
    signal   gt23_rxoutclk_i2                : std_logic;
    signal   gt23_txoutclk_i2                : std_logic;
    signal   gt23_recclk_stable_i            : std_logic;
    signal   gt23_rx_cdrlocked               : std_logic;
    signal   gt23_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt23_rxphaligndone_i            : std_logic;
    signal   gt23_rxdlysreset_i              : std_logic;
    signal   gt23_rxdlysresetdone_i          : std_logic;
    signal   gt23_rxphdlyreset_i             : std_logic;
    signal   gt23_rxphalignen_i              : std_logic;
    signal   gt23_rxdlyen_i                  : std_logic;
    signal   gt23_rxphalign_i                : std_logic;
    signal   gt23_run_rx_phalignment_i       : std_logic;
    signal   gt23_rst_rx_phalignment_i       : std_logic;
    signal   gt23_rx_phalignment_done_i      : std_logic;
    signal   gt23_rxsyncallin_i              : std_logic;
    signal   gt23_rxsyncin_i                 : std_logic;
    signal   gt23_rxsyncmode_i               : std_logic;
    signal   gt23_rxsyncout_i                : std_logic;
    signal   gt23_rxsyncdone_i               : std_logic;
    signal   gt24_txphaligndone_i            : std_logic;
    signal   gt24_txdlysreset_i              : std_logic;
    signal   gt24_txdlysresetdone_i          : std_logic;
    signal   gt24_txphdlyreset_i             : std_logic;
    signal   gt24_txphalignen_i              : std_logic;
    signal   gt24_txdlyen_i                  : std_logic;
    signal   gt24_txphalign_i                : std_logic;
    signal   gt24_txphinit_i                 : std_logic;
    signal   gt24_txphinitdone_i             : std_logic;
    signal   gt24_run_tx_phalignment_i       : std_logic;
    signal   gt24_rst_tx_phalignment_i       : std_logic;
    signal   gt24_tx_phalignment_done_i      : std_logic;
    signal   gt24_txsyncallin_i              : std_logic;
    signal   gt24_txsyncin_i                 : std_logic;
    signal   gt24_txsyncmode_i               : std_logic;
    signal   gt24_txsyncout_i                : std_logic;
    signal   gt24_txsyncdone_i               : std_logic;

    signal   gt24_txoutclk_i                 : std_logic;
    signal   gt24_rxoutclk_i                 : std_logic;
    signal   gt24_rxoutclk_i2                : std_logic;
    signal   gt24_txoutclk_i2                : std_logic;
    signal   gt24_recclk_stable_i            : std_logic;
    signal   gt24_rx_cdrlocked               : std_logic;
    signal   gt24_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt24_rxphaligndone_i            : std_logic;
    signal   gt24_rxdlysreset_i              : std_logic;
    signal   gt24_rxdlysresetdone_i          : std_logic;
    signal   gt24_rxphdlyreset_i             : std_logic;
    signal   gt24_rxphalignen_i              : std_logic;
    signal   gt24_rxdlyen_i                  : std_logic;
    signal   gt24_rxphalign_i                : std_logic;
    signal   gt24_run_rx_phalignment_i       : std_logic;
    signal   gt24_rst_rx_phalignment_i       : std_logic;
    signal   gt24_rx_phalignment_done_i      : std_logic;
    signal   gt24_rxsyncallin_i              : std_logic;
    signal   gt24_rxsyncin_i                 : std_logic;
    signal   gt24_rxsyncmode_i               : std_logic;
    signal   gt24_rxsyncout_i                : std_logic;
    signal   gt24_rxsyncdone_i               : std_logic;
    signal   gt25_txphaligndone_i            : std_logic;
    signal   gt25_txdlysreset_i              : std_logic;
    signal   gt25_txdlysresetdone_i          : std_logic;
    signal   gt25_txphdlyreset_i             : std_logic;
    signal   gt25_txphalignen_i              : std_logic;
    signal   gt25_txdlyen_i                  : std_logic;
    signal   gt25_txphalign_i                : std_logic;
    signal   gt25_txphinit_i                 : std_logic;
    signal   gt25_txphinitdone_i             : std_logic;
    signal   gt25_run_tx_phalignment_i       : std_logic;
    signal   gt25_rst_tx_phalignment_i       : std_logic;
    signal   gt25_tx_phalignment_done_i      : std_logic;
    signal   gt25_txsyncallin_i              : std_logic;
    signal   gt25_txsyncin_i                 : std_logic;
    signal   gt25_txsyncmode_i               : std_logic;
    signal   gt25_txsyncout_i                : std_logic;
    signal   gt25_txsyncdone_i               : std_logic;

    signal   gt25_txoutclk_i                 : std_logic;
    signal   gt25_rxoutclk_i                 : std_logic;
    signal   gt25_rxoutclk_i2                : std_logic;
    signal   gt25_txoutclk_i2                : std_logic;
    signal   gt25_recclk_stable_i            : std_logic;
    signal   gt25_rx_cdrlocked               : std_logic;
    signal   gt25_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt25_rxphaligndone_i            : std_logic;
    signal   gt25_rxdlysreset_i              : std_logic;
    signal   gt25_rxdlysresetdone_i          : std_logic;
    signal   gt25_rxphdlyreset_i             : std_logic;
    signal   gt25_rxphalignen_i              : std_logic;
    signal   gt25_rxdlyen_i                  : std_logic;
    signal   gt25_rxphalign_i                : std_logic;
    signal   gt25_run_rx_phalignment_i       : std_logic;
    signal   gt25_rst_rx_phalignment_i       : std_logic;
    signal   gt25_rx_phalignment_done_i      : std_logic;
    signal   gt25_rxsyncallin_i              : std_logic;
    signal   gt25_rxsyncin_i                 : std_logic;
    signal   gt25_rxsyncmode_i               : std_logic;
    signal   gt25_rxsyncout_i                : std_logic;
    signal   gt25_rxsyncdone_i               : std_logic;
    signal   gt26_txphaligndone_i            : std_logic;
    signal   gt26_txdlysreset_i              : std_logic;
    signal   gt26_txdlysresetdone_i          : std_logic;
    signal   gt26_txphdlyreset_i             : std_logic;
    signal   gt26_txphalignen_i              : std_logic;
    signal   gt26_txdlyen_i                  : std_logic;
    signal   gt26_txphalign_i                : std_logic;
    signal   gt26_txphinit_i                 : std_logic;
    signal   gt26_txphinitdone_i             : std_logic;
    signal   gt26_run_tx_phalignment_i       : std_logic;
    signal   gt26_rst_tx_phalignment_i       : std_logic;
    signal   gt26_tx_phalignment_done_i      : std_logic;
    signal   gt26_txsyncallin_i              : std_logic;
    signal   gt26_txsyncin_i                 : std_logic;
    signal   gt26_txsyncmode_i               : std_logic;
    signal   gt26_txsyncout_i                : std_logic;
    signal   gt26_txsyncdone_i               : std_logic;

    signal   gt26_txoutclk_i                 : std_logic;
    signal   gt26_rxoutclk_i                 : std_logic;
    signal   gt26_rxoutclk_i2                : std_logic;
    signal   gt26_txoutclk_i2                : std_logic;
    signal   gt26_recclk_stable_i            : std_logic;
    signal   gt26_rx_cdrlocked               : std_logic;
    signal   gt26_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt26_rxphaligndone_i            : std_logic;
    signal   gt26_rxdlysreset_i              : std_logic;
    signal   gt26_rxdlysresetdone_i          : std_logic;
    signal   gt26_rxphdlyreset_i             : std_logic;
    signal   gt26_rxphalignen_i              : std_logic;
    signal   gt26_rxdlyen_i                  : std_logic;
    signal   gt26_rxphalign_i                : std_logic;
    signal   gt26_run_rx_phalignment_i       : std_logic;
    signal   gt26_rst_rx_phalignment_i       : std_logic;
    signal   gt26_rx_phalignment_done_i      : std_logic;
    signal   gt26_rxsyncallin_i              : std_logic;
    signal   gt26_rxsyncin_i                 : std_logic;
    signal   gt26_rxsyncmode_i               : std_logic;
    signal   gt26_rxsyncout_i                : std_logic;
    signal   gt26_rxsyncdone_i               : std_logic;
    signal   gt27_txphaligndone_i            : std_logic;
    signal   gt27_txdlysreset_i              : std_logic;
    signal   gt27_txdlysresetdone_i          : std_logic;
    signal   gt27_txphdlyreset_i             : std_logic;
    signal   gt27_txphalignen_i              : std_logic;
    signal   gt27_txdlyen_i                  : std_logic;
    signal   gt27_txphalign_i                : std_logic;
    signal   gt27_txphinit_i                 : std_logic;
    signal   gt27_txphinitdone_i             : std_logic;
    signal   gt27_run_tx_phalignment_i       : std_logic;
    signal   gt27_rst_tx_phalignment_i       : std_logic;
    signal   gt27_tx_phalignment_done_i      : std_logic;
    signal   gt27_txsyncallin_i              : std_logic;
    signal   gt27_txsyncin_i                 : std_logic;
    signal   gt27_txsyncmode_i               : std_logic;
    signal   gt27_txsyncout_i                : std_logic;
    signal   gt27_txsyncdone_i               : std_logic;

    signal   gt27_txoutclk_i                 : std_logic;
    signal   gt27_rxoutclk_i                 : std_logic;
    signal   gt27_rxoutclk_i2                : std_logic;
    signal   gt27_txoutclk_i2                : std_logic;
    signal   gt27_recclk_stable_i            : std_logic;
    signal   gt27_rx_cdrlocked               : std_logic;
    signal   gt27_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt27_rxphaligndone_i            : std_logic;
    signal   gt27_rxdlysreset_i              : std_logic;
    signal   gt27_rxdlysresetdone_i          : std_logic;
    signal   gt27_rxphdlyreset_i             : std_logic;
    signal   gt27_rxphalignen_i              : std_logic;
    signal   gt27_rxdlyen_i                  : std_logic;
    signal   gt27_rxphalign_i                : std_logic;
    signal   gt27_run_rx_phalignment_i       : std_logic;
    signal   gt27_rst_rx_phalignment_i       : std_logic;
    signal   gt27_rx_phalignment_done_i      : std_logic;
    signal   gt27_rxsyncallin_i              : std_logic;
    signal   gt27_rxsyncin_i                 : std_logic;
    signal   gt27_rxsyncmode_i               : std_logic;
    signal   gt27_rxsyncout_i                : std_logic;
    signal   gt27_rxsyncdone_i               : std_logic;
    signal   gt28_txphaligndone_i            : std_logic;
    signal   gt28_txdlysreset_i              : std_logic;
    signal   gt28_txdlysresetdone_i          : std_logic;
    signal   gt28_txphdlyreset_i             : std_logic;
    signal   gt28_txphalignen_i              : std_logic;
    signal   gt28_txdlyen_i                  : std_logic;
    signal   gt28_txphalign_i                : std_logic;
    signal   gt28_txphinit_i                 : std_logic;
    signal   gt28_txphinitdone_i             : std_logic;
    signal   gt28_run_tx_phalignment_i       : std_logic;
    signal   gt28_rst_tx_phalignment_i       : std_logic;
    signal   gt28_tx_phalignment_done_i      : std_logic;
    signal   gt28_txsyncallin_i              : std_logic;
    signal   gt28_txsyncin_i                 : std_logic;
    signal   gt28_txsyncmode_i               : std_logic;
    signal   gt28_txsyncout_i                : std_logic;
    signal   gt28_txsyncdone_i               : std_logic;

    signal   gt28_txoutclk_i                 : std_logic;
    signal   gt28_rxoutclk_i                 : std_logic;
    signal   gt28_rxoutclk_i2                : std_logic;
    signal   gt28_txoutclk_i2                : std_logic;
    signal   gt28_recclk_stable_i            : std_logic;
    signal   gt28_rx_cdrlocked               : std_logic;
    signal   gt28_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt28_rxphaligndone_i            : std_logic;
    signal   gt28_rxdlysreset_i              : std_logic;
    signal   gt28_rxdlysresetdone_i          : std_logic;
    signal   gt28_rxphdlyreset_i             : std_logic;
    signal   gt28_rxphalignen_i              : std_logic;
    signal   gt28_rxdlyen_i                  : std_logic;
    signal   gt28_rxphalign_i                : std_logic;
    signal   gt28_run_rx_phalignment_i       : std_logic;
    signal   gt28_rst_rx_phalignment_i       : std_logic;
    signal   gt28_rx_phalignment_done_i      : std_logic;
    signal   gt28_rxsyncallin_i              : std_logic;
    signal   gt28_rxsyncin_i                 : std_logic;
    signal   gt28_rxsyncmode_i               : std_logic;
    signal   gt28_rxsyncout_i                : std_logic;
    signal   gt28_rxsyncdone_i               : std_logic;
    signal   gt29_txphaligndone_i            : std_logic;
    signal   gt29_txdlysreset_i              : std_logic;
    signal   gt29_txdlysresetdone_i          : std_logic;
    signal   gt29_txphdlyreset_i             : std_logic;
    signal   gt29_txphalignen_i              : std_logic;
    signal   gt29_txdlyen_i                  : std_logic;
    signal   gt29_txphalign_i                : std_logic;
    signal   gt29_txphinit_i                 : std_logic;
    signal   gt29_txphinitdone_i             : std_logic;
    signal   gt29_run_tx_phalignment_i       : std_logic;
    signal   gt29_rst_tx_phalignment_i       : std_logic;
    signal   gt29_tx_phalignment_done_i      : std_logic;
    signal   gt29_txsyncallin_i              : std_logic;
    signal   gt29_txsyncin_i                 : std_logic;
    signal   gt29_txsyncmode_i               : std_logic;
    signal   gt29_txsyncout_i                : std_logic;
    signal   gt29_txsyncdone_i               : std_logic;

    signal   gt29_txoutclk_i                 : std_logic;
    signal   gt29_rxoutclk_i                 : std_logic;
    signal   gt29_rxoutclk_i2                : std_logic;
    signal   gt29_txoutclk_i2                : std_logic;
    signal   gt29_recclk_stable_i            : std_logic;
    signal   gt29_rx_cdrlocked               : std_logic;
    signal   gt29_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt29_rxphaligndone_i            : std_logic;
    signal   gt29_rxdlysreset_i              : std_logic;
    signal   gt29_rxdlysresetdone_i          : std_logic;
    signal   gt29_rxphdlyreset_i             : std_logic;
    signal   gt29_rxphalignen_i              : std_logic;
    signal   gt29_rxdlyen_i                  : std_logic;
    signal   gt29_rxphalign_i                : std_logic;
    signal   gt29_run_rx_phalignment_i       : std_logic;
    signal   gt29_rst_rx_phalignment_i       : std_logic;
    signal   gt29_rx_phalignment_done_i      : std_logic;
    signal   gt29_rxsyncallin_i              : std_logic;
    signal   gt29_rxsyncin_i                 : std_logic;
    signal   gt29_rxsyncmode_i               : std_logic;
    signal   gt29_rxsyncout_i                : std_logic;
    signal   gt29_rxsyncdone_i               : std_logic;
    signal   gt30_txphaligndone_i            : std_logic;
    signal   gt30_txdlysreset_i              : std_logic;
    signal   gt30_txdlysresetdone_i          : std_logic;
    signal   gt30_txphdlyreset_i             : std_logic;
    signal   gt30_txphalignen_i              : std_logic;
    signal   gt30_txdlyen_i                  : std_logic;
    signal   gt30_txphalign_i                : std_logic;
    signal   gt30_txphinit_i                 : std_logic;
    signal   gt30_txphinitdone_i             : std_logic;
    signal   gt30_run_tx_phalignment_i       : std_logic;
    signal   gt30_rst_tx_phalignment_i       : std_logic;
    signal   gt30_tx_phalignment_done_i      : std_logic;
    signal   gt30_txsyncallin_i              : std_logic;
    signal   gt30_txsyncin_i                 : std_logic;
    signal   gt30_txsyncmode_i               : std_logic;
    signal   gt30_txsyncout_i                : std_logic;
    signal   gt30_txsyncdone_i               : std_logic;

    signal   gt30_txoutclk_i                 : std_logic;
    signal   gt30_rxoutclk_i                 : std_logic;
    signal   gt30_rxoutclk_i2                : std_logic;
    signal   gt30_txoutclk_i2                : std_logic;
    signal   gt30_recclk_stable_i            : std_logic;
    signal   gt30_rx_cdrlocked               : std_logic;
    signal   gt30_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt30_rxphaligndone_i            : std_logic;
    signal   gt30_rxdlysreset_i              : std_logic;
    signal   gt30_rxdlysresetdone_i          : std_logic;
    signal   gt30_rxphdlyreset_i             : std_logic;
    signal   gt30_rxphalignen_i              : std_logic;
    signal   gt30_rxdlyen_i                  : std_logic;
    signal   gt30_rxphalign_i                : std_logic;
    signal   gt30_run_rx_phalignment_i       : std_logic;
    signal   gt30_rst_rx_phalignment_i       : std_logic;
    signal   gt30_rx_phalignment_done_i      : std_logic;
    signal   gt30_rxsyncallin_i              : std_logic;
    signal   gt30_rxsyncin_i                 : std_logic;
    signal   gt30_rxsyncmode_i               : std_logic;
    signal   gt30_rxsyncout_i                : std_logic;
    signal   gt30_rxsyncdone_i               : std_logic;
    signal   gt31_txphaligndone_i            : std_logic;
    signal   gt31_txdlysreset_i              : std_logic;
    signal   gt31_txdlysresetdone_i          : std_logic;
    signal   gt31_txphdlyreset_i             : std_logic;
    signal   gt31_txphalignen_i              : std_logic;
    signal   gt31_txdlyen_i                  : std_logic;
    signal   gt31_txphalign_i                : std_logic;
    signal   gt31_txphinit_i                 : std_logic;
    signal   gt31_txphinitdone_i             : std_logic;
    signal   gt31_run_tx_phalignment_i       : std_logic;
    signal   gt31_rst_tx_phalignment_i       : std_logic;
    signal   gt31_tx_phalignment_done_i      : std_logic;
    signal   gt31_txsyncallin_i              : std_logic;
    signal   gt31_txsyncin_i                 : std_logic;
    signal   gt31_txsyncmode_i               : std_logic;
    signal   gt31_txsyncout_i                : std_logic;
    signal   gt31_txsyncdone_i               : std_logic;

    signal   gt31_txoutclk_i                 : std_logic;
    signal   gt31_rxoutclk_i                 : std_logic;
    signal   gt31_rxoutclk_i2                : std_logic;
    signal   gt31_txoutclk_i2                : std_logic;
    signal   gt31_recclk_stable_i            : std_logic;
    signal   gt31_rx_cdrlocked               : std_logic;
    signal   gt31_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal   gt31_rxphaligndone_i            : std_logic;
    signal   gt31_rxdlysreset_i              : std_logic;
    signal   gt31_rxdlysresetdone_i          : std_logic;
    signal   gt31_rxphdlyreset_i             : std_logic;
    signal   gt31_rxphalignen_i              : std_logic;
    signal   gt31_rxdlyen_i                  : std_logic;
    signal   gt31_rxphalign_i                : std_logic;
    signal   gt31_run_rx_phalignment_i       : std_logic;
    signal   gt31_rst_rx_phalignment_i       : std_logic;
    signal   gt31_rx_phalignment_done_i      : std_logic;
    signal   gt31_rxsyncallin_i              : std_logic;
    signal   gt31_rxsyncin_i                 : std_logic;
    signal   gt31_rxsyncmode_i               : std_logic;
    signal   gt31_rxsyncout_i                : std_logic;
    signal   gt31_rxsyncdone_i               : std_logic;



    --------------------------- TX Buffer Bypass Signals --------------------
    signal  mstr0_txsyncallin_i  :   std_logic;
    signal  U0_TXDLYEN           :   std_logic_vector(11 downto 0);
    signal  U0_TXDLYSRESET       :   std_logic_vector(11 downto 0);
    signal  U0_TXDLYSRESETDONE   :   std_logic_vector(11 downto 0);
    signal  U0_TXPHINIT          :   std_logic_vector(11 downto 0);
    signal  U0_TXPHINITDONE      :   std_logic_vector(11 downto 0);
    signal  U0_TXPHALIGN         :   std_logic_vector(11 downto 0);
    signal  U0_TXPHALIGNDONE     :   std_logic_vector(11 downto 0);
    signal  U0_run_tx_phalignment_i :   std_logic;
    signal  U0_rst_tx_phalignment_i :   std_logic;

    signal  mstr12_txsyncallin_i  :   std_logic;
    signal  U12_TXDLYEN           :   std_logic_vector(11 downto 0);
    signal  U12_TXDLYSRESET       :   std_logic_vector(11 downto 0);
    signal  U12_TXDLYSRESETDONE   :   std_logic_vector(11 downto 0);
    signal  U12_TXPHINIT          :   std_logic_vector(11 downto 0);
    signal  U12_TXPHINITDONE      :   std_logic_vector(11 downto 0);
    signal  U12_TXPHALIGN         :   std_logic_vector(11 downto 0);
    signal  U12_TXPHALIGNDONE     :   std_logic_vector(11 downto 0);
    signal  U12_run_tx_phalignment_i :   std_logic;
    signal  U12_rst_tx_phalignment_i :   std_logic;

    signal  mstr24_txsyncallin_i  :   std_logic;
    signal  U24_TXDLYEN           :   std_logic_vector(7 downto 0);
    signal  U24_TXDLYSRESET       :   std_logic_vector(7 downto 0);
    signal  U24_TXDLYSRESETDONE   :   std_logic_vector(7 downto 0);
    signal  U24_TXPHINIT          :   std_logic_vector(7 downto 0);
    signal  U24_TXPHINITDONE      :   std_logic_vector(7 downto 0);
    signal  U24_TXPHALIGN         :   std_logic_vector(7 downto 0);
    signal  U24_TXPHALIGNDONE     :   std_logic_vector(7 downto 0);
    signal  U24_run_tx_phalignment_i :   std_logic;
    signal  U24_rst_tx_phalignment_i :   std_logic;


    --------------------------- RX Buffer Bypass Signals --------------------
    signal   rxmstr0_rxsyncallin_i :   std_logic;
    signal  U0_RXDLYEN           :   std_logic_vector(11 downto 0);
    signal  U0_RXDLYSRESET       :   std_logic_vector(11 downto 0);
    signal  U0_RXDLYSRESETDONE   :   std_logic_vector(11 downto 0);
    signal  U0_RXPHALIGN         :   std_logic_vector(11 downto 0);
    signal  U0_RXPHALIGNDONE     :   std_logic_vector(11 downto 0);
    signal  U0_run_rx_phalignment_i :   std_logic;
    signal  U0_rst_rx_phalignment_i :   std_logic;

    signal   rxmstr12_rxsyncallin_i :   std_logic;
    signal  U12_RXDLYEN           :   std_logic_vector(11 downto 0);
    signal  U12_RXDLYSRESET       :   std_logic_vector(11 downto 0);
    signal  U12_RXDLYSRESETDONE   :   std_logic_vector(11 downto 0);
    signal  U12_RXPHALIGN         :   std_logic_vector(11 downto 0);
    signal  U12_RXPHALIGNDONE     :   std_logic_vector(11 downto 0);
    signal  U12_run_rx_phalignment_i :   std_logic;
    signal  U12_rst_rx_phalignment_i :   std_logic;

    signal   rxmstr24_rxsyncallin_i :   std_logic;
    signal  U24_RXDLYEN           :   std_logic_vector(7 downto 0);
    signal  U24_RXDLYSRESET       :   std_logic_vector(7 downto 0);
    signal  U24_RXDLYSRESETDONE   :   std_logic_vector(7 downto 0);
    signal  U24_RXPHALIGN         :   std_logic_vector(7 downto 0);
    signal  U24_RXPHALIGNDONE     :   std_logic_vector(7 downto 0);
    signal  U24_run_rx_phalignment_i :   std_logic;
    signal  U24_rst_rx_phalignment_i :   std_logic;



    signal      rx_cdrlocked                    : std_logic;


 


--**************************** Main Body of Code *******************************
begin
    --  Static signal Assigments
    tied_to_ground_i                             <= '0';
    tied_to_vcc_i                                <= '1';

    ----------------------------- The GT Wrapper -----------------------------
    
    -- Use the instantiation template in the example directory to add the GT wrapper to your design.
    -- In this example, the wrapper is wired up for basic operation with a frame generator and frame 
    -- checker. The GTs will reset, then attempt to align and transmit data. If channel bonding is 
    -- enabled, bonding should occur after alignment.


    gtwizard_0_i : gtwizard_0_multi_gt
    generic map
    (
        EXAMPLE_SIMULATION              =>      EXAMPLE_SIMULATION,
        WRAPPER_SIM_GTRESET_SPEEDUP     =>      EXAMPLE_SIM_GTRESET_SPEEDUP
    )
    port map
    (
        GT0_DRP_BUSY_OUT                =>      GT0_DRP_BUSY_OUT,
        GT0_RXPMARESETDONE_OUT          =>      gt0_rxpmaresetdone_i,
        GT0_TXPMARESETDONE_OUT          =>      gt0_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT0  (X1Y4)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt0_drpaddr_in                  =>      gt0_drpaddr_in,
        gt0_drpclk_in                   =>      gt0_drpclk_in,
        gt0_drpdi_in                    =>      gt0_drpdi_in,
        gt0_drpdo_out                   =>      gt0_drpdo_out,
        gt0_drpen_in                    =>      gt0_drpen_in,
        gt0_drprdy_out                  =>      gt0_drprdy_out,
        gt0_drpwe_in                    =>      gt0_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt0_eyescanreset_in             =>      gt0_eyescanreset_in,
        gt0_rxuserrdy_in                =>      gt0_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt0_eyescandataerror_out        =>      gt0_eyescandataerror_out,
        gt0_eyescantrigger_in           =>      gt0_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt0_rxslide_in                  =>      gt0_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt0_dmonitorout_out             =>      gt0_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt0_rxusrclk_in                 =>      gt0_rxusrclk_in,
        gt0_rxusrclk2_in                =>      gt0_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt0_rxdata_out                  =>      gt0_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt0_rxdisperr_out               =>      gt0_rxdisperr_out,
        gt0_rxnotintable_out            =>      gt0_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt0_gthrxn_in                   =>      gt0_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt0_rxdlyen_in                  =>      gt0_rxdlyen_i,
        gt0_rxdlysreset_in              =>      gt0_rxdlysreset_i,
        gt0_rxdlysresetdone_out         =>      gt0_rxdlysresetdone_i,
        gt0_rxphalign_in                =>      gt0_rxphalign_i,
        gt0_rxphaligndone_out           =>      gt0_rxphaligndone_i,
        gt0_rxphalignen_in              =>      gt0_rxphalignen_i,
        gt0_rxphdlyreset_in             =>      gt0_rxphdlyreset_i,
        gt0_rxphmonitor_out             =>      gt0_rxphmonitor_out,
        gt0_rxphslipmonitor_out         =>      gt0_rxphslipmonitor_out,
        gt0_rxsyncallin_in              =>      gt0_rxsyncallin_i,
        gt0_rxsyncdone_out              =>      gt0_rxsyncdone_i,
        gt0_rxsyncin_in                 =>      gt0_rxsyncin_i,
        gt0_rxsyncmode_in               =>      gt0_rxsyncmode_i,
        gt0_rxsyncout_out               =>      gt0_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt0_rxbyteisaligned_out         =>      gt0_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt0_rxlpmhfhold_in              =>      gt0_rxlpmhfhold_i,
        gt0_rxlpmlfhold_in              =>      gt0_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt0_rxmonitorout_out            =>      gt0_rxmonitorout_out,
        gt0_rxmonitorsel_in             =>      gt0_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt0_rxoutclk_out                =>      gt0_rxoutclk_i,
        gt0_rxoutclkfabric_out          =>      gt0_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt0_gtrxreset_in                =>      gt0_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt0_rxcharisk_out               =>      gt0_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt0_gthrxp_in                   =>      gt0_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt0_rxresetdone_out             =>      gt0_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt0_gttxreset_in                =>      gt0_gttxreset_i,
        gt0_txuserrdy_in                =>      gt0_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt0_txusrclk_in                 =>      gt0_txusrclk_in,
        gt0_txusrclk2_in                =>      gt0_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt0_txdlyen_in                  =>      gt0_txdlyen_i,
        gt0_txdlysreset_in              =>      gt0_txdlysreset_i,
        gt0_txdlysresetdone_out         =>      gt0_txdlysresetdone_i,
        gt0_txphalign_in                =>      gt0_txphalign_i,
        gt0_txphaligndone_out           =>      gt0_txphaligndone_i,
        gt0_txphalignen_in              =>      gt0_txphalignen_i,
        gt0_txphdlyreset_in             =>      gt0_txphdlyreset_i,
        gt0_txphinit_in                 =>      gt0_txphinit_i,
        gt0_txphinitdone_out            =>      gt0_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt0_txdata_in                   =>      gt0_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt0_gthtxn_out                  =>      gt0_gthtxn_out,
        gt0_gthtxp_out                  =>      gt0_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt0_txoutclk_out                =>      gt0_txoutclk_i,
        gt0_txoutclkfabric_out          =>      gt0_txoutclkfabric_out,
        gt0_txoutclkpcs_out             =>      gt0_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt0_txresetdone_out             =>      gt0_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt0_txcharisk_in                =>      gt0_txcharisk_in,


        GT1_DRP_BUSY_OUT                =>      GT1_DRP_BUSY_OUT,
        GT1_RXPMARESETDONE_OUT          =>      gt1_rxpmaresetdone_i,
        GT1_TXPMARESETDONE_OUT          =>      gt1_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT1  (X1Y5)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt1_drpaddr_in                  =>      gt1_drpaddr_in,
        gt1_drpclk_in                   =>      gt1_drpclk_in,
        gt1_drpdi_in                    =>      gt1_drpdi_in,
        gt1_drpdo_out                   =>      gt1_drpdo_out,
        gt1_drpen_in                    =>      gt1_drpen_in,
        gt1_drprdy_out                  =>      gt1_drprdy_out,
        gt1_drpwe_in                    =>      gt1_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt1_eyescanreset_in             =>      gt1_eyescanreset_in,
        gt1_rxuserrdy_in                =>      gt1_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt1_eyescandataerror_out        =>      gt1_eyescandataerror_out,
        gt1_eyescantrigger_in           =>      gt1_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt1_rxslide_in                  =>      gt1_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt1_dmonitorout_out             =>      gt1_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt1_rxusrclk_in                 =>      gt1_rxusrclk_in,
        gt1_rxusrclk2_in                =>      gt1_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt1_rxdata_out                  =>      gt1_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt1_rxdisperr_out               =>      gt1_rxdisperr_out,
        gt1_rxnotintable_out            =>      gt1_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt1_gthrxn_in                   =>      gt1_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt1_rxdlyen_in                  =>      gt1_rxdlyen_i,
        gt1_rxdlysreset_in              =>      gt1_rxdlysreset_i,
        gt1_rxdlysresetdone_out         =>      gt1_rxdlysresetdone_i,
        gt1_rxphalign_in                =>      gt1_rxphalign_i,
        gt1_rxphaligndone_out           =>      gt1_rxphaligndone_i,
        gt1_rxphalignen_in              =>      gt1_rxphalignen_i,
        gt1_rxphdlyreset_in             =>      gt1_rxphdlyreset_i,
        gt1_rxphmonitor_out             =>      gt1_rxphmonitor_out,
        gt1_rxphslipmonitor_out         =>      gt1_rxphslipmonitor_out,
        gt1_rxsyncallin_in              =>      gt1_rxsyncallin_i,
        gt1_rxsyncdone_out              =>      gt1_rxsyncdone_i,
        gt1_rxsyncin_in                 =>      gt1_rxsyncin_i,
        gt1_rxsyncmode_in               =>      gt1_rxsyncmode_i,
        gt1_rxsyncout_out               =>      gt1_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt1_rxbyteisaligned_out         =>      gt1_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt1_rxlpmhfhold_in              =>      gt1_rxlpmhfhold_i,
        gt1_rxlpmlfhold_in              =>      gt1_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt1_rxmonitorout_out            =>      gt1_rxmonitorout_out,
        gt1_rxmonitorsel_in             =>      gt1_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt1_rxoutclk_out                =>      gt1_rxoutclk_i,
        gt1_rxoutclkfabric_out          =>      gt1_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt1_gtrxreset_in                =>      gt1_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt1_rxcharisk_out               =>      gt1_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt1_gthrxp_in                   =>      gt1_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt1_rxresetdone_out             =>      gt1_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt1_gttxreset_in                =>      gt1_gttxreset_i,
        gt1_txuserrdy_in                =>      gt1_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt1_txusrclk_in                 =>      gt1_txusrclk_in,
        gt1_txusrclk2_in                =>      gt1_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt1_txdlyen_in                  =>      gt1_txdlyen_i,
        gt1_txdlysreset_in              =>      gt1_txdlysreset_i,
        gt1_txdlysresetdone_out         =>      gt1_txdlysresetdone_i,
        gt1_txphalign_in                =>      gt1_txphalign_i,
        gt1_txphaligndone_out           =>      gt1_txphaligndone_i,
        gt1_txphalignen_in              =>      gt1_txphalignen_i,
        gt1_txphdlyreset_in             =>      gt1_txphdlyreset_i,
        gt1_txphinit_in                 =>      gt1_txphinit_i,
        gt1_txphinitdone_out            =>      gt1_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt1_txdata_in                   =>      gt1_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt1_gthtxn_out                  =>      gt1_gthtxn_out,
        gt1_gthtxp_out                  =>      gt1_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt1_txoutclk_out                =>      gt1_txoutclk_i,
        gt1_txoutclkfabric_out          =>      gt1_txoutclkfabric_out,
        gt1_txoutclkpcs_out             =>      gt1_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt1_txresetdone_out             =>      gt1_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt1_txcharisk_in                =>      gt1_txcharisk_in,


        GT2_DRP_BUSY_OUT                =>      GT2_DRP_BUSY_OUT,
        GT2_RXPMARESETDONE_OUT          =>      gt2_rxpmaresetdone_i,
        GT2_TXPMARESETDONE_OUT          =>      gt2_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT2  (X1Y6)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt2_drpaddr_in                  =>      gt2_drpaddr_in,
        gt2_drpclk_in                   =>      gt2_drpclk_in,
        gt2_drpdi_in                    =>      gt2_drpdi_in,
        gt2_drpdo_out                   =>      gt2_drpdo_out,
        gt2_drpen_in                    =>      gt2_drpen_in,
        gt2_drprdy_out                  =>      gt2_drprdy_out,
        gt2_drpwe_in                    =>      gt2_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt2_eyescanreset_in             =>      gt2_eyescanreset_in,
        gt2_rxuserrdy_in                =>      gt2_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt2_eyescandataerror_out        =>      gt2_eyescandataerror_out,
        gt2_eyescantrigger_in           =>      gt2_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt2_rxslide_in                  =>      gt2_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt2_dmonitorout_out             =>      gt2_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt2_rxusrclk_in                 =>      gt2_rxusrclk_in,
        gt2_rxusrclk2_in                =>      gt2_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt2_rxdata_out                  =>      gt2_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt2_rxdisperr_out               =>      gt2_rxdisperr_out,
        gt2_rxnotintable_out            =>      gt2_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt2_gthrxn_in                   =>      gt2_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt2_rxdlyen_in                  =>      gt2_rxdlyen_i,
        gt2_rxdlysreset_in              =>      gt2_rxdlysreset_i,
        gt2_rxdlysresetdone_out         =>      gt2_rxdlysresetdone_i,
        gt2_rxphalign_in                =>      gt2_rxphalign_i,
        gt2_rxphaligndone_out           =>      gt2_rxphaligndone_i,
        gt2_rxphalignen_in              =>      gt2_rxphalignen_i,
        gt2_rxphdlyreset_in             =>      gt2_rxphdlyreset_i,
        gt2_rxphmonitor_out             =>      gt2_rxphmonitor_out,
        gt2_rxphslipmonitor_out         =>      gt2_rxphslipmonitor_out,
        gt2_rxsyncallin_in              =>      gt2_rxsyncallin_i,
        gt2_rxsyncdone_out              =>      gt2_rxsyncdone_i,
        gt2_rxsyncin_in                 =>      gt2_rxsyncin_i,
        gt2_rxsyncmode_in               =>      gt2_rxsyncmode_i,
        gt2_rxsyncout_out               =>      gt2_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt2_rxbyteisaligned_out         =>      gt2_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt2_rxlpmhfhold_in              =>      gt2_rxlpmhfhold_i,
        gt2_rxlpmlfhold_in              =>      gt2_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt2_rxmonitorout_out            =>      gt2_rxmonitorout_out,
        gt2_rxmonitorsel_in             =>      gt2_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt2_rxoutclk_out                =>      gt2_rxoutclk_i,
        gt2_rxoutclkfabric_out          =>      gt2_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt2_gtrxreset_in                =>      gt2_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt2_rxcharisk_out               =>      gt2_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt2_gthrxp_in                   =>      gt2_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt2_rxresetdone_out             =>      gt2_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt2_gttxreset_in                =>      gt2_gttxreset_i,
        gt2_txuserrdy_in                =>      gt2_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt2_txusrclk_in                 =>      gt2_txusrclk_in,
        gt2_txusrclk2_in                =>      gt2_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt2_txdlyen_in                  =>      gt2_txdlyen_i,
        gt2_txdlysreset_in              =>      gt2_txdlysreset_i,
        gt2_txdlysresetdone_out         =>      gt2_txdlysresetdone_i,
        gt2_txphalign_in                =>      gt2_txphalign_i,
        gt2_txphaligndone_out           =>      gt2_txphaligndone_i,
        gt2_txphalignen_in              =>      gt2_txphalignen_i,
        gt2_txphdlyreset_in             =>      gt2_txphdlyreset_i,
        gt2_txphinit_in                 =>      gt2_txphinit_i,
        gt2_txphinitdone_out            =>      gt2_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt2_txdata_in                   =>      gt2_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt2_gthtxn_out                  =>      gt2_gthtxn_out,
        gt2_gthtxp_out                  =>      gt2_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt2_txoutclk_out                =>      gt2_txoutclk_i,
        gt2_txoutclkfabric_out          =>      gt2_txoutclkfabric_out,
        gt2_txoutclkpcs_out             =>      gt2_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt2_txresetdone_out             =>      gt2_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt2_txcharisk_in                =>      gt2_txcharisk_in,


        GT3_DRP_BUSY_OUT                =>      GT3_DRP_BUSY_OUT,
        GT3_RXPMARESETDONE_OUT          =>      gt3_rxpmaresetdone_i,
        GT3_TXPMARESETDONE_OUT          =>      gt3_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT3  (X1Y7)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt3_drpaddr_in                  =>      gt3_drpaddr_in,
        gt3_drpclk_in                   =>      gt3_drpclk_in,
        gt3_drpdi_in                    =>      gt3_drpdi_in,
        gt3_drpdo_out                   =>      gt3_drpdo_out,
        gt3_drpen_in                    =>      gt3_drpen_in,
        gt3_drprdy_out                  =>      gt3_drprdy_out,
        gt3_drpwe_in                    =>      gt3_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt3_eyescanreset_in             =>      gt3_eyescanreset_in,
        gt3_rxuserrdy_in                =>      gt3_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt3_eyescandataerror_out        =>      gt3_eyescandataerror_out,
        gt3_eyescantrigger_in           =>      gt3_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt3_rxslide_in                  =>      gt3_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt3_dmonitorout_out             =>      gt3_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt3_rxusrclk_in                 =>      gt3_rxusrclk_in,
        gt3_rxusrclk2_in                =>      gt3_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt3_rxdata_out                  =>      gt3_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt3_rxdisperr_out               =>      gt3_rxdisperr_out,
        gt3_rxnotintable_out            =>      gt3_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt3_gthrxn_in                   =>      gt3_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt3_rxdlyen_in                  =>      gt3_rxdlyen_i,
        gt3_rxdlysreset_in              =>      gt3_rxdlysreset_i,
        gt3_rxdlysresetdone_out         =>      gt3_rxdlysresetdone_i,
        gt3_rxphalign_in                =>      gt3_rxphalign_i,
        gt3_rxphaligndone_out           =>      gt3_rxphaligndone_i,
        gt3_rxphalignen_in              =>      gt3_rxphalignen_i,
        gt3_rxphdlyreset_in             =>      gt3_rxphdlyreset_i,
        gt3_rxphmonitor_out             =>      gt3_rxphmonitor_out,
        gt3_rxphslipmonitor_out         =>      gt3_rxphslipmonitor_out,
        gt3_rxsyncallin_in              =>      gt3_rxsyncallin_i,
        gt3_rxsyncdone_out              =>      gt3_rxsyncdone_i,
        gt3_rxsyncin_in                 =>      gt3_rxsyncin_i,
        gt3_rxsyncmode_in               =>      gt3_rxsyncmode_i,
        gt3_rxsyncout_out               =>      gt3_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt3_rxbyteisaligned_out         =>      gt3_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt3_rxlpmhfhold_in              =>      gt3_rxlpmhfhold_i,
        gt3_rxlpmlfhold_in              =>      gt3_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt3_rxmonitorout_out            =>      gt3_rxmonitorout_out,
        gt3_rxmonitorsel_in             =>      gt3_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt3_rxoutclk_out                =>      gt3_rxoutclk_i,
        gt3_rxoutclkfabric_out          =>      gt3_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt3_gtrxreset_in                =>      gt3_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt3_rxcharisk_out               =>      gt3_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt3_gthrxp_in                   =>      gt3_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt3_rxresetdone_out             =>      gt3_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt3_gttxreset_in                =>      gt3_gttxreset_i,
        gt3_txuserrdy_in                =>      gt3_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt3_txusrclk_in                 =>      gt3_txusrclk_in,
        gt3_txusrclk2_in                =>      gt3_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt3_txdlyen_in                  =>      gt3_txdlyen_i,
        gt3_txdlysreset_in              =>      gt3_txdlysreset_i,
        gt3_txdlysresetdone_out         =>      gt3_txdlysresetdone_i,
        gt3_txphalign_in                =>      gt3_txphalign_i,
        gt3_txphaligndone_out           =>      gt3_txphaligndone_i,
        gt3_txphalignen_in              =>      gt3_txphalignen_i,
        gt3_txphdlyreset_in             =>      gt3_txphdlyreset_i,
        gt3_txphinit_in                 =>      gt3_txphinit_i,
        gt3_txphinitdone_out            =>      gt3_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt3_txdata_in                   =>      gt3_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt3_gthtxn_out                  =>      gt3_gthtxn_out,
        gt3_gthtxp_out                  =>      gt3_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt3_txoutclk_out                =>      gt3_txoutclk_i,
        gt3_txoutclkfabric_out          =>      gt3_txoutclkfabric_out,
        gt3_txoutclkpcs_out             =>      gt3_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt3_txresetdone_out             =>      gt3_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt3_txcharisk_in                =>      gt3_txcharisk_in,


        GT4_DRP_BUSY_OUT                =>      GT4_DRP_BUSY_OUT,
        GT4_RXPMARESETDONE_OUT          =>      gt4_rxpmaresetdone_i,
        GT4_TXPMARESETDONE_OUT          =>      gt4_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT4  (X1Y8)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt4_drpaddr_in                  =>      gt4_drpaddr_in,
        gt4_drpclk_in                   =>      gt4_drpclk_in,
        gt4_drpdi_in                    =>      gt4_drpdi_in,
        gt4_drpdo_out                   =>      gt4_drpdo_out,
        gt4_drpen_in                    =>      gt4_drpen_in,
        gt4_drprdy_out                  =>      gt4_drprdy_out,
        gt4_drpwe_in                    =>      gt4_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt4_eyescanreset_in             =>      gt4_eyescanreset_in,
        gt4_rxuserrdy_in                =>      gt4_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt4_eyescandataerror_out        =>      gt4_eyescandataerror_out,
        gt4_eyescantrigger_in           =>      gt4_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt4_rxslide_in                  =>      gt4_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt4_dmonitorout_out             =>      gt4_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt4_rxusrclk_in                 =>      gt4_rxusrclk_in,
        gt4_rxusrclk2_in                =>      gt4_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt4_rxdata_out                  =>      gt4_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt4_rxdisperr_out               =>      gt4_rxdisperr_out,
        gt4_rxnotintable_out            =>      gt4_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt4_gthrxn_in                   =>      gt4_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt4_rxdlyen_in                  =>      gt4_rxdlyen_i,
        gt4_rxdlysreset_in              =>      gt4_rxdlysreset_i,
        gt4_rxdlysresetdone_out         =>      gt4_rxdlysresetdone_i,
        gt4_rxphalign_in                =>      gt4_rxphalign_i,
        gt4_rxphaligndone_out           =>      gt4_rxphaligndone_i,
        gt4_rxphalignen_in              =>      gt4_rxphalignen_i,
        gt4_rxphdlyreset_in             =>      gt4_rxphdlyreset_i,
        gt4_rxphmonitor_out             =>      gt4_rxphmonitor_out,
        gt4_rxphslipmonitor_out         =>      gt4_rxphslipmonitor_out,
        gt4_rxsyncallin_in              =>      gt4_rxsyncallin_i,
        gt4_rxsyncdone_out              =>      gt4_rxsyncdone_i,
        gt4_rxsyncin_in                 =>      gt4_rxsyncin_i,
        gt4_rxsyncmode_in               =>      gt4_rxsyncmode_i,
        gt4_rxsyncout_out               =>      gt4_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt4_rxbyteisaligned_out         =>      gt4_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt4_rxlpmhfhold_in              =>      gt4_rxlpmhfhold_i,
        gt4_rxlpmlfhold_in              =>      gt4_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt4_rxmonitorout_out            =>      gt4_rxmonitorout_out,
        gt4_rxmonitorsel_in             =>      gt4_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt4_rxoutclk_out                =>      gt4_rxoutclk_i,
        gt4_rxoutclkfabric_out          =>      gt4_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt4_gtrxreset_in                =>      gt4_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt4_rxcharisk_out               =>      gt4_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt4_gthrxp_in                   =>      gt4_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt4_rxresetdone_out             =>      gt4_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt4_gttxreset_in                =>      gt4_gttxreset_i,
        gt4_txuserrdy_in                =>      gt4_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt4_txusrclk_in                 =>      gt4_txusrclk_in,
        gt4_txusrclk2_in                =>      gt4_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt4_txdlyen_in                  =>      gt4_txdlyen_i,
        gt4_txdlysreset_in              =>      gt4_txdlysreset_i,
        gt4_txdlysresetdone_out         =>      gt4_txdlysresetdone_i,
        gt4_txphalign_in                =>      gt4_txphalign_i,
        gt4_txphaligndone_out           =>      gt4_txphaligndone_i,
        gt4_txphalignen_in              =>      gt4_txphalignen_i,
        gt4_txphdlyreset_in             =>      gt4_txphdlyreset_i,
        gt4_txphinit_in                 =>      gt4_txphinit_i,
        gt4_txphinitdone_out            =>      gt4_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt4_txdata_in                   =>      gt4_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt4_gthtxn_out                  =>      gt4_gthtxn_out,
        gt4_gthtxp_out                  =>      gt4_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt4_txoutclk_out                =>      gt4_txoutclk_i,
        gt4_txoutclkfabric_out          =>      gt4_txoutclkfabric_out,
        gt4_txoutclkpcs_out             =>      gt4_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt4_txresetdone_out             =>      gt4_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt4_txcharisk_in                =>      gt4_txcharisk_in,


        GT5_DRP_BUSY_OUT                =>      GT5_DRP_BUSY_OUT,
        GT5_RXPMARESETDONE_OUT          =>      gt5_rxpmaresetdone_i,
        GT5_TXPMARESETDONE_OUT          =>      gt5_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT5  (X1Y9)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt5_drpaddr_in                  =>      gt5_drpaddr_in,
        gt5_drpclk_in                   =>      gt5_drpclk_in,
        gt5_drpdi_in                    =>      gt5_drpdi_in,
        gt5_drpdo_out                   =>      gt5_drpdo_out,
        gt5_drpen_in                    =>      gt5_drpen_in,
        gt5_drprdy_out                  =>      gt5_drprdy_out,
        gt5_drpwe_in                    =>      gt5_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt5_eyescanreset_in             =>      gt5_eyescanreset_in,
        gt5_rxuserrdy_in                =>      gt5_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt5_eyescandataerror_out        =>      gt5_eyescandataerror_out,
        gt5_eyescantrigger_in           =>      gt5_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt5_rxslide_in                  =>      gt5_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt5_dmonitorout_out             =>      gt5_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt5_rxusrclk_in                 =>      gt5_rxusrclk_in,
        gt5_rxusrclk2_in                =>      gt5_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt5_rxdata_out                  =>      gt5_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt5_rxdisperr_out               =>      gt5_rxdisperr_out,
        gt5_rxnotintable_out            =>      gt5_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt5_gthrxn_in                   =>      gt5_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt5_rxdlyen_in                  =>      gt5_rxdlyen_i,
        gt5_rxdlysreset_in              =>      gt5_rxdlysreset_i,
        gt5_rxdlysresetdone_out         =>      gt5_rxdlysresetdone_i,
        gt5_rxphalign_in                =>      gt5_rxphalign_i,
        gt5_rxphaligndone_out           =>      gt5_rxphaligndone_i,
        gt5_rxphalignen_in              =>      gt5_rxphalignen_i,
        gt5_rxphdlyreset_in             =>      gt5_rxphdlyreset_i,
        gt5_rxphmonitor_out             =>      gt5_rxphmonitor_out,
        gt5_rxphslipmonitor_out         =>      gt5_rxphslipmonitor_out,
        gt5_rxsyncallin_in              =>      gt5_rxsyncallin_i,
        gt5_rxsyncdone_out              =>      gt5_rxsyncdone_i,
        gt5_rxsyncin_in                 =>      gt5_rxsyncin_i,
        gt5_rxsyncmode_in               =>      gt5_rxsyncmode_i,
        gt5_rxsyncout_out               =>      gt5_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt5_rxbyteisaligned_out         =>      gt5_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt5_rxlpmhfhold_in              =>      gt5_rxlpmhfhold_i,
        gt5_rxlpmlfhold_in              =>      gt5_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt5_rxmonitorout_out            =>      gt5_rxmonitorout_out,
        gt5_rxmonitorsel_in             =>      gt5_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt5_rxoutclk_out                =>      gt5_rxoutclk_i,
        gt5_rxoutclkfabric_out          =>      gt5_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt5_gtrxreset_in                =>      gt5_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt5_rxcharisk_out               =>      gt5_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt5_gthrxp_in                   =>      gt5_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt5_rxresetdone_out             =>      gt5_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt5_gttxreset_in                =>      gt5_gttxreset_i,
        gt5_txuserrdy_in                =>      gt5_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt5_txusrclk_in                 =>      gt5_txusrclk_in,
        gt5_txusrclk2_in                =>      gt5_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt5_txdlyen_in                  =>      gt5_txdlyen_i,
        gt5_txdlysreset_in              =>      gt5_txdlysreset_i,
        gt5_txdlysresetdone_out         =>      gt5_txdlysresetdone_i,
        gt5_txphalign_in                =>      gt5_txphalign_i,
        gt5_txphaligndone_out           =>      gt5_txphaligndone_i,
        gt5_txphalignen_in              =>      gt5_txphalignen_i,
        gt5_txphdlyreset_in             =>      gt5_txphdlyreset_i,
        gt5_txphinit_in                 =>      gt5_txphinit_i,
        gt5_txphinitdone_out            =>      gt5_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt5_txdata_in                   =>      gt5_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt5_gthtxn_out                  =>      gt5_gthtxn_out,
        gt5_gthtxp_out                  =>      gt5_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt5_txoutclk_out                =>      gt5_txoutclk_i,
        gt5_txoutclkfabric_out          =>      gt5_txoutclkfabric_out,
        gt5_txoutclkpcs_out             =>      gt5_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt5_txresetdone_out             =>      gt5_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt5_txcharisk_in                =>      gt5_txcharisk_in,


        GT6_DRP_BUSY_OUT                =>      GT6_DRP_BUSY_OUT,
        GT6_RXPMARESETDONE_OUT          =>      gt6_rxpmaresetdone_i,
        GT6_TXPMARESETDONE_OUT          =>      gt6_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT6  (X1Y10)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt6_drpaddr_in                  =>      gt6_drpaddr_in,
        gt6_drpclk_in                   =>      gt6_drpclk_in,
        gt6_drpdi_in                    =>      gt6_drpdi_in,
        gt6_drpdo_out                   =>      gt6_drpdo_out,
        gt6_drpen_in                    =>      gt6_drpen_in,
        gt6_drprdy_out                  =>      gt6_drprdy_out,
        gt6_drpwe_in                    =>      gt6_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt6_eyescanreset_in             =>      gt6_eyescanreset_in,
        gt6_rxuserrdy_in                =>      gt6_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt6_eyescandataerror_out        =>      gt6_eyescandataerror_out,
        gt6_eyescantrigger_in           =>      gt6_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt6_rxslide_in                  =>      gt6_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt6_dmonitorout_out             =>      gt6_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt6_rxusrclk_in                 =>      gt6_rxusrclk_in,
        gt6_rxusrclk2_in                =>      gt6_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt6_rxdata_out                  =>      gt6_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt6_rxdisperr_out               =>      gt6_rxdisperr_out,
        gt6_rxnotintable_out            =>      gt6_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt6_gthrxn_in                   =>      gt6_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt6_rxdlyen_in                  =>      gt6_rxdlyen_i,
        gt6_rxdlysreset_in              =>      gt6_rxdlysreset_i,
        gt6_rxdlysresetdone_out         =>      gt6_rxdlysresetdone_i,
        gt6_rxphalign_in                =>      gt6_rxphalign_i,
        gt6_rxphaligndone_out           =>      gt6_rxphaligndone_i,
        gt6_rxphalignen_in              =>      gt6_rxphalignen_i,
        gt6_rxphdlyreset_in             =>      gt6_rxphdlyreset_i,
        gt6_rxphmonitor_out             =>      gt6_rxphmonitor_out,
        gt6_rxphslipmonitor_out         =>      gt6_rxphslipmonitor_out,
        gt6_rxsyncallin_in              =>      gt6_rxsyncallin_i,
        gt6_rxsyncdone_out              =>      gt6_rxsyncdone_i,
        gt6_rxsyncin_in                 =>      gt6_rxsyncin_i,
        gt6_rxsyncmode_in               =>      gt6_rxsyncmode_i,
        gt6_rxsyncout_out               =>      gt6_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt6_rxbyteisaligned_out         =>      gt6_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt6_rxlpmhfhold_in              =>      gt6_rxlpmhfhold_i,
        gt6_rxlpmlfhold_in              =>      gt6_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt6_rxmonitorout_out            =>      gt6_rxmonitorout_out,
        gt6_rxmonitorsel_in             =>      gt6_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt6_rxoutclk_out                =>      gt6_rxoutclk_i,
        gt6_rxoutclkfabric_out          =>      gt6_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt6_gtrxreset_in                =>      gt6_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt6_rxcharisk_out               =>      gt6_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt6_gthrxp_in                   =>      gt6_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt6_rxresetdone_out             =>      gt6_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt6_gttxreset_in                =>      gt6_gttxreset_i,
        gt6_txuserrdy_in                =>      gt6_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt6_txusrclk_in                 =>      gt6_txusrclk_in,
        gt6_txusrclk2_in                =>      gt6_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt6_txdlyen_in                  =>      gt6_txdlyen_i,
        gt6_txdlysreset_in              =>      gt6_txdlysreset_i,
        gt6_txdlysresetdone_out         =>      gt6_txdlysresetdone_i,
        gt6_txphalign_in                =>      gt6_txphalign_i,
        gt6_txphaligndone_out           =>      gt6_txphaligndone_i,
        gt6_txphalignen_in              =>      gt6_txphalignen_i,
        gt6_txphdlyreset_in             =>      gt6_txphdlyreset_i,
        gt6_txphinit_in                 =>      gt6_txphinit_i,
        gt6_txphinitdone_out            =>      gt6_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt6_txdata_in                   =>      gt6_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt6_gthtxn_out                  =>      gt6_gthtxn_out,
        gt6_gthtxp_out                  =>      gt6_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt6_txoutclk_out                =>      gt6_txoutclk_i,
        gt6_txoutclkfabric_out          =>      gt6_txoutclkfabric_out,
        gt6_txoutclkpcs_out             =>      gt6_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt6_txresetdone_out             =>      gt6_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt6_txcharisk_in                =>      gt6_txcharisk_in,


        GT7_DRP_BUSY_OUT                =>      GT7_DRP_BUSY_OUT,
        GT7_RXPMARESETDONE_OUT          =>      gt7_rxpmaresetdone_i,
        GT7_TXPMARESETDONE_OUT          =>      gt7_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT7  (X1Y11)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt7_drpaddr_in                  =>      gt7_drpaddr_in,
        gt7_drpclk_in                   =>      gt7_drpclk_in,
        gt7_drpdi_in                    =>      gt7_drpdi_in,
        gt7_drpdo_out                   =>      gt7_drpdo_out,
        gt7_drpen_in                    =>      gt7_drpen_in,
        gt7_drprdy_out                  =>      gt7_drprdy_out,
        gt7_drpwe_in                    =>      gt7_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt7_eyescanreset_in             =>      gt7_eyescanreset_in,
        gt7_rxuserrdy_in                =>      gt7_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt7_eyescandataerror_out        =>      gt7_eyescandataerror_out,
        gt7_eyescantrigger_in           =>      gt7_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt7_rxslide_in                  =>      gt7_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt7_dmonitorout_out             =>      gt7_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt7_rxusrclk_in                 =>      gt7_rxusrclk_in,
        gt7_rxusrclk2_in                =>      gt7_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt7_rxdata_out                  =>      gt7_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt7_rxdisperr_out               =>      gt7_rxdisperr_out,
        gt7_rxnotintable_out            =>      gt7_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt7_gthrxn_in                   =>      gt7_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt7_rxdlyen_in                  =>      gt7_rxdlyen_i,
        gt7_rxdlysreset_in              =>      gt7_rxdlysreset_i,
        gt7_rxdlysresetdone_out         =>      gt7_rxdlysresetdone_i,
        gt7_rxphalign_in                =>      gt7_rxphalign_i,
        gt7_rxphaligndone_out           =>      gt7_rxphaligndone_i,
        gt7_rxphalignen_in              =>      gt7_rxphalignen_i,
        gt7_rxphdlyreset_in             =>      gt7_rxphdlyreset_i,
        gt7_rxphmonitor_out             =>      gt7_rxphmonitor_out,
        gt7_rxphslipmonitor_out         =>      gt7_rxphslipmonitor_out,
        gt7_rxsyncallin_in              =>      gt7_rxsyncallin_i,
        gt7_rxsyncdone_out              =>      gt7_rxsyncdone_i,
        gt7_rxsyncin_in                 =>      gt7_rxsyncin_i,
        gt7_rxsyncmode_in               =>      gt7_rxsyncmode_i,
        gt7_rxsyncout_out               =>      gt7_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt7_rxbyteisaligned_out         =>      gt7_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt7_rxlpmhfhold_in              =>      gt7_rxlpmhfhold_i,
        gt7_rxlpmlfhold_in              =>      gt7_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt7_rxmonitorout_out            =>      gt7_rxmonitorout_out,
        gt7_rxmonitorsel_in             =>      gt7_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt7_rxoutclk_out                =>      gt7_rxoutclk_i,
        gt7_rxoutclkfabric_out          =>      gt7_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt7_gtrxreset_in                =>      gt7_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt7_rxcharisk_out               =>      gt7_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt7_gthrxp_in                   =>      gt7_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt7_rxresetdone_out             =>      gt7_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt7_gttxreset_in                =>      gt7_gttxreset_i,
        gt7_txuserrdy_in                =>      gt7_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt7_txusrclk_in                 =>      gt7_txusrclk_in,
        gt7_txusrclk2_in                =>      gt7_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt7_txdlyen_in                  =>      gt7_txdlyen_i,
        gt7_txdlysreset_in              =>      gt7_txdlysreset_i,
        gt7_txdlysresetdone_out         =>      gt7_txdlysresetdone_i,
        gt7_txphalign_in                =>      gt7_txphalign_i,
        gt7_txphaligndone_out           =>      gt7_txphaligndone_i,
        gt7_txphalignen_in              =>      gt7_txphalignen_i,
        gt7_txphdlyreset_in             =>      gt7_txphdlyreset_i,
        gt7_txphinit_in                 =>      gt7_txphinit_i,
        gt7_txphinitdone_out            =>      gt7_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt7_txdata_in                   =>      gt7_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt7_gthtxn_out                  =>      gt7_gthtxn_out,
        gt7_gthtxp_out                  =>      gt7_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt7_txoutclk_out                =>      gt7_txoutclk_i,
        gt7_txoutclkfabric_out          =>      gt7_txoutclkfabric_out,
        gt7_txoutclkpcs_out             =>      gt7_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt7_txresetdone_out             =>      gt7_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt7_txcharisk_in                =>      gt7_txcharisk_in,


        GT8_DRP_BUSY_OUT                =>      GT8_DRP_BUSY_OUT,
        GT8_RXPMARESETDONE_OUT          =>      gt8_rxpmaresetdone_i,
        GT8_TXPMARESETDONE_OUT          =>      gt8_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT8  (X1Y12)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt8_drpaddr_in                  =>      gt8_drpaddr_in,
        gt8_drpclk_in                   =>      gt8_drpclk_in,
        gt8_drpdi_in                    =>      gt8_drpdi_in,
        gt8_drpdo_out                   =>      gt8_drpdo_out,
        gt8_drpen_in                    =>      gt8_drpen_in,
        gt8_drprdy_out                  =>      gt8_drprdy_out,
        gt8_drpwe_in                    =>      gt8_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt8_eyescanreset_in             =>      gt8_eyescanreset_in,
        gt8_rxuserrdy_in                =>      gt8_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt8_eyescandataerror_out        =>      gt8_eyescandataerror_out,
        gt8_eyescantrigger_in           =>      gt8_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt8_rxslide_in                  =>      gt8_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt8_dmonitorout_out             =>      gt8_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt8_rxusrclk_in                 =>      gt8_rxusrclk_in,
        gt8_rxusrclk2_in                =>      gt8_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt8_rxdata_out                  =>      gt8_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt8_rxdisperr_out               =>      gt8_rxdisperr_out,
        gt8_rxnotintable_out            =>      gt8_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt8_gthrxn_in                   =>      gt8_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt8_rxdlyen_in                  =>      gt8_rxdlyen_i,
        gt8_rxdlysreset_in              =>      gt8_rxdlysreset_i,
        gt8_rxdlysresetdone_out         =>      gt8_rxdlysresetdone_i,
        gt8_rxphalign_in                =>      gt8_rxphalign_i,
        gt8_rxphaligndone_out           =>      gt8_rxphaligndone_i,
        gt8_rxphalignen_in              =>      gt8_rxphalignen_i,
        gt8_rxphdlyreset_in             =>      gt8_rxphdlyreset_i,
        gt8_rxphmonitor_out             =>      gt8_rxphmonitor_out,
        gt8_rxphslipmonitor_out         =>      gt8_rxphslipmonitor_out,
        gt8_rxsyncallin_in              =>      gt8_rxsyncallin_i,
        gt8_rxsyncdone_out              =>      gt8_rxsyncdone_i,
        gt8_rxsyncin_in                 =>      gt8_rxsyncin_i,
        gt8_rxsyncmode_in               =>      gt8_rxsyncmode_i,
        gt8_rxsyncout_out               =>      gt8_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt8_rxbyteisaligned_out         =>      gt8_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt8_rxlpmhfhold_in              =>      gt8_rxlpmhfhold_i,
        gt8_rxlpmlfhold_in              =>      gt8_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt8_rxmonitorout_out            =>      gt8_rxmonitorout_out,
        gt8_rxmonitorsel_in             =>      gt8_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt8_rxoutclk_out                =>      gt8_rxoutclk_i,
        gt8_rxoutclkfabric_out          =>      gt8_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt8_gtrxreset_in                =>      gt8_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt8_rxcharisk_out               =>      gt8_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt8_gthrxp_in                   =>      gt8_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt8_rxresetdone_out             =>      gt8_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt8_gttxreset_in                =>      gt8_gttxreset_i,
        gt8_txuserrdy_in                =>      gt8_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt8_txusrclk_in                 =>      gt8_txusrclk_in,
        gt8_txusrclk2_in                =>      gt8_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt8_txdlyen_in                  =>      gt8_txdlyen_i,
        gt8_txdlysreset_in              =>      gt8_txdlysreset_i,
        gt8_txdlysresetdone_out         =>      gt8_txdlysresetdone_i,
        gt8_txphalign_in                =>      gt8_txphalign_i,
        gt8_txphaligndone_out           =>      gt8_txphaligndone_i,
        gt8_txphalignen_in              =>      gt8_txphalignen_i,
        gt8_txphdlyreset_in             =>      gt8_txphdlyreset_i,
        gt8_txphinit_in                 =>      gt8_txphinit_i,
        gt8_txphinitdone_out            =>      gt8_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt8_txdata_in                   =>      gt8_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt8_gthtxn_out                  =>      gt8_gthtxn_out,
        gt8_gthtxp_out                  =>      gt8_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt8_txoutclk_out                =>      gt8_txoutclk_i,
        gt8_txoutclkfabric_out          =>      gt8_txoutclkfabric_out,
        gt8_txoutclkpcs_out             =>      gt8_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt8_txresetdone_out             =>      gt8_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt8_txcharisk_in                =>      gt8_txcharisk_in,


        GT9_DRP_BUSY_OUT                =>      GT9_DRP_BUSY_OUT,
        GT9_RXPMARESETDONE_OUT          =>      gt9_rxpmaresetdone_i,
        GT9_TXPMARESETDONE_OUT          =>      gt9_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT9  (X1Y13)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt9_drpaddr_in                  =>      gt9_drpaddr_in,
        gt9_drpclk_in                   =>      gt9_drpclk_in,
        gt9_drpdi_in                    =>      gt9_drpdi_in,
        gt9_drpdo_out                   =>      gt9_drpdo_out,
        gt9_drpen_in                    =>      gt9_drpen_in,
        gt9_drprdy_out                  =>      gt9_drprdy_out,
        gt9_drpwe_in                    =>      gt9_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt9_eyescanreset_in             =>      gt9_eyescanreset_in,
        gt9_rxuserrdy_in                =>      gt9_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt9_eyescandataerror_out        =>      gt9_eyescandataerror_out,
        gt9_eyescantrigger_in           =>      gt9_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt9_rxslide_in                  =>      gt9_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt9_dmonitorout_out             =>      gt9_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt9_rxusrclk_in                 =>      gt9_rxusrclk_in,
        gt9_rxusrclk2_in                =>      gt9_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt9_rxdata_out                  =>      gt9_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt9_rxdisperr_out               =>      gt9_rxdisperr_out,
        gt9_rxnotintable_out            =>      gt9_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt9_gthrxn_in                   =>      gt9_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt9_rxdlyen_in                  =>      gt9_rxdlyen_i,
        gt9_rxdlysreset_in              =>      gt9_rxdlysreset_i,
        gt9_rxdlysresetdone_out         =>      gt9_rxdlysresetdone_i,
        gt9_rxphalign_in                =>      gt9_rxphalign_i,
        gt9_rxphaligndone_out           =>      gt9_rxphaligndone_i,
        gt9_rxphalignen_in              =>      gt9_rxphalignen_i,
        gt9_rxphdlyreset_in             =>      gt9_rxphdlyreset_i,
        gt9_rxphmonitor_out             =>      gt9_rxphmonitor_out,
        gt9_rxphslipmonitor_out         =>      gt9_rxphslipmonitor_out,
        gt9_rxsyncallin_in              =>      gt9_rxsyncallin_i,
        gt9_rxsyncdone_out              =>      gt9_rxsyncdone_i,
        gt9_rxsyncin_in                 =>      gt9_rxsyncin_i,
        gt9_rxsyncmode_in               =>      gt9_rxsyncmode_i,
        gt9_rxsyncout_out               =>      gt9_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt9_rxbyteisaligned_out         =>      gt9_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt9_rxlpmhfhold_in              =>      gt9_rxlpmhfhold_i,
        gt9_rxlpmlfhold_in              =>      gt9_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt9_rxmonitorout_out            =>      gt9_rxmonitorout_out,
        gt9_rxmonitorsel_in             =>      gt9_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt9_rxoutclk_out                =>      gt9_rxoutclk_i,
        gt9_rxoutclkfabric_out          =>      gt9_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt9_gtrxreset_in                =>      gt9_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt9_rxcharisk_out               =>      gt9_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt9_gthrxp_in                   =>      gt9_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt9_rxresetdone_out             =>      gt9_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt9_gttxreset_in                =>      gt9_gttxreset_i,
        gt9_txuserrdy_in                =>      gt9_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt9_txusrclk_in                 =>      gt9_txusrclk_in,
        gt9_txusrclk2_in                =>      gt9_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt9_txdlyen_in                  =>      gt9_txdlyen_i,
        gt9_txdlysreset_in              =>      gt9_txdlysreset_i,
        gt9_txdlysresetdone_out         =>      gt9_txdlysresetdone_i,
        gt9_txphalign_in                =>      gt9_txphalign_i,
        gt9_txphaligndone_out           =>      gt9_txphaligndone_i,
        gt9_txphalignen_in              =>      gt9_txphalignen_i,
        gt9_txphdlyreset_in             =>      gt9_txphdlyreset_i,
        gt9_txphinit_in                 =>      gt9_txphinit_i,
        gt9_txphinitdone_out            =>      gt9_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt9_txdata_in                   =>      gt9_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt9_gthtxn_out                  =>      gt9_gthtxn_out,
        gt9_gthtxp_out                  =>      gt9_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt9_txoutclk_out                =>      gt9_txoutclk_i,
        gt9_txoutclkfabric_out          =>      gt9_txoutclkfabric_out,
        gt9_txoutclkpcs_out             =>      gt9_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt9_txresetdone_out             =>      gt9_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt9_txcharisk_in                =>      gt9_txcharisk_in,


        GT10_DRP_BUSY_OUT               =>      GT10_DRP_BUSY_OUT,
        GT10_RXPMARESETDONE_OUT         =>      gt10_rxpmaresetdone_i,
        GT10_TXPMARESETDONE_OUT         =>      gt10_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT10  (X1Y14)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt10_drpaddr_in                 =>      gt10_drpaddr_in,
        gt10_drpclk_in                  =>      gt10_drpclk_in,
        gt10_drpdi_in                   =>      gt10_drpdi_in,
        gt10_drpdo_out                  =>      gt10_drpdo_out,
        gt10_drpen_in                   =>      gt10_drpen_in,
        gt10_drprdy_out                 =>      gt10_drprdy_out,
        gt10_drpwe_in                   =>      gt10_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt10_eyescanreset_in            =>      gt10_eyescanreset_in,
        gt10_rxuserrdy_in               =>      gt10_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt10_eyescandataerror_out       =>      gt10_eyescandataerror_out,
        gt10_eyescantrigger_in          =>      gt10_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt10_rxslide_in                 =>      gt10_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt10_dmonitorout_out            =>      gt10_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt10_rxusrclk_in                =>      gt10_rxusrclk_in,
        gt10_rxusrclk2_in               =>      gt10_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt10_rxdata_out                 =>      gt10_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt10_rxdisperr_out              =>      gt10_rxdisperr_out,
        gt10_rxnotintable_out           =>      gt10_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt10_gthrxn_in                  =>      gt10_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt10_rxdlyen_in                 =>      gt10_rxdlyen_i,
        gt10_rxdlysreset_in             =>      gt10_rxdlysreset_i,
        gt10_rxdlysresetdone_out        =>      gt10_rxdlysresetdone_i,
        gt10_rxphalign_in               =>      gt10_rxphalign_i,
        gt10_rxphaligndone_out          =>      gt10_rxphaligndone_i,
        gt10_rxphalignen_in             =>      gt10_rxphalignen_i,
        gt10_rxphdlyreset_in            =>      gt10_rxphdlyreset_i,
        gt10_rxphmonitor_out            =>      gt10_rxphmonitor_out,
        gt10_rxphslipmonitor_out        =>      gt10_rxphslipmonitor_out,
        gt10_rxsyncallin_in             =>      gt10_rxsyncallin_i,
        gt10_rxsyncdone_out             =>      gt10_rxsyncdone_i,
        gt10_rxsyncin_in                =>      gt10_rxsyncin_i,
        gt10_rxsyncmode_in              =>      gt10_rxsyncmode_i,
        gt10_rxsyncout_out              =>      gt10_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt10_rxbyteisaligned_out        =>      gt10_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt10_rxlpmhfhold_in             =>      gt10_rxlpmhfhold_i,
        gt10_rxlpmlfhold_in             =>      gt10_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt10_rxmonitorout_out           =>      gt10_rxmonitorout_out,
        gt10_rxmonitorsel_in            =>      gt10_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt10_rxoutclk_out               =>      gt10_rxoutclk_i,
        gt10_rxoutclkfabric_out         =>      gt10_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt10_gtrxreset_in               =>      gt10_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt10_rxcharisk_out              =>      gt10_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt10_gthrxp_in                  =>      gt10_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt10_rxresetdone_out            =>      gt10_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt10_gttxreset_in               =>      gt10_gttxreset_i,
        gt10_txuserrdy_in               =>      gt10_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt10_txusrclk_in                =>      gt10_txusrclk_in,
        gt10_txusrclk2_in               =>      gt10_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt10_txdlyen_in                 =>      gt10_txdlyen_i,
        gt10_txdlysreset_in             =>      gt10_txdlysreset_i,
        gt10_txdlysresetdone_out        =>      gt10_txdlysresetdone_i,
        gt10_txphalign_in               =>      gt10_txphalign_i,
        gt10_txphaligndone_out          =>      gt10_txphaligndone_i,
        gt10_txphalignen_in             =>      gt10_txphalignen_i,
        gt10_txphdlyreset_in            =>      gt10_txphdlyreset_i,
        gt10_txphinit_in                =>      gt10_txphinit_i,
        gt10_txphinitdone_out           =>      gt10_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt10_txdata_in                  =>      gt10_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt10_gthtxn_out                 =>      gt10_gthtxn_out,
        gt10_gthtxp_out                 =>      gt10_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt10_txoutclk_out               =>      gt10_txoutclk_i,
        gt10_txoutclkfabric_out         =>      gt10_txoutclkfabric_out,
        gt10_txoutclkpcs_out            =>      gt10_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt10_txresetdone_out            =>      gt10_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt10_txcharisk_in               =>      gt10_txcharisk_in,


        GT11_DRP_BUSY_OUT               =>      GT11_DRP_BUSY_OUT,
        GT11_RXPMARESETDONE_OUT         =>      gt11_rxpmaresetdone_i,
        GT11_TXPMARESETDONE_OUT         =>      gt11_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT11  (X1Y15)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt11_drpaddr_in                 =>      gt11_drpaddr_in,
        gt11_drpclk_in                  =>      gt11_drpclk_in,
        gt11_drpdi_in                   =>      gt11_drpdi_in,
        gt11_drpdo_out                  =>      gt11_drpdo_out,
        gt11_drpen_in                   =>      gt11_drpen_in,
        gt11_drprdy_out                 =>      gt11_drprdy_out,
        gt11_drpwe_in                   =>      gt11_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt11_eyescanreset_in            =>      gt11_eyescanreset_in,
        gt11_rxuserrdy_in               =>      gt11_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt11_eyescandataerror_out       =>      gt11_eyescandataerror_out,
        gt11_eyescantrigger_in          =>      gt11_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt11_rxslide_in                 =>      gt11_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt11_dmonitorout_out            =>      gt11_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt11_rxusrclk_in                =>      gt11_rxusrclk_in,
        gt11_rxusrclk2_in               =>      gt11_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt11_rxdata_out                 =>      gt11_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt11_rxdisperr_out              =>      gt11_rxdisperr_out,
        gt11_rxnotintable_out           =>      gt11_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt11_gthrxn_in                  =>      gt11_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt11_rxdlyen_in                 =>      gt11_rxdlyen_i,
        gt11_rxdlysreset_in             =>      gt11_rxdlysreset_i,
        gt11_rxdlysresetdone_out        =>      gt11_rxdlysresetdone_i,
        gt11_rxphalign_in               =>      gt11_rxphalign_i,
        gt11_rxphaligndone_out          =>      gt11_rxphaligndone_i,
        gt11_rxphalignen_in             =>      gt11_rxphalignen_i,
        gt11_rxphdlyreset_in            =>      gt11_rxphdlyreset_i,
        gt11_rxphmonitor_out            =>      gt11_rxphmonitor_out,
        gt11_rxphslipmonitor_out        =>      gt11_rxphslipmonitor_out,
        gt11_rxsyncallin_in             =>      gt11_rxsyncallin_i,
        gt11_rxsyncdone_out             =>      gt11_rxsyncdone_i,
        gt11_rxsyncin_in                =>      gt11_rxsyncin_i,
        gt11_rxsyncmode_in              =>      gt11_rxsyncmode_i,
        gt11_rxsyncout_out              =>      gt11_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt11_rxbyteisaligned_out        =>      gt11_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt11_rxlpmhfhold_in             =>      gt11_rxlpmhfhold_i,
        gt11_rxlpmlfhold_in             =>      gt11_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt11_rxmonitorout_out           =>      gt11_rxmonitorout_out,
        gt11_rxmonitorsel_in            =>      gt11_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt11_rxoutclk_out               =>      gt11_rxoutclk_i,
        gt11_rxoutclkfabric_out         =>      gt11_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt11_gtrxreset_in               =>      gt11_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt11_rxcharisk_out              =>      gt11_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt11_gthrxp_in                  =>      gt11_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt11_rxresetdone_out            =>      gt11_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt11_gttxreset_in               =>      gt11_gttxreset_i,
        gt11_txuserrdy_in               =>      gt11_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt11_txusrclk_in                =>      gt11_txusrclk_in,
        gt11_txusrclk2_in               =>      gt11_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt11_txdlyen_in                 =>      gt11_txdlyen_i,
        gt11_txdlysreset_in             =>      gt11_txdlysreset_i,
        gt11_txdlysresetdone_out        =>      gt11_txdlysresetdone_i,
        gt11_txphalign_in               =>      gt11_txphalign_i,
        gt11_txphaligndone_out          =>      gt11_txphaligndone_i,
        gt11_txphalignen_in             =>      gt11_txphalignen_i,
        gt11_txphdlyreset_in            =>      gt11_txphdlyreset_i,
        gt11_txphinit_in                =>      gt11_txphinit_i,
        gt11_txphinitdone_out           =>      gt11_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt11_txdata_in                  =>      gt11_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt11_gthtxn_out                 =>      gt11_gthtxn_out,
        gt11_gthtxp_out                 =>      gt11_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt11_txoutclk_out               =>      gt11_txoutclk_i,
        gt11_txoutclkfabric_out         =>      gt11_txoutclkfabric_out,
        gt11_txoutclkpcs_out            =>      gt11_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt11_txresetdone_out            =>      gt11_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt11_txcharisk_in               =>      gt11_txcharisk_in,


        GT12_DRP_BUSY_OUT               =>      GT12_DRP_BUSY_OUT,
        GT12_RXPMARESETDONE_OUT         =>      gt12_rxpmaresetdone_i,
        GT12_TXPMARESETDONE_OUT         =>      gt12_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT12  (X1Y16)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt12_drpaddr_in                 =>      gt12_drpaddr_in,
        gt12_drpclk_in                  =>      gt12_drpclk_in,
        gt12_drpdi_in                   =>      gt12_drpdi_in,
        gt12_drpdo_out                  =>      gt12_drpdo_out,
        gt12_drpen_in                   =>      gt12_drpen_in,
        gt12_drprdy_out                 =>      gt12_drprdy_out,
        gt12_drpwe_in                   =>      gt12_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt12_eyescanreset_in            =>      gt12_eyescanreset_in,
        gt12_rxuserrdy_in               =>      gt12_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt12_eyescandataerror_out       =>      gt12_eyescandataerror_out,
        gt12_eyescantrigger_in          =>      gt12_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt12_rxslide_in                 =>      gt12_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt12_dmonitorout_out            =>      gt12_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt12_rxusrclk_in                =>      gt12_rxusrclk_in,
        gt12_rxusrclk2_in               =>      gt12_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt12_rxdata_out                 =>      gt12_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt12_rxdisperr_out              =>      gt12_rxdisperr_out,
        gt12_rxnotintable_out           =>      gt12_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt12_gthrxn_in                  =>      gt12_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt12_rxdlyen_in                 =>      gt12_rxdlyen_i,
        gt12_rxdlysreset_in             =>      gt12_rxdlysreset_i,
        gt12_rxdlysresetdone_out        =>      gt12_rxdlysresetdone_i,
        gt12_rxphalign_in               =>      gt12_rxphalign_i,
        gt12_rxphaligndone_out          =>      gt12_rxphaligndone_i,
        gt12_rxphalignen_in             =>      gt12_rxphalignen_i,
        gt12_rxphdlyreset_in            =>      gt12_rxphdlyreset_i,
        gt12_rxphmonitor_out            =>      gt12_rxphmonitor_out,
        gt12_rxphslipmonitor_out        =>      gt12_rxphslipmonitor_out,
        gt12_rxsyncallin_in             =>      gt12_rxsyncallin_i,
        gt12_rxsyncdone_out             =>      gt12_rxsyncdone_i,
        gt12_rxsyncin_in                =>      gt12_rxsyncin_i,
        gt12_rxsyncmode_in              =>      gt12_rxsyncmode_i,
        gt12_rxsyncout_out              =>      gt12_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt12_rxbyteisaligned_out        =>      gt12_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt12_rxlpmhfhold_in             =>      gt12_rxlpmhfhold_i,
        gt12_rxlpmlfhold_in             =>      gt12_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt12_rxmonitorout_out           =>      gt12_rxmonitorout_out,
        gt12_rxmonitorsel_in            =>      gt12_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt12_rxoutclk_out               =>      gt12_rxoutclk_i,
        gt12_rxoutclkfabric_out         =>      gt12_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt12_gtrxreset_in               =>      gt12_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt12_rxcharisk_out              =>      gt12_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt12_gthrxp_in                  =>      gt12_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt12_rxresetdone_out            =>      gt12_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt12_gttxreset_in               =>      gt12_gttxreset_i,
        gt12_txuserrdy_in               =>      gt12_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt12_txusrclk_in                =>      gt12_txusrclk_in,
        gt12_txusrclk2_in               =>      gt12_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt12_txdlyen_in                 =>      gt12_txdlyen_i,
        gt12_txdlysreset_in             =>      gt12_txdlysreset_i,
        gt12_txdlysresetdone_out        =>      gt12_txdlysresetdone_i,
        gt12_txphalign_in               =>      gt12_txphalign_i,
        gt12_txphaligndone_out          =>      gt12_txphaligndone_i,
        gt12_txphalignen_in             =>      gt12_txphalignen_i,
        gt12_txphdlyreset_in            =>      gt12_txphdlyreset_i,
        gt12_txphinit_in                =>      gt12_txphinit_i,
        gt12_txphinitdone_out           =>      gt12_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt12_txdata_in                  =>      gt12_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt12_gthtxn_out                 =>      gt12_gthtxn_out,
        gt12_gthtxp_out                 =>      gt12_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt12_txoutclk_out               =>      gt12_txoutclk_i,
        gt12_txoutclkfabric_out         =>      gt12_txoutclkfabric_out,
        gt12_txoutclkpcs_out            =>      gt12_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt12_txresetdone_out            =>      gt12_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt12_txcharisk_in               =>      gt12_txcharisk_in,


        GT13_DRP_BUSY_OUT               =>      GT13_DRP_BUSY_OUT,
        GT13_RXPMARESETDONE_OUT         =>      gt13_rxpmaresetdone_i,
        GT13_TXPMARESETDONE_OUT         =>      gt13_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT13  (X1Y17)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt13_drpaddr_in                 =>      gt13_drpaddr_in,
        gt13_drpclk_in                  =>      gt13_drpclk_in,
        gt13_drpdi_in                   =>      gt13_drpdi_in,
        gt13_drpdo_out                  =>      gt13_drpdo_out,
        gt13_drpen_in                   =>      gt13_drpen_in,
        gt13_drprdy_out                 =>      gt13_drprdy_out,
        gt13_drpwe_in                   =>      gt13_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt13_eyescanreset_in            =>      gt13_eyescanreset_in,
        gt13_rxuserrdy_in               =>      gt13_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt13_eyescandataerror_out       =>      gt13_eyescandataerror_out,
        gt13_eyescantrigger_in          =>      gt13_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt13_rxslide_in                 =>      gt13_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt13_dmonitorout_out            =>      gt13_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt13_rxusrclk_in                =>      gt13_rxusrclk_in,
        gt13_rxusrclk2_in               =>      gt13_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt13_rxdata_out                 =>      gt13_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt13_rxdisperr_out              =>      gt13_rxdisperr_out,
        gt13_rxnotintable_out           =>      gt13_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt13_gthrxn_in                  =>      gt13_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt13_rxdlyen_in                 =>      gt13_rxdlyen_i,
        gt13_rxdlysreset_in             =>      gt13_rxdlysreset_i,
        gt13_rxdlysresetdone_out        =>      gt13_rxdlysresetdone_i,
        gt13_rxphalign_in               =>      gt13_rxphalign_i,
        gt13_rxphaligndone_out          =>      gt13_rxphaligndone_i,
        gt13_rxphalignen_in             =>      gt13_rxphalignen_i,
        gt13_rxphdlyreset_in            =>      gt13_rxphdlyreset_i,
        gt13_rxphmonitor_out            =>      gt13_rxphmonitor_out,
        gt13_rxphslipmonitor_out        =>      gt13_rxphslipmonitor_out,
        gt13_rxsyncallin_in             =>      gt13_rxsyncallin_i,
        gt13_rxsyncdone_out             =>      gt13_rxsyncdone_i,
        gt13_rxsyncin_in                =>      gt13_rxsyncin_i,
        gt13_rxsyncmode_in              =>      gt13_rxsyncmode_i,
        gt13_rxsyncout_out              =>      gt13_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt13_rxbyteisaligned_out        =>      gt13_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt13_rxlpmhfhold_in             =>      gt13_rxlpmhfhold_i,
        gt13_rxlpmlfhold_in             =>      gt13_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt13_rxmonitorout_out           =>      gt13_rxmonitorout_out,
        gt13_rxmonitorsel_in            =>      gt13_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt13_rxoutclk_out               =>      gt13_rxoutclk_i,
        gt13_rxoutclkfabric_out         =>      gt13_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt13_gtrxreset_in               =>      gt13_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt13_rxcharisk_out              =>      gt13_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt13_gthrxp_in                  =>      gt13_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt13_rxresetdone_out            =>      gt13_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt13_gttxreset_in               =>      gt13_gttxreset_i,
        gt13_txuserrdy_in               =>      gt13_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt13_txusrclk_in                =>      gt13_txusrclk_in,
        gt13_txusrclk2_in               =>      gt13_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt13_txdlyen_in                 =>      gt13_txdlyen_i,
        gt13_txdlysreset_in             =>      gt13_txdlysreset_i,
        gt13_txdlysresetdone_out        =>      gt13_txdlysresetdone_i,
        gt13_txphalign_in               =>      gt13_txphalign_i,
        gt13_txphaligndone_out          =>      gt13_txphaligndone_i,
        gt13_txphalignen_in             =>      gt13_txphalignen_i,
        gt13_txphdlyreset_in            =>      gt13_txphdlyreset_i,
        gt13_txphinit_in                =>      gt13_txphinit_i,
        gt13_txphinitdone_out           =>      gt13_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt13_txdata_in                  =>      gt13_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt13_gthtxn_out                 =>      gt13_gthtxn_out,
        gt13_gthtxp_out                 =>      gt13_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt13_txoutclk_out               =>      gt13_txoutclk_i,
        gt13_txoutclkfabric_out         =>      gt13_txoutclkfabric_out,
        gt13_txoutclkpcs_out            =>      gt13_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt13_txresetdone_out            =>      gt13_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt13_txcharisk_in               =>      gt13_txcharisk_in,


        GT14_DRP_BUSY_OUT               =>      GT14_DRP_BUSY_OUT,
        GT14_RXPMARESETDONE_OUT         =>      gt14_rxpmaresetdone_i,
        GT14_TXPMARESETDONE_OUT         =>      gt14_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT14  (X1Y18)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt14_drpaddr_in                 =>      gt14_drpaddr_in,
        gt14_drpclk_in                  =>      gt14_drpclk_in,
        gt14_drpdi_in                   =>      gt14_drpdi_in,
        gt14_drpdo_out                  =>      gt14_drpdo_out,
        gt14_drpen_in                   =>      gt14_drpen_in,
        gt14_drprdy_out                 =>      gt14_drprdy_out,
        gt14_drpwe_in                   =>      gt14_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt14_eyescanreset_in            =>      gt14_eyescanreset_in,
        gt14_rxuserrdy_in               =>      gt14_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt14_eyescandataerror_out       =>      gt14_eyescandataerror_out,
        gt14_eyescantrigger_in          =>      gt14_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt14_rxslide_in                 =>      gt14_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt14_dmonitorout_out            =>      gt14_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt14_rxusrclk_in                =>      gt14_rxusrclk_in,
        gt14_rxusrclk2_in               =>      gt14_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt14_rxdata_out                 =>      gt14_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt14_rxdisperr_out              =>      gt14_rxdisperr_out,
        gt14_rxnotintable_out           =>      gt14_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt14_gthrxn_in                  =>      gt14_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt14_rxdlyen_in                 =>      gt14_rxdlyen_i,
        gt14_rxdlysreset_in             =>      gt14_rxdlysreset_i,
        gt14_rxdlysresetdone_out        =>      gt14_rxdlysresetdone_i,
        gt14_rxphalign_in               =>      gt14_rxphalign_i,
        gt14_rxphaligndone_out          =>      gt14_rxphaligndone_i,
        gt14_rxphalignen_in             =>      gt14_rxphalignen_i,
        gt14_rxphdlyreset_in            =>      gt14_rxphdlyreset_i,
        gt14_rxphmonitor_out            =>      gt14_rxphmonitor_out,
        gt14_rxphslipmonitor_out        =>      gt14_rxphslipmonitor_out,
        gt14_rxsyncallin_in             =>      gt14_rxsyncallin_i,
        gt14_rxsyncdone_out             =>      gt14_rxsyncdone_i,
        gt14_rxsyncin_in                =>      gt14_rxsyncin_i,
        gt14_rxsyncmode_in              =>      gt14_rxsyncmode_i,
        gt14_rxsyncout_out              =>      gt14_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt14_rxbyteisaligned_out        =>      gt14_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt14_rxlpmhfhold_in             =>      gt14_rxlpmhfhold_i,
        gt14_rxlpmlfhold_in             =>      gt14_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt14_rxmonitorout_out           =>      gt14_rxmonitorout_out,
        gt14_rxmonitorsel_in            =>      gt14_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt14_rxoutclk_out               =>      gt14_rxoutclk_i,
        gt14_rxoutclkfabric_out         =>      gt14_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt14_gtrxreset_in               =>      gt14_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt14_rxcharisk_out              =>      gt14_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt14_gthrxp_in                  =>      gt14_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt14_rxresetdone_out            =>      gt14_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt14_gttxreset_in               =>      gt14_gttxreset_i,
        gt14_txuserrdy_in               =>      gt14_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt14_txusrclk_in                =>      gt14_txusrclk_in,
        gt14_txusrclk2_in               =>      gt14_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt14_txdlyen_in                 =>      gt14_txdlyen_i,
        gt14_txdlysreset_in             =>      gt14_txdlysreset_i,
        gt14_txdlysresetdone_out        =>      gt14_txdlysresetdone_i,
        gt14_txphalign_in               =>      gt14_txphalign_i,
        gt14_txphaligndone_out          =>      gt14_txphaligndone_i,
        gt14_txphalignen_in             =>      gt14_txphalignen_i,
        gt14_txphdlyreset_in            =>      gt14_txphdlyreset_i,
        gt14_txphinit_in                =>      gt14_txphinit_i,
        gt14_txphinitdone_out           =>      gt14_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt14_txdata_in                  =>      gt14_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt14_gthtxn_out                 =>      gt14_gthtxn_out,
        gt14_gthtxp_out                 =>      gt14_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt14_txoutclk_out               =>      gt14_txoutclk_i,
        gt14_txoutclkfabric_out         =>      gt14_txoutclkfabric_out,
        gt14_txoutclkpcs_out            =>      gt14_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt14_txresetdone_out            =>      gt14_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt14_txcharisk_in               =>      gt14_txcharisk_in,


        GT15_DRP_BUSY_OUT               =>      GT15_DRP_BUSY_OUT,
        GT15_RXPMARESETDONE_OUT         =>      gt15_rxpmaresetdone_i,
        GT15_TXPMARESETDONE_OUT         =>      gt15_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT15  (X1Y19)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt15_drpaddr_in                 =>      gt15_drpaddr_in,
        gt15_drpclk_in                  =>      gt15_drpclk_in,
        gt15_drpdi_in                   =>      gt15_drpdi_in,
        gt15_drpdo_out                  =>      gt15_drpdo_out,
        gt15_drpen_in                   =>      gt15_drpen_in,
        gt15_drprdy_out                 =>      gt15_drprdy_out,
        gt15_drpwe_in                   =>      gt15_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt15_eyescanreset_in            =>      gt15_eyescanreset_in,
        gt15_rxuserrdy_in               =>      gt15_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt15_eyescandataerror_out       =>      gt15_eyescandataerror_out,
        gt15_eyescantrigger_in          =>      gt15_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt15_rxslide_in                 =>      gt15_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt15_dmonitorout_out            =>      gt15_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt15_rxusrclk_in                =>      gt15_rxusrclk_in,
        gt15_rxusrclk2_in               =>      gt15_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt15_rxdata_out                 =>      gt15_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt15_rxdisperr_out              =>      gt15_rxdisperr_out,
        gt15_rxnotintable_out           =>      gt15_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt15_gthrxn_in                  =>      gt15_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt15_rxdlyen_in                 =>      gt15_rxdlyen_i,
        gt15_rxdlysreset_in             =>      gt15_rxdlysreset_i,
        gt15_rxdlysresetdone_out        =>      gt15_rxdlysresetdone_i,
        gt15_rxphalign_in               =>      gt15_rxphalign_i,
        gt15_rxphaligndone_out          =>      gt15_rxphaligndone_i,
        gt15_rxphalignen_in             =>      gt15_rxphalignen_i,
        gt15_rxphdlyreset_in            =>      gt15_rxphdlyreset_i,
        gt15_rxphmonitor_out            =>      gt15_rxphmonitor_out,
        gt15_rxphslipmonitor_out        =>      gt15_rxphslipmonitor_out,
        gt15_rxsyncallin_in             =>      gt15_rxsyncallin_i,
        gt15_rxsyncdone_out             =>      gt15_rxsyncdone_i,
        gt15_rxsyncin_in                =>      gt15_rxsyncin_i,
        gt15_rxsyncmode_in              =>      gt15_rxsyncmode_i,
        gt15_rxsyncout_out              =>      gt15_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt15_rxbyteisaligned_out        =>      gt15_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt15_rxlpmhfhold_in             =>      gt15_rxlpmhfhold_i,
        gt15_rxlpmlfhold_in             =>      gt15_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt15_rxmonitorout_out           =>      gt15_rxmonitorout_out,
        gt15_rxmonitorsel_in            =>      gt15_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt15_rxoutclk_out               =>      gt15_rxoutclk_i,
        gt15_rxoutclkfabric_out         =>      gt15_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt15_gtrxreset_in               =>      gt15_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt15_rxcharisk_out              =>      gt15_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt15_gthrxp_in                  =>      gt15_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt15_rxresetdone_out            =>      gt15_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt15_gttxreset_in               =>      gt15_gttxreset_i,
        gt15_txuserrdy_in               =>      gt15_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt15_txusrclk_in                =>      gt15_txusrclk_in,
        gt15_txusrclk2_in               =>      gt15_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt15_txdlyen_in                 =>      gt15_txdlyen_i,
        gt15_txdlysreset_in             =>      gt15_txdlysreset_i,
        gt15_txdlysresetdone_out        =>      gt15_txdlysresetdone_i,
        gt15_txphalign_in               =>      gt15_txphalign_i,
        gt15_txphaligndone_out          =>      gt15_txphaligndone_i,
        gt15_txphalignen_in             =>      gt15_txphalignen_i,
        gt15_txphdlyreset_in            =>      gt15_txphdlyreset_i,
        gt15_txphinit_in                =>      gt15_txphinit_i,
        gt15_txphinitdone_out           =>      gt15_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt15_txdata_in                  =>      gt15_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt15_gthtxn_out                 =>      gt15_gthtxn_out,
        gt15_gthtxp_out                 =>      gt15_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt15_txoutclk_out               =>      gt15_txoutclk_i,
        gt15_txoutclkfabric_out         =>      gt15_txoutclkfabric_out,
        gt15_txoutclkpcs_out            =>      gt15_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt15_txresetdone_out            =>      gt15_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt15_txcharisk_in               =>      gt15_txcharisk_in,


        GT16_DRP_BUSY_OUT               =>      GT16_DRP_BUSY_OUT,
        GT16_RXPMARESETDONE_OUT         =>      gt16_rxpmaresetdone_i,
        GT16_TXPMARESETDONE_OUT         =>      gt16_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT16  (X1Y20)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt16_drpaddr_in                 =>      gt16_drpaddr_in,
        gt16_drpclk_in                  =>      gt16_drpclk_in,
        gt16_drpdi_in                   =>      gt16_drpdi_in,
        gt16_drpdo_out                  =>      gt16_drpdo_out,
        gt16_drpen_in                   =>      gt16_drpen_in,
        gt16_drprdy_out                 =>      gt16_drprdy_out,
        gt16_drpwe_in                   =>      gt16_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt16_eyescanreset_in            =>      gt16_eyescanreset_in,
        gt16_rxuserrdy_in               =>      gt16_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt16_eyescandataerror_out       =>      gt16_eyescandataerror_out,
        gt16_eyescantrigger_in          =>      gt16_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt16_rxslide_in                 =>      gt16_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt16_dmonitorout_out            =>      gt16_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt16_rxusrclk_in                =>      gt16_rxusrclk_in,
        gt16_rxusrclk2_in               =>      gt16_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt16_rxdata_out                 =>      gt16_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt16_rxdisperr_out              =>      gt16_rxdisperr_out,
        gt16_rxnotintable_out           =>      gt16_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt16_gthrxn_in                  =>      gt16_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt16_rxdlyen_in                 =>      gt16_rxdlyen_i,
        gt16_rxdlysreset_in             =>      gt16_rxdlysreset_i,
        gt16_rxdlysresetdone_out        =>      gt16_rxdlysresetdone_i,
        gt16_rxphalign_in               =>      gt16_rxphalign_i,
        gt16_rxphaligndone_out          =>      gt16_rxphaligndone_i,
        gt16_rxphalignen_in             =>      gt16_rxphalignen_i,
        gt16_rxphdlyreset_in            =>      gt16_rxphdlyreset_i,
        gt16_rxphmonitor_out            =>      gt16_rxphmonitor_out,
        gt16_rxphslipmonitor_out        =>      gt16_rxphslipmonitor_out,
        gt16_rxsyncallin_in             =>      gt16_rxsyncallin_i,
        gt16_rxsyncdone_out             =>      gt16_rxsyncdone_i,
        gt16_rxsyncin_in                =>      gt16_rxsyncin_i,
        gt16_rxsyncmode_in              =>      gt16_rxsyncmode_i,
        gt16_rxsyncout_out              =>      gt16_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt16_rxbyteisaligned_out        =>      gt16_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt16_rxlpmhfhold_in             =>      gt16_rxlpmhfhold_i,
        gt16_rxlpmlfhold_in             =>      gt16_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt16_rxmonitorout_out           =>      gt16_rxmonitorout_out,
        gt16_rxmonitorsel_in            =>      gt16_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt16_rxoutclk_out               =>      gt16_rxoutclk_i,
        gt16_rxoutclkfabric_out         =>      gt16_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt16_gtrxreset_in               =>      gt16_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt16_rxcharisk_out              =>      gt16_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt16_gthrxp_in                  =>      gt16_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt16_rxresetdone_out            =>      gt16_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt16_gttxreset_in               =>      gt16_gttxreset_i,
        gt16_txuserrdy_in               =>      gt16_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt16_txusrclk_in                =>      gt16_txusrclk_in,
        gt16_txusrclk2_in               =>      gt16_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt16_txdlyen_in                 =>      gt16_txdlyen_i,
        gt16_txdlysreset_in             =>      gt16_txdlysreset_i,
        gt16_txdlysresetdone_out        =>      gt16_txdlysresetdone_i,
        gt16_txphalign_in               =>      gt16_txphalign_i,
        gt16_txphaligndone_out          =>      gt16_txphaligndone_i,
        gt16_txphalignen_in             =>      gt16_txphalignen_i,
        gt16_txphdlyreset_in            =>      gt16_txphdlyreset_i,
        gt16_txphinit_in                =>      gt16_txphinit_i,
        gt16_txphinitdone_out           =>      gt16_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt16_txdata_in                  =>      gt16_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt16_gthtxn_out                 =>      gt16_gthtxn_out,
        gt16_gthtxp_out                 =>      gt16_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt16_txoutclk_out               =>      gt16_txoutclk_i,
        gt16_txoutclkfabric_out         =>      gt16_txoutclkfabric_out,
        gt16_txoutclkpcs_out            =>      gt16_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt16_txresetdone_out            =>      gt16_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt16_txcharisk_in               =>      gt16_txcharisk_in,


        GT17_DRP_BUSY_OUT               =>      GT17_DRP_BUSY_OUT,
        GT17_RXPMARESETDONE_OUT         =>      gt17_rxpmaresetdone_i,
        GT17_TXPMARESETDONE_OUT         =>      gt17_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT17  (X1Y21)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt17_drpaddr_in                 =>      gt17_drpaddr_in,
        gt17_drpclk_in                  =>      gt17_drpclk_in,
        gt17_drpdi_in                   =>      gt17_drpdi_in,
        gt17_drpdo_out                  =>      gt17_drpdo_out,
        gt17_drpen_in                   =>      gt17_drpen_in,
        gt17_drprdy_out                 =>      gt17_drprdy_out,
        gt17_drpwe_in                   =>      gt17_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt17_eyescanreset_in            =>      gt17_eyescanreset_in,
        gt17_rxuserrdy_in               =>      gt17_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt17_eyescandataerror_out       =>      gt17_eyescandataerror_out,
        gt17_eyescantrigger_in          =>      gt17_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt17_rxslide_in                 =>      gt17_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt17_dmonitorout_out            =>      gt17_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt17_rxusrclk_in                =>      gt17_rxusrclk_in,
        gt17_rxusrclk2_in               =>      gt17_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt17_rxdata_out                 =>      gt17_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt17_rxdisperr_out              =>      gt17_rxdisperr_out,
        gt17_rxnotintable_out           =>      gt17_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt17_gthrxn_in                  =>      gt17_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt17_rxdlyen_in                 =>      gt17_rxdlyen_i,
        gt17_rxdlysreset_in             =>      gt17_rxdlysreset_i,
        gt17_rxdlysresetdone_out        =>      gt17_rxdlysresetdone_i,
        gt17_rxphalign_in               =>      gt17_rxphalign_i,
        gt17_rxphaligndone_out          =>      gt17_rxphaligndone_i,
        gt17_rxphalignen_in             =>      gt17_rxphalignen_i,
        gt17_rxphdlyreset_in            =>      gt17_rxphdlyreset_i,
        gt17_rxphmonitor_out            =>      gt17_rxphmonitor_out,
        gt17_rxphslipmonitor_out        =>      gt17_rxphslipmonitor_out,
        gt17_rxsyncallin_in             =>      gt17_rxsyncallin_i,
        gt17_rxsyncdone_out             =>      gt17_rxsyncdone_i,
        gt17_rxsyncin_in                =>      gt17_rxsyncin_i,
        gt17_rxsyncmode_in              =>      gt17_rxsyncmode_i,
        gt17_rxsyncout_out              =>      gt17_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt17_rxbyteisaligned_out        =>      gt17_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt17_rxlpmhfhold_in             =>      gt17_rxlpmhfhold_i,
        gt17_rxlpmlfhold_in             =>      gt17_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt17_rxmonitorout_out           =>      gt17_rxmonitorout_out,
        gt17_rxmonitorsel_in            =>      gt17_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt17_rxoutclk_out               =>      gt17_rxoutclk_i,
        gt17_rxoutclkfabric_out         =>      gt17_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt17_gtrxreset_in               =>      gt17_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt17_rxcharisk_out              =>      gt17_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt17_gthrxp_in                  =>      gt17_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt17_rxresetdone_out            =>      gt17_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt17_gttxreset_in               =>      gt17_gttxreset_i,
        gt17_txuserrdy_in               =>      gt17_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt17_txusrclk_in                =>      gt17_txusrclk_in,
        gt17_txusrclk2_in               =>      gt17_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt17_txdlyen_in                 =>      gt17_txdlyen_i,
        gt17_txdlysreset_in             =>      gt17_txdlysreset_i,
        gt17_txdlysresetdone_out        =>      gt17_txdlysresetdone_i,
        gt17_txphalign_in               =>      gt17_txphalign_i,
        gt17_txphaligndone_out          =>      gt17_txphaligndone_i,
        gt17_txphalignen_in             =>      gt17_txphalignen_i,
        gt17_txphdlyreset_in            =>      gt17_txphdlyreset_i,
        gt17_txphinit_in                =>      gt17_txphinit_i,
        gt17_txphinitdone_out           =>      gt17_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt17_txdata_in                  =>      gt17_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt17_gthtxn_out                 =>      gt17_gthtxn_out,
        gt17_gthtxp_out                 =>      gt17_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt17_txoutclk_out               =>      gt17_txoutclk_i,
        gt17_txoutclkfabric_out         =>      gt17_txoutclkfabric_out,
        gt17_txoutclkpcs_out            =>      gt17_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt17_txresetdone_out            =>      gt17_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt17_txcharisk_in               =>      gt17_txcharisk_in,


        GT18_DRP_BUSY_OUT               =>      GT18_DRP_BUSY_OUT,
        GT18_RXPMARESETDONE_OUT         =>      gt18_rxpmaresetdone_i,
        GT18_TXPMARESETDONE_OUT         =>      gt18_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT18  (X1Y22)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt18_drpaddr_in                 =>      gt18_drpaddr_in,
        gt18_drpclk_in                  =>      gt18_drpclk_in,
        gt18_drpdi_in                   =>      gt18_drpdi_in,
        gt18_drpdo_out                  =>      gt18_drpdo_out,
        gt18_drpen_in                   =>      gt18_drpen_in,
        gt18_drprdy_out                 =>      gt18_drprdy_out,
        gt18_drpwe_in                   =>      gt18_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt18_eyescanreset_in            =>      gt18_eyescanreset_in,
        gt18_rxuserrdy_in               =>      gt18_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt18_eyescandataerror_out       =>      gt18_eyescandataerror_out,
        gt18_eyescantrigger_in          =>      gt18_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt18_rxslide_in                 =>      gt18_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt18_dmonitorout_out            =>      gt18_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt18_rxusrclk_in                =>      gt18_rxusrclk_in,
        gt18_rxusrclk2_in               =>      gt18_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt18_rxdata_out                 =>      gt18_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt18_rxdisperr_out              =>      gt18_rxdisperr_out,
        gt18_rxnotintable_out           =>      gt18_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt18_gthrxn_in                  =>      gt18_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt18_rxdlyen_in                 =>      gt18_rxdlyen_i,
        gt18_rxdlysreset_in             =>      gt18_rxdlysreset_i,
        gt18_rxdlysresetdone_out        =>      gt18_rxdlysresetdone_i,
        gt18_rxphalign_in               =>      gt18_rxphalign_i,
        gt18_rxphaligndone_out          =>      gt18_rxphaligndone_i,
        gt18_rxphalignen_in             =>      gt18_rxphalignen_i,
        gt18_rxphdlyreset_in            =>      gt18_rxphdlyreset_i,
        gt18_rxphmonitor_out            =>      gt18_rxphmonitor_out,
        gt18_rxphslipmonitor_out        =>      gt18_rxphslipmonitor_out,
        gt18_rxsyncallin_in             =>      gt18_rxsyncallin_i,
        gt18_rxsyncdone_out             =>      gt18_rxsyncdone_i,
        gt18_rxsyncin_in                =>      gt18_rxsyncin_i,
        gt18_rxsyncmode_in              =>      gt18_rxsyncmode_i,
        gt18_rxsyncout_out              =>      gt18_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt18_rxbyteisaligned_out        =>      gt18_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt18_rxlpmhfhold_in             =>      gt18_rxlpmhfhold_i,
        gt18_rxlpmlfhold_in             =>      gt18_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt18_rxmonitorout_out           =>      gt18_rxmonitorout_out,
        gt18_rxmonitorsel_in            =>      gt18_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt18_rxoutclk_out               =>      gt18_rxoutclk_i,
        gt18_rxoutclkfabric_out         =>      gt18_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt18_gtrxreset_in               =>      gt18_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt18_rxcharisk_out              =>      gt18_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt18_gthrxp_in                  =>      gt18_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt18_rxresetdone_out            =>      gt18_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt18_gttxreset_in               =>      gt18_gttxreset_i,
        gt18_txuserrdy_in               =>      gt18_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt18_txusrclk_in                =>      gt18_txusrclk_in,
        gt18_txusrclk2_in               =>      gt18_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt18_txdlyen_in                 =>      gt18_txdlyen_i,
        gt18_txdlysreset_in             =>      gt18_txdlysreset_i,
        gt18_txdlysresetdone_out        =>      gt18_txdlysresetdone_i,
        gt18_txphalign_in               =>      gt18_txphalign_i,
        gt18_txphaligndone_out          =>      gt18_txphaligndone_i,
        gt18_txphalignen_in             =>      gt18_txphalignen_i,
        gt18_txphdlyreset_in            =>      gt18_txphdlyreset_i,
        gt18_txphinit_in                =>      gt18_txphinit_i,
        gt18_txphinitdone_out           =>      gt18_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt18_txdata_in                  =>      gt18_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt18_gthtxn_out                 =>      gt18_gthtxn_out,
        gt18_gthtxp_out                 =>      gt18_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt18_txoutclk_out               =>      gt18_txoutclk_i,
        gt18_txoutclkfabric_out         =>      gt18_txoutclkfabric_out,
        gt18_txoutclkpcs_out            =>      gt18_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt18_txresetdone_out            =>      gt18_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt18_txcharisk_in               =>      gt18_txcharisk_in,


        GT19_DRP_BUSY_OUT               =>      GT19_DRP_BUSY_OUT,
        GT19_RXPMARESETDONE_OUT         =>      gt19_rxpmaresetdone_i,
        GT19_TXPMARESETDONE_OUT         =>      gt19_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT19  (X1Y23)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt19_drpaddr_in                 =>      gt19_drpaddr_in,
        gt19_drpclk_in                  =>      gt19_drpclk_in,
        gt19_drpdi_in                   =>      gt19_drpdi_in,
        gt19_drpdo_out                  =>      gt19_drpdo_out,
        gt19_drpen_in                   =>      gt19_drpen_in,
        gt19_drprdy_out                 =>      gt19_drprdy_out,
        gt19_drpwe_in                   =>      gt19_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt19_eyescanreset_in            =>      gt19_eyescanreset_in,
        gt19_rxuserrdy_in               =>      gt19_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt19_eyescandataerror_out       =>      gt19_eyescandataerror_out,
        gt19_eyescantrigger_in          =>      gt19_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt19_rxslide_in                 =>      gt19_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt19_dmonitorout_out            =>      gt19_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt19_rxusrclk_in                =>      gt19_rxusrclk_in,
        gt19_rxusrclk2_in               =>      gt19_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt19_rxdata_out                 =>      gt19_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt19_rxdisperr_out              =>      gt19_rxdisperr_out,
        gt19_rxnotintable_out           =>      gt19_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt19_gthrxn_in                  =>      gt19_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt19_rxdlyen_in                 =>      gt19_rxdlyen_i,
        gt19_rxdlysreset_in             =>      gt19_rxdlysreset_i,
        gt19_rxdlysresetdone_out        =>      gt19_rxdlysresetdone_i,
        gt19_rxphalign_in               =>      gt19_rxphalign_i,
        gt19_rxphaligndone_out          =>      gt19_rxphaligndone_i,
        gt19_rxphalignen_in             =>      gt19_rxphalignen_i,
        gt19_rxphdlyreset_in            =>      gt19_rxphdlyreset_i,
        gt19_rxphmonitor_out            =>      gt19_rxphmonitor_out,
        gt19_rxphslipmonitor_out        =>      gt19_rxphslipmonitor_out,
        gt19_rxsyncallin_in             =>      gt19_rxsyncallin_i,
        gt19_rxsyncdone_out             =>      gt19_rxsyncdone_i,
        gt19_rxsyncin_in                =>      gt19_rxsyncin_i,
        gt19_rxsyncmode_in              =>      gt19_rxsyncmode_i,
        gt19_rxsyncout_out              =>      gt19_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt19_rxbyteisaligned_out        =>      gt19_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt19_rxlpmhfhold_in             =>      gt19_rxlpmhfhold_i,
        gt19_rxlpmlfhold_in             =>      gt19_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt19_rxmonitorout_out           =>      gt19_rxmonitorout_out,
        gt19_rxmonitorsel_in            =>      gt19_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt19_rxoutclk_out               =>      gt19_rxoutclk_i,
        gt19_rxoutclkfabric_out         =>      gt19_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt19_gtrxreset_in               =>      gt19_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt19_rxcharisk_out              =>      gt19_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt19_gthrxp_in                  =>      gt19_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt19_rxresetdone_out            =>      gt19_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt19_gttxreset_in               =>      gt19_gttxreset_i,
        gt19_txuserrdy_in               =>      gt19_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt19_txusrclk_in                =>      gt19_txusrclk_in,
        gt19_txusrclk2_in               =>      gt19_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt19_txdlyen_in                 =>      gt19_txdlyen_i,
        gt19_txdlysreset_in             =>      gt19_txdlysreset_i,
        gt19_txdlysresetdone_out        =>      gt19_txdlysresetdone_i,
        gt19_txphalign_in               =>      gt19_txphalign_i,
        gt19_txphaligndone_out          =>      gt19_txphaligndone_i,
        gt19_txphalignen_in             =>      gt19_txphalignen_i,
        gt19_txphdlyreset_in            =>      gt19_txphdlyreset_i,
        gt19_txphinit_in                =>      gt19_txphinit_i,
        gt19_txphinitdone_out           =>      gt19_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt19_txdata_in                  =>      gt19_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt19_gthtxn_out                 =>      gt19_gthtxn_out,
        gt19_gthtxp_out                 =>      gt19_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt19_txoutclk_out               =>      gt19_txoutclk_i,
        gt19_txoutclkfabric_out         =>      gt19_txoutclkfabric_out,
        gt19_txoutclkpcs_out            =>      gt19_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt19_txresetdone_out            =>      gt19_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt19_txcharisk_in               =>      gt19_txcharisk_in,


        GT20_DRP_BUSY_OUT               =>      GT20_DRP_BUSY_OUT,
        GT20_RXPMARESETDONE_OUT         =>      gt20_rxpmaresetdone_i,
        GT20_TXPMARESETDONE_OUT         =>      gt20_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT20  (X1Y24)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt20_drpaddr_in                 =>      gt20_drpaddr_in,
        gt20_drpclk_in                  =>      gt20_drpclk_in,
        gt20_drpdi_in                   =>      gt20_drpdi_in,
        gt20_drpdo_out                  =>      gt20_drpdo_out,
        gt20_drpen_in                   =>      gt20_drpen_in,
        gt20_drprdy_out                 =>      gt20_drprdy_out,
        gt20_drpwe_in                   =>      gt20_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt20_eyescanreset_in            =>      gt20_eyescanreset_in,
        gt20_rxuserrdy_in               =>      gt20_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt20_eyescandataerror_out       =>      gt20_eyescandataerror_out,
        gt20_eyescantrigger_in          =>      gt20_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt20_rxslide_in                 =>      gt20_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt20_dmonitorout_out            =>      gt20_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt20_rxusrclk_in                =>      gt20_rxusrclk_in,
        gt20_rxusrclk2_in               =>      gt20_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt20_rxdata_out                 =>      gt20_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt20_rxdisperr_out              =>      gt20_rxdisperr_out,
        gt20_rxnotintable_out           =>      gt20_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt20_gthrxn_in                  =>      gt20_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt20_rxdlyen_in                 =>      gt20_rxdlyen_i,
        gt20_rxdlysreset_in             =>      gt20_rxdlysreset_i,
        gt20_rxdlysresetdone_out        =>      gt20_rxdlysresetdone_i,
        gt20_rxphalign_in               =>      gt20_rxphalign_i,
        gt20_rxphaligndone_out          =>      gt20_rxphaligndone_i,
        gt20_rxphalignen_in             =>      gt20_rxphalignen_i,
        gt20_rxphdlyreset_in            =>      gt20_rxphdlyreset_i,
        gt20_rxphmonitor_out            =>      gt20_rxphmonitor_out,
        gt20_rxphslipmonitor_out        =>      gt20_rxphslipmonitor_out,
        gt20_rxsyncallin_in             =>      gt20_rxsyncallin_i,
        gt20_rxsyncdone_out             =>      gt20_rxsyncdone_i,
        gt20_rxsyncin_in                =>      gt20_rxsyncin_i,
        gt20_rxsyncmode_in              =>      gt20_rxsyncmode_i,
        gt20_rxsyncout_out              =>      gt20_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt20_rxbyteisaligned_out        =>      gt20_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt20_rxlpmhfhold_in             =>      gt20_rxlpmhfhold_i,
        gt20_rxlpmlfhold_in             =>      gt20_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt20_rxmonitorout_out           =>      gt20_rxmonitorout_out,
        gt20_rxmonitorsel_in            =>      gt20_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt20_rxoutclk_out               =>      gt20_rxoutclk_i,
        gt20_rxoutclkfabric_out         =>      gt20_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt20_gtrxreset_in               =>      gt20_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt20_rxcharisk_out              =>      gt20_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt20_gthrxp_in                  =>      gt20_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt20_rxresetdone_out            =>      gt20_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt20_gttxreset_in               =>      gt20_gttxreset_i,
        gt20_txuserrdy_in               =>      gt20_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt20_txusrclk_in                =>      gt20_txusrclk_in,
        gt20_txusrclk2_in               =>      gt20_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt20_txdlyen_in                 =>      gt20_txdlyen_i,
        gt20_txdlysreset_in             =>      gt20_txdlysreset_i,
        gt20_txdlysresetdone_out        =>      gt20_txdlysresetdone_i,
        gt20_txphalign_in               =>      gt20_txphalign_i,
        gt20_txphaligndone_out          =>      gt20_txphaligndone_i,
        gt20_txphalignen_in             =>      gt20_txphalignen_i,
        gt20_txphdlyreset_in            =>      gt20_txphdlyreset_i,
        gt20_txphinit_in                =>      gt20_txphinit_i,
        gt20_txphinitdone_out           =>      gt20_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt20_txdata_in                  =>      gt20_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt20_gthtxn_out                 =>      gt20_gthtxn_out,
        gt20_gthtxp_out                 =>      gt20_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt20_txoutclk_out               =>      gt20_txoutclk_i,
        gt20_txoutclkfabric_out         =>      gt20_txoutclkfabric_out,
        gt20_txoutclkpcs_out            =>      gt20_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt20_txresetdone_out            =>      gt20_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt20_txcharisk_in               =>      gt20_txcharisk_in,


        GT21_DRP_BUSY_OUT               =>      GT21_DRP_BUSY_OUT,
        GT21_RXPMARESETDONE_OUT         =>      gt21_rxpmaresetdone_i,
        GT21_TXPMARESETDONE_OUT         =>      gt21_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT21  (X1Y25)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt21_drpaddr_in                 =>      gt21_drpaddr_in,
        gt21_drpclk_in                  =>      gt21_drpclk_in,
        gt21_drpdi_in                   =>      gt21_drpdi_in,
        gt21_drpdo_out                  =>      gt21_drpdo_out,
        gt21_drpen_in                   =>      gt21_drpen_in,
        gt21_drprdy_out                 =>      gt21_drprdy_out,
        gt21_drpwe_in                   =>      gt21_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt21_eyescanreset_in            =>      gt21_eyescanreset_in,
        gt21_rxuserrdy_in               =>      gt21_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt21_eyescandataerror_out       =>      gt21_eyescandataerror_out,
        gt21_eyescantrigger_in          =>      gt21_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt21_rxslide_in                 =>      gt21_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt21_dmonitorout_out            =>      gt21_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt21_rxusrclk_in                =>      gt21_rxusrclk_in,
        gt21_rxusrclk2_in               =>      gt21_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt21_rxdata_out                 =>      gt21_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt21_rxdisperr_out              =>      gt21_rxdisperr_out,
        gt21_rxnotintable_out           =>      gt21_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt21_gthrxn_in                  =>      gt21_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt21_rxdlyen_in                 =>      gt21_rxdlyen_i,
        gt21_rxdlysreset_in             =>      gt21_rxdlysreset_i,
        gt21_rxdlysresetdone_out        =>      gt21_rxdlysresetdone_i,
        gt21_rxphalign_in               =>      gt21_rxphalign_i,
        gt21_rxphaligndone_out          =>      gt21_rxphaligndone_i,
        gt21_rxphalignen_in             =>      gt21_rxphalignen_i,
        gt21_rxphdlyreset_in            =>      gt21_rxphdlyreset_i,
        gt21_rxphmonitor_out            =>      gt21_rxphmonitor_out,
        gt21_rxphslipmonitor_out        =>      gt21_rxphslipmonitor_out,
        gt21_rxsyncallin_in             =>      gt21_rxsyncallin_i,
        gt21_rxsyncdone_out             =>      gt21_rxsyncdone_i,
        gt21_rxsyncin_in                =>      gt21_rxsyncin_i,
        gt21_rxsyncmode_in              =>      gt21_rxsyncmode_i,
        gt21_rxsyncout_out              =>      gt21_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt21_rxbyteisaligned_out        =>      gt21_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt21_rxlpmhfhold_in             =>      gt21_rxlpmhfhold_i,
        gt21_rxlpmlfhold_in             =>      gt21_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt21_rxmonitorout_out           =>      gt21_rxmonitorout_out,
        gt21_rxmonitorsel_in            =>      gt21_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt21_rxoutclk_out               =>      gt21_rxoutclk_i,
        gt21_rxoutclkfabric_out         =>      gt21_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt21_gtrxreset_in               =>      gt21_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt21_rxcharisk_out              =>      gt21_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt21_gthrxp_in                  =>      gt21_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt21_rxresetdone_out            =>      gt21_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt21_gttxreset_in               =>      gt21_gttxreset_i,
        gt21_txuserrdy_in               =>      gt21_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt21_txusrclk_in                =>      gt21_txusrclk_in,
        gt21_txusrclk2_in               =>      gt21_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt21_txdlyen_in                 =>      gt21_txdlyen_i,
        gt21_txdlysreset_in             =>      gt21_txdlysreset_i,
        gt21_txdlysresetdone_out        =>      gt21_txdlysresetdone_i,
        gt21_txphalign_in               =>      gt21_txphalign_i,
        gt21_txphaligndone_out          =>      gt21_txphaligndone_i,
        gt21_txphalignen_in             =>      gt21_txphalignen_i,
        gt21_txphdlyreset_in            =>      gt21_txphdlyreset_i,
        gt21_txphinit_in                =>      gt21_txphinit_i,
        gt21_txphinitdone_out           =>      gt21_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt21_txdata_in                  =>      gt21_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt21_gthtxn_out                 =>      gt21_gthtxn_out,
        gt21_gthtxp_out                 =>      gt21_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt21_txoutclk_out               =>      gt21_txoutclk_i,
        gt21_txoutclkfabric_out         =>      gt21_txoutclkfabric_out,
        gt21_txoutclkpcs_out            =>      gt21_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt21_txresetdone_out            =>      gt21_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt21_txcharisk_in               =>      gt21_txcharisk_in,


        GT22_DRP_BUSY_OUT               =>      GT22_DRP_BUSY_OUT,
        GT22_RXPMARESETDONE_OUT         =>      gt22_rxpmaresetdone_i,
        GT22_TXPMARESETDONE_OUT         =>      gt22_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT22  (X1Y26)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt22_drpaddr_in                 =>      gt22_drpaddr_in,
        gt22_drpclk_in                  =>      gt22_drpclk_in,
        gt22_drpdi_in                   =>      gt22_drpdi_in,
        gt22_drpdo_out                  =>      gt22_drpdo_out,
        gt22_drpen_in                   =>      gt22_drpen_in,
        gt22_drprdy_out                 =>      gt22_drprdy_out,
        gt22_drpwe_in                   =>      gt22_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt22_eyescanreset_in            =>      gt22_eyescanreset_in,
        gt22_rxuserrdy_in               =>      gt22_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt22_eyescandataerror_out       =>      gt22_eyescandataerror_out,
        gt22_eyescantrigger_in          =>      gt22_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt22_rxslide_in                 =>      gt22_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt22_dmonitorout_out            =>      gt22_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt22_rxusrclk_in                =>      gt22_rxusrclk_in,
        gt22_rxusrclk2_in               =>      gt22_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt22_rxdata_out                 =>      gt22_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt22_rxdisperr_out              =>      gt22_rxdisperr_out,
        gt22_rxnotintable_out           =>      gt22_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt22_gthrxn_in                  =>      gt22_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt22_rxdlyen_in                 =>      gt22_rxdlyen_i,
        gt22_rxdlysreset_in             =>      gt22_rxdlysreset_i,
        gt22_rxdlysresetdone_out        =>      gt22_rxdlysresetdone_i,
        gt22_rxphalign_in               =>      gt22_rxphalign_i,
        gt22_rxphaligndone_out          =>      gt22_rxphaligndone_i,
        gt22_rxphalignen_in             =>      gt22_rxphalignen_i,
        gt22_rxphdlyreset_in            =>      gt22_rxphdlyreset_i,
        gt22_rxphmonitor_out            =>      gt22_rxphmonitor_out,
        gt22_rxphslipmonitor_out        =>      gt22_rxphslipmonitor_out,
        gt22_rxsyncallin_in             =>      gt22_rxsyncallin_i,
        gt22_rxsyncdone_out             =>      gt22_rxsyncdone_i,
        gt22_rxsyncin_in                =>      gt22_rxsyncin_i,
        gt22_rxsyncmode_in              =>      gt22_rxsyncmode_i,
        gt22_rxsyncout_out              =>      gt22_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt22_rxbyteisaligned_out        =>      gt22_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt22_rxlpmhfhold_in             =>      gt22_rxlpmhfhold_i,
        gt22_rxlpmlfhold_in             =>      gt22_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt22_rxmonitorout_out           =>      gt22_rxmonitorout_out,
        gt22_rxmonitorsel_in            =>      gt22_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt22_rxoutclk_out               =>      gt22_rxoutclk_i,
        gt22_rxoutclkfabric_out         =>      gt22_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt22_gtrxreset_in               =>      gt22_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt22_rxcharisk_out              =>      gt22_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt22_gthrxp_in                  =>      gt22_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt22_rxresetdone_out            =>      gt22_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt22_gttxreset_in               =>      gt22_gttxreset_i,
        gt22_txuserrdy_in               =>      gt22_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt22_txusrclk_in                =>      gt22_txusrclk_in,
        gt22_txusrclk2_in               =>      gt22_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt22_txdlyen_in                 =>      gt22_txdlyen_i,
        gt22_txdlysreset_in             =>      gt22_txdlysreset_i,
        gt22_txdlysresetdone_out        =>      gt22_txdlysresetdone_i,
        gt22_txphalign_in               =>      gt22_txphalign_i,
        gt22_txphaligndone_out          =>      gt22_txphaligndone_i,
        gt22_txphalignen_in             =>      gt22_txphalignen_i,
        gt22_txphdlyreset_in            =>      gt22_txphdlyreset_i,
        gt22_txphinit_in                =>      gt22_txphinit_i,
        gt22_txphinitdone_out           =>      gt22_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt22_txdata_in                  =>      gt22_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt22_gthtxn_out                 =>      gt22_gthtxn_out,
        gt22_gthtxp_out                 =>      gt22_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt22_txoutclk_out               =>      gt22_txoutclk_i,
        gt22_txoutclkfabric_out         =>      gt22_txoutclkfabric_out,
        gt22_txoutclkpcs_out            =>      gt22_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt22_txresetdone_out            =>      gt22_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt22_txcharisk_in               =>      gt22_txcharisk_in,


        GT23_DRP_BUSY_OUT               =>      GT23_DRP_BUSY_OUT,
        GT23_RXPMARESETDONE_OUT         =>      gt23_rxpmaresetdone_i,
        GT23_TXPMARESETDONE_OUT         =>      gt23_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT23  (X1Y27)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt23_drpaddr_in                 =>      gt23_drpaddr_in,
        gt23_drpclk_in                  =>      gt23_drpclk_in,
        gt23_drpdi_in                   =>      gt23_drpdi_in,
        gt23_drpdo_out                  =>      gt23_drpdo_out,
        gt23_drpen_in                   =>      gt23_drpen_in,
        gt23_drprdy_out                 =>      gt23_drprdy_out,
        gt23_drpwe_in                   =>      gt23_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt23_eyescanreset_in            =>      gt23_eyescanreset_in,
        gt23_rxuserrdy_in               =>      gt23_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt23_eyescandataerror_out       =>      gt23_eyescandataerror_out,
        gt23_eyescantrigger_in          =>      gt23_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt23_rxslide_in                 =>      gt23_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt23_dmonitorout_out            =>      gt23_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt23_rxusrclk_in                =>      gt23_rxusrclk_in,
        gt23_rxusrclk2_in               =>      gt23_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt23_rxdata_out                 =>      gt23_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt23_rxdisperr_out              =>      gt23_rxdisperr_out,
        gt23_rxnotintable_out           =>      gt23_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt23_gthrxn_in                  =>      gt23_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt23_rxdlyen_in                 =>      gt23_rxdlyen_i,
        gt23_rxdlysreset_in             =>      gt23_rxdlysreset_i,
        gt23_rxdlysresetdone_out        =>      gt23_rxdlysresetdone_i,
        gt23_rxphalign_in               =>      gt23_rxphalign_i,
        gt23_rxphaligndone_out          =>      gt23_rxphaligndone_i,
        gt23_rxphalignen_in             =>      gt23_rxphalignen_i,
        gt23_rxphdlyreset_in            =>      gt23_rxphdlyreset_i,
        gt23_rxphmonitor_out            =>      gt23_rxphmonitor_out,
        gt23_rxphslipmonitor_out        =>      gt23_rxphslipmonitor_out,
        gt23_rxsyncallin_in             =>      gt23_rxsyncallin_i,
        gt23_rxsyncdone_out             =>      gt23_rxsyncdone_i,
        gt23_rxsyncin_in                =>      gt23_rxsyncin_i,
        gt23_rxsyncmode_in              =>      gt23_rxsyncmode_i,
        gt23_rxsyncout_out              =>      gt23_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt23_rxbyteisaligned_out        =>      gt23_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt23_rxlpmhfhold_in             =>      gt23_rxlpmhfhold_i,
        gt23_rxlpmlfhold_in             =>      gt23_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt23_rxmonitorout_out           =>      gt23_rxmonitorout_out,
        gt23_rxmonitorsel_in            =>      gt23_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt23_rxoutclk_out               =>      gt23_rxoutclk_i,
        gt23_rxoutclkfabric_out         =>      gt23_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt23_gtrxreset_in               =>      gt23_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt23_rxcharisk_out              =>      gt23_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt23_gthrxp_in                  =>      gt23_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt23_rxresetdone_out            =>      gt23_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt23_gttxreset_in               =>      gt23_gttxreset_i,
        gt23_txuserrdy_in               =>      gt23_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt23_txusrclk_in                =>      gt23_txusrclk_in,
        gt23_txusrclk2_in               =>      gt23_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt23_txdlyen_in                 =>      gt23_txdlyen_i,
        gt23_txdlysreset_in             =>      gt23_txdlysreset_i,
        gt23_txdlysresetdone_out        =>      gt23_txdlysresetdone_i,
        gt23_txphalign_in               =>      gt23_txphalign_i,
        gt23_txphaligndone_out          =>      gt23_txphaligndone_i,
        gt23_txphalignen_in             =>      gt23_txphalignen_i,
        gt23_txphdlyreset_in            =>      gt23_txphdlyreset_i,
        gt23_txphinit_in                =>      gt23_txphinit_i,
        gt23_txphinitdone_out           =>      gt23_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt23_txdata_in                  =>      gt23_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt23_gthtxn_out                 =>      gt23_gthtxn_out,
        gt23_gthtxp_out                 =>      gt23_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt23_txoutclk_out               =>      gt23_txoutclk_i,
        gt23_txoutclkfabric_out         =>      gt23_txoutclkfabric_out,
        gt23_txoutclkpcs_out            =>      gt23_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt23_txresetdone_out            =>      gt23_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt23_txcharisk_in               =>      gt23_txcharisk_in,


        GT24_DRP_BUSY_OUT               =>      GT24_DRP_BUSY_OUT,
        GT24_RXPMARESETDONE_OUT         =>      gt24_rxpmaresetdone_i,
        GT24_TXPMARESETDONE_OUT         =>      gt24_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT24  (X1Y28)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt24_drpaddr_in                 =>      gt24_drpaddr_in,
        gt24_drpclk_in                  =>      gt24_drpclk_in,
        gt24_drpdi_in                   =>      gt24_drpdi_in,
        gt24_drpdo_out                  =>      gt24_drpdo_out,
        gt24_drpen_in                   =>      gt24_drpen_in,
        gt24_drprdy_out                 =>      gt24_drprdy_out,
        gt24_drpwe_in                   =>      gt24_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt24_eyescanreset_in            =>      gt24_eyescanreset_in,
        gt24_rxuserrdy_in               =>      gt24_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt24_eyescandataerror_out       =>      gt24_eyescandataerror_out,
        gt24_eyescantrigger_in          =>      gt24_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt24_rxslide_in                 =>      gt24_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt24_dmonitorout_out            =>      gt24_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt24_rxusrclk_in                =>      gt24_rxusrclk_in,
        gt24_rxusrclk2_in               =>      gt24_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt24_rxdata_out                 =>      gt24_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt24_rxdisperr_out              =>      gt24_rxdisperr_out,
        gt24_rxnotintable_out           =>      gt24_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt24_gthrxn_in                  =>      gt24_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt24_rxdlyen_in                 =>      gt24_rxdlyen_i,
        gt24_rxdlysreset_in             =>      gt24_rxdlysreset_i,
        gt24_rxdlysresetdone_out        =>      gt24_rxdlysresetdone_i,
        gt24_rxphalign_in               =>      gt24_rxphalign_i,
        gt24_rxphaligndone_out          =>      gt24_rxphaligndone_i,
        gt24_rxphalignen_in             =>      gt24_rxphalignen_i,
        gt24_rxphdlyreset_in            =>      gt24_rxphdlyreset_i,
        gt24_rxphmonitor_out            =>      gt24_rxphmonitor_out,
        gt24_rxphslipmonitor_out        =>      gt24_rxphslipmonitor_out,
        gt24_rxsyncallin_in             =>      gt24_rxsyncallin_i,
        gt24_rxsyncdone_out             =>      gt24_rxsyncdone_i,
        gt24_rxsyncin_in                =>      gt24_rxsyncin_i,
        gt24_rxsyncmode_in              =>      gt24_rxsyncmode_i,
        gt24_rxsyncout_out              =>      gt24_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt24_rxbyteisaligned_out        =>      gt24_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt24_rxlpmhfhold_in             =>      gt24_rxlpmhfhold_i,
        gt24_rxlpmlfhold_in             =>      gt24_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt24_rxmonitorout_out           =>      gt24_rxmonitorout_out,
        gt24_rxmonitorsel_in            =>      gt24_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt24_rxoutclk_out               =>      gt24_rxoutclk_i,
        gt24_rxoutclkfabric_out         =>      gt24_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt24_gtrxreset_in               =>      gt24_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt24_rxcharisk_out              =>      gt24_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt24_gthrxp_in                  =>      gt24_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt24_rxresetdone_out            =>      gt24_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt24_gttxreset_in               =>      gt24_gttxreset_i,
        gt24_txuserrdy_in               =>      gt24_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt24_txusrclk_in                =>      gt24_txusrclk_in,
        gt24_txusrclk2_in               =>      gt24_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt24_txdlyen_in                 =>      gt24_txdlyen_i,
        gt24_txdlysreset_in             =>      gt24_txdlysreset_i,
        gt24_txdlysresetdone_out        =>      gt24_txdlysresetdone_i,
        gt24_txphalign_in               =>      gt24_txphalign_i,
        gt24_txphaligndone_out          =>      gt24_txphaligndone_i,
        gt24_txphalignen_in             =>      gt24_txphalignen_i,
        gt24_txphdlyreset_in            =>      gt24_txphdlyreset_i,
        gt24_txphinit_in                =>      gt24_txphinit_i,
        gt24_txphinitdone_out           =>      gt24_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt24_txdata_in                  =>      gt24_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt24_gthtxn_out                 =>      gt24_gthtxn_out,
        gt24_gthtxp_out                 =>      gt24_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt24_txoutclk_out               =>      gt24_txoutclk_i,
        gt24_txoutclkfabric_out         =>      gt24_txoutclkfabric_out,
        gt24_txoutclkpcs_out            =>      gt24_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt24_txresetdone_out            =>      gt24_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt24_txcharisk_in               =>      gt24_txcharisk_in,


        GT25_DRP_BUSY_OUT               =>      GT25_DRP_BUSY_OUT,
        GT25_RXPMARESETDONE_OUT         =>      gt25_rxpmaresetdone_i,
        GT25_TXPMARESETDONE_OUT         =>      gt25_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT25  (X1Y29)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt25_drpaddr_in                 =>      gt25_drpaddr_in,
        gt25_drpclk_in                  =>      gt25_drpclk_in,
        gt25_drpdi_in                   =>      gt25_drpdi_in,
        gt25_drpdo_out                  =>      gt25_drpdo_out,
        gt25_drpen_in                   =>      gt25_drpen_in,
        gt25_drprdy_out                 =>      gt25_drprdy_out,
        gt25_drpwe_in                   =>      gt25_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt25_eyescanreset_in            =>      gt25_eyescanreset_in,
        gt25_rxuserrdy_in               =>      gt25_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt25_eyescandataerror_out       =>      gt25_eyescandataerror_out,
        gt25_eyescantrigger_in          =>      gt25_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt25_rxslide_in                 =>      gt25_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt25_dmonitorout_out            =>      gt25_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt25_rxusrclk_in                =>      gt25_rxusrclk_in,
        gt25_rxusrclk2_in               =>      gt25_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt25_rxdata_out                 =>      gt25_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt25_rxdisperr_out              =>      gt25_rxdisperr_out,
        gt25_rxnotintable_out           =>      gt25_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt25_gthrxn_in                  =>      gt25_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt25_rxdlyen_in                 =>      gt25_rxdlyen_i,
        gt25_rxdlysreset_in             =>      gt25_rxdlysreset_i,
        gt25_rxdlysresetdone_out        =>      gt25_rxdlysresetdone_i,
        gt25_rxphalign_in               =>      gt25_rxphalign_i,
        gt25_rxphaligndone_out          =>      gt25_rxphaligndone_i,
        gt25_rxphalignen_in             =>      gt25_rxphalignen_i,
        gt25_rxphdlyreset_in            =>      gt25_rxphdlyreset_i,
        gt25_rxphmonitor_out            =>      gt25_rxphmonitor_out,
        gt25_rxphslipmonitor_out        =>      gt25_rxphslipmonitor_out,
        gt25_rxsyncallin_in             =>      gt25_rxsyncallin_i,
        gt25_rxsyncdone_out             =>      gt25_rxsyncdone_i,
        gt25_rxsyncin_in                =>      gt25_rxsyncin_i,
        gt25_rxsyncmode_in              =>      gt25_rxsyncmode_i,
        gt25_rxsyncout_out              =>      gt25_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt25_rxbyteisaligned_out        =>      gt25_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt25_rxlpmhfhold_in             =>      gt25_rxlpmhfhold_i,
        gt25_rxlpmlfhold_in             =>      gt25_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt25_rxmonitorout_out           =>      gt25_rxmonitorout_out,
        gt25_rxmonitorsel_in            =>      gt25_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt25_rxoutclk_out               =>      gt25_rxoutclk_i,
        gt25_rxoutclkfabric_out         =>      gt25_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt25_gtrxreset_in               =>      gt25_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt25_rxcharisk_out              =>      gt25_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt25_gthrxp_in                  =>      gt25_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt25_rxresetdone_out            =>      gt25_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt25_gttxreset_in               =>      gt25_gttxreset_i,
        gt25_txuserrdy_in               =>      gt25_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt25_txusrclk_in                =>      gt25_txusrclk_in,
        gt25_txusrclk2_in               =>      gt25_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt25_txdlyen_in                 =>      gt25_txdlyen_i,
        gt25_txdlysreset_in             =>      gt25_txdlysreset_i,
        gt25_txdlysresetdone_out        =>      gt25_txdlysresetdone_i,
        gt25_txphalign_in               =>      gt25_txphalign_i,
        gt25_txphaligndone_out          =>      gt25_txphaligndone_i,
        gt25_txphalignen_in             =>      gt25_txphalignen_i,
        gt25_txphdlyreset_in            =>      gt25_txphdlyreset_i,
        gt25_txphinit_in                =>      gt25_txphinit_i,
        gt25_txphinitdone_out           =>      gt25_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt25_txdata_in                  =>      gt25_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt25_gthtxn_out                 =>      gt25_gthtxn_out,
        gt25_gthtxp_out                 =>      gt25_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt25_txoutclk_out               =>      gt25_txoutclk_i,
        gt25_txoutclkfabric_out         =>      gt25_txoutclkfabric_out,
        gt25_txoutclkpcs_out            =>      gt25_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt25_txresetdone_out            =>      gt25_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt25_txcharisk_in               =>      gt25_txcharisk_in,


        GT26_DRP_BUSY_OUT               =>      GT26_DRP_BUSY_OUT,
        GT26_RXPMARESETDONE_OUT         =>      gt26_rxpmaresetdone_i,
        GT26_TXPMARESETDONE_OUT         =>      gt26_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT26  (X1Y30)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt26_drpaddr_in                 =>      gt26_drpaddr_in,
        gt26_drpclk_in                  =>      gt26_drpclk_in,
        gt26_drpdi_in                   =>      gt26_drpdi_in,
        gt26_drpdo_out                  =>      gt26_drpdo_out,
        gt26_drpen_in                   =>      gt26_drpen_in,
        gt26_drprdy_out                 =>      gt26_drprdy_out,
        gt26_drpwe_in                   =>      gt26_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt26_eyescanreset_in            =>      gt26_eyescanreset_in,
        gt26_rxuserrdy_in               =>      gt26_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt26_eyescandataerror_out       =>      gt26_eyescandataerror_out,
        gt26_eyescantrigger_in          =>      gt26_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt26_rxslide_in                 =>      gt26_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt26_dmonitorout_out            =>      gt26_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt26_rxusrclk_in                =>      gt26_rxusrclk_in,
        gt26_rxusrclk2_in               =>      gt26_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt26_rxdata_out                 =>      gt26_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt26_rxdisperr_out              =>      gt26_rxdisperr_out,
        gt26_rxnotintable_out           =>      gt26_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt26_gthrxn_in                  =>      gt26_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt26_rxdlyen_in                 =>      gt26_rxdlyen_i,
        gt26_rxdlysreset_in             =>      gt26_rxdlysreset_i,
        gt26_rxdlysresetdone_out        =>      gt26_rxdlysresetdone_i,
        gt26_rxphalign_in               =>      gt26_rxphalign_i,
        gt26_rxphaligndone_out          =>      gt26_rxphaligndone_i,
        gt26_rxphalignen_in             =>      gt26_rxphalignen_i,
        gt26_rxphdlyreset_in            =>      gt26_rxphdlyreset_i,
        gt26_rxphmonitor_out            =>      gt26_rxphmonitor_out,
        gt26_rxphslipmonitor_out        =>      gt26_rxphslipmonitor_out,
        gt26_rxsyncallin_in             =>      gt26_rxsyncallin_i,
        gt26_rxsyncdone_out             =>      gt26_rxsyncdone_i,
        gt26_rxsyncin_in                =>      gt26_rxsyncin_i,
        gt26_rxsyncmode_in              =>      gt26_rxsyncmode_i,
        gt26_rxsyncout_out              =>      gt26_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt26_rxbyteisaligned_out        =>      gt26_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt26_rxlpmhfhold_in             =>      gt26_rxlpmhfhold_i,
        gt26_rxlpmlfhold_in             =>      gt26_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt26_rxmonitorout_out           =>      gt26_rxmonitorout_out,
        gt26_rxmonitorsel_in            =>      gt26_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt26_rxoutclk_out               =>      gt26_rxoutclk_i,
        gt26_rxoutclkfabric_out         =>      gt26_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt26_gtrxreset_in               =>      gt26_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt26_rxcharisk_out              =>      gt26_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt26_gthrxp_in                  =>      gt26_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt26_rxresetdone_out            =>      gt26_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt26_gttxreset_in               =>      gt26_gttxreset_i,
        gt26_txuserrdy_in               =>      gt26_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt26_txusrclk_in                =>      gt26_txusrclk_in,
        gt26_txusrclk2_in               =>      gt26_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt26_txdlyen_in                 =>      gt26_txdlyen_i,
        gt26_txdlysreset_in             =>      gt26_txdlysreset_i,
        gt26_txdlysresetdone_out        =>      gt26_txdlysresetdone_i,
        gt26_txphalign_in               =>      gt26_txphalign_i,
        gt26_txphaligndone_out          =>      gt26_txphaligndone_i,
        gt26_txphalignen_in             =>      gt26_txphalignen_i,
        gt26_txphdlyreset_in            =>      gt26_txphdlyreset_i,
        gt26_txphinit_in                =>      gt26_txphinit_i,
        gt26_txphinitdone_out           =>      gt26_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt26_txdata_in                  =>      gt26_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt26_gthtxn_out                 =>      gt26_gthtxn_out,
        gt26_gthtxp_out                 =>      gt26_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt26_txoutclk_out               =>      gt26_txoutclk_i,
        gt26_txoutclkfabric_out         =>      gt26_txoutclkfabric_out,
        gt26_txoutclkpcs_out            =>      gt26_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt26_txresetdone_out            =>      gt26_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt26_txcharisk_in               =>      gt26_txcharisk_in,


        GT27_DRP_BUSY_OUT               =>      GT27_DRP_BUSY_OUT,
        GT27_RXPMARESETDONE_OUT         =>      gt27_rxpmaresetdone_i,
        GT27_TXPMARESETDONE_OUT         =>      gt27_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT27  (X1Y31)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt27_drpaddr_in                 =>      gt27_drpaddr_in,
        gt27_drpclk_in                  =>      gt27_drpclk_in,
        gt27_drpdi_in                   =>      gt27_drpdi_in,
        gt27_drpdo_out                  =>      gt27_drpdo_out,
        gt27_drpen_in                   =>      gt27_drpen_in,
        gt27_drprdy_out                 =>      gt27_drprdy_out,
        gt27_drpwe_in                   =>      gt27_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt27_eyescanreset_in            =>      gt27_eyescanreset_in,
        gt27_rxuserrdy_in               =>      gt27_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt27_eyescandataerror_out       =>      gt27_eyescandataerror_out,
        gt27_eyescantrigger_in          =>      gt27_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt27_rxslide_in                 =>      gt27_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt27_dmonitorout_out            =>      gt27_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt27_rxusrclk_in                =>      gt27_rxusrclk_in,
        gt27_rxusrclk2_in               =>      gt27_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt27_rxdata_out                 =>      gt27_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt27_rxdisperr_out              =>      gt27_rxdisperr_out,
        gt27_rxnotintable_out           =>      gt27_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt27_gthrxn_in                  =>      gt27_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt27_rxdlyen_in                 =>      gt27_rxdlyen_i,
        gt27_rxdlysreset_in             =>      gt27_rxdlysreset_i,
        gt27_rxdlysresetdone_out        =>      gt27_rxdlysresetdone_i,
        gt27_rxphalign_in               =>      gt27_rxphalign_i,
        gt27_rxphaligndone_out          =>      gt27_rxphaligndone_i,
        gt27_rxphalignen_in             =>      gt27_rxphalignen_i,
        gt27_rxphdlyreset_in            =>      gt27_rxphdlyreset_i,
        gt27_rxphmonitor_out            =>      gt27_rxphmonitor_out,
        gt27_rxphslipmonitor_out        =>      gt27_rxphslipmonitor_out,
        gt27_rxsyncallin_in             =>      gt27_rxsyncallin_i,
        gt27_rxsyncdone_out             =>      gt27_rxsyncdone_i,
        gt27_rxsyncin_in                =>      gt27_rxsyncin_i,
        gt27_rxsyncmode_in              =>      gt27_rxsyncmode_i,
        gt27_rxsyncout_out              =>      gt27_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt27_rxbyteisaligned_out        =>      gt27_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt27_rxlpmhfhold_in             =>      gt27_rxlpmhfhold_i,
        gt27_rxlpmlfhold_in             =>      gt27_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt27_rxmonitorout_out           =>      gt27_rxmonitorout_out,
        gt27_rxmonitorsel_in            =>      gt27_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt27_rxoutclk_out               =>      gt27_rxoutclk_i,
        gt27_rxoutclkfabric_out         =>      gt27_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt27_gtrxreset_in               =>      gt27_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt27_rxcharisk_out              =>      gt27_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt27_gthrxp_in                  =>      gt27_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt27_rxresetdone_out            =>      gt27_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt27_gttxreset_in               =>      gt27_gttxreset_i,
        gt27_txuserrdy_in               =>      gt27_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt27_txusrclk_in                =>      gt27_txusrclk_in,
        gt27_txusrclk2_in               =>      gt27_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt27_txdlyen_in                 =>      gt27_txdlyen_i,
        gt27_txdlysreset_in             =>      gt27_txdlysreset_i,
        gt27_txdlysresetdone_out        =>      gt27_txdlysresetdone_i,
        gt27_txphalign_in               =>      gt27_txphalign_i,
        gt27_txphaligndone_out          =>      gt27_txphaligndone_i,
        gt27_txphalignen_in             =>      gt27_txphalignen_i,
        gt27_txphdlyreset_in            =>      gt27_txphdlyreset_i,
        gt27_txphinit_in                =>      gt27_txphinit_i,
        gt27_txphinitdone_out           =>      gt27_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt27_txdata_in                  =>      gt27_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt27_gthtxn_out                 =>      gt27_gthtxn_out,
        gt27_gthtxp_out                 =>      gt27_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt27_txoutclk_out               =>      gt27_txoutclk_i,
        gt27_txoutclkfabric_out         =>      gt27_txoutclkfabric_out,
        gt27_txoutclkpcs_out            =>      gt27_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt27_txresetdone_out            =>      gt27_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt27_txcharisk_in               =>      gt27_txcharisk_in,


        GT28_DRP_BUSY_OUT               =>      GT28_DRP_BUSY_OUT,
        GT28_RXPMARESETDONE_OUT         =>      gt28_rxpmaresetdone_i,
        GT28_TXPMARESETDONE_OUT         =>      gt28_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT28  (X1Y32)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt28_drpaddr_in                 =>      gt28_drpaddr_in,
        gt28_drpclk_in                  =>      gt28_drpclk_in,
        gt28_drpdi_in                   =>      gt28_drpdi_in,
        gt28_drpdo_out                  =>      gt28_drpdo_out,
        gt28_drpen_in                   =>      gt28_drpen_in,
        gt28_drprdy_out                 =>      gt28_drprdy_out,
        gt28_drpwe_in                   =>      gt28_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt28_eyescanreset_in            =>      gt28_eyescanreset_in,
        gt28_rxuserrdy_in               =>      gt28_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt28_eyescandataerror_out       =>      gt28_eyescandataerror_out,
        gt28_eyescantrigger_in          =>      gt28_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt28_rxslide_in                 =>      gt28_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt28_dmonitorout_out            =>      gt28_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt28_rxusrclk_in                =>      gt28_rxusrclk_in,
        gt28_rxusrclk2_in               =>      gt28_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt28_rxdata_out                 =>      gt28_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt28_rxdisperr_out              =>      gt28_rxdisperr_out,
        gt28_rxnotintable_out           =>      gt28_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt28_gthrxn_in                  =>      gt28_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt28_rxdlyen_in                 =>      gt28_rxdlyen_i,
        gt28_rxdlysreset_in             =>      gt28_rxdlysreset_i,
        gt28_rxdlysresetdone_out        =>      gt28_rxdlysresetdone_i,
        gt28_rxphalign_in               =>      gt28_rxphalign_i,
        gt28_rxphaligndone_out          =>      gt28_rxphaligndone_i,
        gt28_rxphalignen_in             =>      gt28_rxphalignen_i,
        gt28_rxphdlyreset_in            =>      gt28_rxphdlyreset_i,
        gt28_rxphmonitor_out            =>      gt28_rxphmonitor_out,
        gt28_rxphslipmonitor_out        =>      gt28_rxphslipmonitor_out,
        gt28_rxsyncallin_in             =>      gt28_rxsyncallin_i,
        gt28_rxsyncdone_out             =>      gt28_rxsyncdone_i,
        gt28_rxsyncin_in                =>      gt28_rxsyncin_i,
        gt28_rxsyncmode_in              =>      gt28_rxsyncmode_i,
        gt28_rxsyncout_out              =>      gt28_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt28_rxbyteisaligned_out        =>      gt28_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt28_rxlpmhfhold_in             =>      gt28_rxlpmhfhold_i,
        gt28_rxlpmlfhold_in             =>      gt28_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt28_rxmonitorout_out           =>      gt28_rxmonitorout_out,
        gt28_rxmonitorsel_in            =>      gt28_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt28_rxoutclk_out               =>      gt28_rxoutclk_i,
        gt28_rxoutclkfabric_out         =>      gt28_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt28_gtrxreset_in               =>      gt28_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt28_rxcharisk_out              =>      gt28_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt28_gthrxp_in                  =>      gt28_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt28_rxresetdone_out            =>      gt28_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt28_gttxreset_in               =>      gt28_gttxreset_i,
        gt28_txuserrdy_in               =>      gt28_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt28_txusrclk_in                =>      gt28_txusrclk_in,
        gt28_txusrclk2_in               =>      gt28_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt28_txdlyen_in                 =>      gt28_txdlyen_i,
        gt28_txdlysreset_in             =>      gt28_txdlysreset_i,
        gt28_txdlysresetdone_out        =>      gt28_txdlysresetdone_i,
        gt28_txphalign_in               =>      gt28_txphalign_i,
        gt28_txphaligndone_out          =>      gt28_txphaligndone_i,
        gt28_txphalignen_in             =>      gt28_txphalignen_i,
        gt28_txphdlyreset_in            =>      gt28_txphdlyreset_i,
        gt28_txphinit_in                =>      gt28_txphinit_i,
        gt28_txphinitdone_out           =>      gt28_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt28_txdata_in                  =>      gt28_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt28_gthtxn_out                 =>      gt28_gthtxn_out,
        gt28_gthtxp_out                 =>      gt28_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt28_txoutclk_out               =>      gt28_txoutclk_i,
        gt28_txoutclkfabric_out         =>      gt28_txoutclkfabric_out,
        gt28_txoutclkpcs_out            =>      gt28_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt28_txresetdone_out            =>      gt28_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt28_txcharisk_in               =>      gt28_txcharisk_in,


        GT29_DRP_BUSY_OUT               =>      GT29_DRP_BUSY_OUT,
        GT29_RXPMARESETDONE_OUT         =>      gt29_rxpmaresetdone_i,
        GT29_TXPMARESETDONE_OUT         =>      gt29_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT29  (X1Y33)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt29_drpaddr_in                 =>      gt29_drpaddr_in,
        gt29_drpclk_in                  =>      gt29_drpclk_in,
        gt29_drpdi_in                   =>      gt29_drpdi_in,
        gt29_drpdo_out                  =>      gt29_drpdo_out,
        gt29_drpen_in                   =>      gt29_drpen_in,
        gt29_drprdy_out                 =>      gt29_drprdy_out,
        gt29_drpwe_in                   =>      gt29_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt29_eyescanreset_in            =>      gt29_eyescanreset_in,
        gt29_rxuserrdy_in               =>      gt29_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt29_eyescandataerror_out       =>      gt29_eyescandataerror_out,
        gt29_eyescantrigger_in          =>      gt29_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt29_rxslide_in                 =>      gt29_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt29_dmonitorout_out            =>      gt29_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt29_rxusrclk_in                =>      gt29_rxusrclk_in,
        gt29_rxusrclk2_in               =>      gt29_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt29_rxdata_out                 =>      gt29_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt29_rxdisperr_out              =>      gt29_rxdisperr_out,
        gt29_rxnotintable_out           =>      gt29_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt29_gthrxn_in                  =>      gt29_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt29_rxdlyen_in                 =>      gt29_rxdlyen_i,
        gt29_rxdlysreset_in             =>      gt29_rxdlysreset_i,
        gt29_rxdlysresetdone_out        =>      gt29_rxdlysresetdone_i,
        gt29_rxphalign_in               =>      gt29_rxphalign_i,
        gt29_rxphaligndone_out          =>      gt29_rxphaligndone_i,
        gt29_rxphalignen_in             =>      gt29_rxphalignen_i,
        gt29_rxphdlyreset_in            =>      gt29_rxphdlyreset_i,
        gt29_rxphmonitor_out            =>      gt29_rxphmonitor_out,
        gt29_rxphslipmonitor_out        =>      gt29_rxphslipmonitor_out,
        gt29_rxsyncallin_in             =>      gt29_rxsyncallin_i,
        gt29_rxsyncdone_out             =>      gt29_rxsyncdone_i,
        gt29_rxsyncin_in                =>      gt29_rxsyncin_i,
        gt29_rxsyncmode_in              =>      gt29_rxsyncmode_i,
        gt29_rxsyncout_out              =>      gt29_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt29_rxbyteisaligned_out        =>      gt29_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt29_rxlpmhfhold_in             =>      gt29_rxlpmhfhold_i,
        gt29_rxlpmlfhold_in             =>      gt29_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt29_rxmonitorout_out           =>      gt29_rxmonitorout_out,
        gt29_rxmonitorsel_in            =>      gt29_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt29_rxoutclk_out               =>      gt29_rxoutclk_i,
        gt29_rxoutclkfabric_out         =>      gt29_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt29_gtrxreset_in               =>      gt29_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt29_rxcharisk_out              =>      gt29_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt29_gthrxp_in                  =>      gt29_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt29_rxresetdone_out            =>      gt29_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt29_gttxreset_in               =>      gt29_gttxreset_i,
        gt29_txuserrdy_in               =>      gt29_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt29_txusrclk_in                =>      gt29_txusrclk_in,
        gt29_txusrclk2_in               =>      gt29_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt29_txdlyen_in                 =>      gt29_txdlyen_i,
        gt29_txdlysreset_in             =>      gt29_txdlysreset_i,
        gt29_txdlysresetdone_out        =>      gt29_txdlysresetdone_i,
        gt29_txphalign_in               =>      gt29_txphalign_i,
        gt29_txphaligndone_out          =>      gt29_txphaligndone_i,
        gt29_txphalignen_in             =>      gt29_txphalignen_i,
        gt29_txphdlyreset_in            =>      gt29_txphdlyreset_i,
        gt29_txphinit_in                =>      gt29_txphinit_i,
        gt29_txphinitdone_out           =>      gt29_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt29_txdata_in                  =>      gt29_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt29_gthtxn_out                 =>      gt29_gthtxn_out,
        gt29_gthtxp_out                 =>      gt29_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt29_txoutclk_out               =>      gt29_txoutclk_i,
        gt29_txoutclkfabric_out         =>      gt29_txoutclkfabric_out,
        gt29_txoutclkpcs_out            =>      gt29_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt29_txresetdone_out            =>      gt29_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt29_txcharisk_in               =>      gt29_txcharisk_in,


        GT30_DRP_BUSY_OUT               =>      GT30_DRP_BUSY_OUT,
        GT30_RXPMARESETDONE_OUT         =>      gt30_rxpmaresetdone_i,
        GT30_TXPMARESETDONE_OUT         =>      gt30_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT30  (X1Y34)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt30_drpaddr_in                 =>      gt30_drpaddr_in,
        gt30_drpclk_in                  =>      gt30_drpclk_in,
        gt30_drpdi_in                   =>      gt30_drpdi_in,
        gt30_drpdo_out                  =>      gt30_drpdo_out,
        gt30_drpen_in                   =>      gt30_drpen_in,
        gt30_drprdy_out                 =>      gt30_drprdy_out,
        gt30_drpwe_in                   =>      gt30_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt30_eyescanreset_in            =>      gt30_eyescanreset_in,
        gt30_rxuserrdy_in               =>      gt30_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt30_eyescandataerror_out       =>      gt30_eyescandataerror_out,
        gt30_eyescantrigger_in          =>      gt30_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt30_rxslide_in                 =>      gt30_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt30_dmonitorout_out            =>      gt30_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt30_rxusrclk_in                =>      gt30_rxusrclk_in,
        gt30_rxusrclk2_in               =>      gt30_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt30_rxdata_out                 =>      gt30_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt30_rxdisperr_out              =>      gt30_rxdisperr_out,
        gt30_rxnotintable_out           =>      gt30_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt30_gthrxn_in                  =>      gt30_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt30_rxdlyen_in                 =>      gt30_rxdlyen_i,
        gt30_rxdlysreset_in             =>      gt30_rxdlysreset_i,
        gt30_rxdlysresetdone_out        =>      gt30_rxdlysresetdone_i,
        gt30_rxphalign_in               =>      gt30_rxphalign_i,
        gt30_rxphaligndone_out          =>      gt30_rxphaligndone_i,
        gt30_rxphalignen_in             =>      gt30_rxphalignen_i,
        gt30_rxphdlyreset_in            =>      gt30_rxphdlyreset_i,
        gt30_rxphmonitor_out            =>      gt30_rxphmonitor_out,
        gt30_rxphslipmonitor_out        =>      gt30_rxphslipmonitor_out,
        gt30_rxsyncallin_in             =>      gt30_rxsyncallin_i,
        gt30_rxsyncdone_out             =>      gt30_rxsyncdone_i,
        gt30_rxsyncin_in                =>      gt30_rxsyncin_i,
        gt30_rxsyncmode_in              =>      gt30_rxsyncmode_i,
        gt30_rxsyncout_out              =>      gt30_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt30_rxbyteisaligned_out        =>      gt30_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt30_rxlpmhfhold_in             =>      gt30_rxlpmhfhold_i,
        gt30_rxlpmlfhold_in             =>      gt30_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt30_rxmonitorout_out           =>      gt30_rxmonitorout_out,
        gt30_rxmonitorsel_in            =>      gt30_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt30_rxoutclk_out               =>      gt30_rxoutclk_i,
        gt30_rxoutclkfabric_out         =>      gt30_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt30_gtrxreset_in               =>      gt30_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt30_rxcharisk_out              =>      gt30_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt30_gthrxp_in                  =>      gt30_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt30_rxresetdone_out            =>      gt30_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt30_gttxreset_in               =>      gt30_gttxreset_i,
        gt30_txuserrdy_in               =>      gt30_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt30_txusrclk_in                =>      gt30_txusrclk_in,
        gt30_txusrclk2_in               =>      gt30_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt30_txdlyen_in                 =>      gt30_txdlyen_i,
        gt30_txdlysreset_in             =>      gt30_txdlysreset_i,
        gt30_txdlysresetdone_out        =>      gt30_txdlysresetdone_i,
        gt30_txphalign_in               =>      gt30_txphalign_i,
        gt30_txphaligndone_out          =>      gt30_txphaligndone_i,
        gt30_txphalignen_in             =>      gt30_txphalignen_i,
        gt30_txphdlyreset_in            =>      gt30_txphdlyreset_i,
        gt30_txphinit_in                =>      gt30_txphinit_i,
        gt30_txphinitdone_out           =>      gt30_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt30_txdata_in                  =>      gt30_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt30_gthtxn_out                 =>      gt30_gthtxn_out,
        gt30_gthtxp_out                 =>      gt30_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt30_txoutclk_out               =>      gt30_txoutclk_i,
        gt30_txoutclkfabric_out         =>      gt30_txoutclkfabric_out,
        gt30_txoutclkpcs_out            =>      gt30_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt30_txresetdone_out            =>      gt30_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt30_txcharisk_in               =>      gt30_txcharisk_in,


        GT31_DRP_BUSY_OUT               =>      GT31_DRP_BUSY_OUT,
        GT31_RXPMARESETDONE_OUT         =>      gt31_rxpmaresetdone_i,
        GT31_TXPMARESETDONE_OUT         =>      gt31_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT31  (X1Y35)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt31_drpaddr_in                 =>      gt31_drpaddr_in,
        gt31_drpclk_in                  =>      gt31_drpclk_in,
        gt31_drpdi_in                   =>      gt31_drpdi_in,
        gt31_drpdo_out                  =>      gt31_drpdo_out,
        gt31_drpen_in                   =>      gt31_drpen_in,
        gt31_drprdy_out                 =>      gt31_drprdy_out,
        gt31_drpwe_in                   =>      gt31_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt31_eyescanreset_in            =>      gt31_eyescanreset_in,
        gt31_rxuserrdy_in               =>      gt31_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt31_eyescandataerror_out       =>      gt31_eyescandataerror_out,
        gt31_eyescantrigger_in          =>      gt31_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt31_rxslide_in                 =>      gt31_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt31_dmonitorout_out            =>      gt31_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt31_rxusrclk_in                =>      gt31_rxusrclk_in,
        gt31_rxusrclk2_in               =>      gt31_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt31_rxdata_out                 =>      gt31_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt31_rxdisperr_out              =>      gt31_rxdisperr_out,
        gt31_rxnotintable_out           =>      gt31_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt31_gthrxn_in                  =>      gt31_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt31_rxdlyen_in                 =>      gt31_rxdlyen_i,
        gt31_rxdlysreset_in             =>      gt31_rxdlysreset_i,
        gt31_rxdlysresetdone_out        =>      gt31_rxdlysresetdone_i,
        gt31_rxphalign_in               =>      gt31_rxphalign_i,
        gt31_rxphaligndone_out          =>      gt31_rxphaligndone_i,
        gt31_rxphalignen_in             =>      gt31_rxphalignen_i,
        gt31_rxphdlyreset_in            =>      gt31_rxphdlyreset_i,
        gt31_rxphmonitor_out            =>      gt31_rxphmonitor_out,
        gt31_rxphslipmonitor_out        =>      gt31_rxphslipmonitor_out,
        gt31_rxsyncallin_in             =>      gt31_rxsyncallin_i,
        gt31_rxsyncdone_out             =>      gt31_rxsyncdone_i,
        gt31_rxsyncin_in                =>      gt31_rxsyncin_i,
        gt31_rxsyncmode_in              =>      gt31_rxsyncmode_i,
        gt31_rxsyncout_out              =>      gt31_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt31_rxbyteisaligned_out        =>      gt31_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt31_rxlpmhfhold_in             =>      gt31_rxlpmhfhold_i,
        gt31_rxlpmlfhold_in             =>      gt31_rxlpmlfhold_i,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt31_rxmonitorout_out           =>      gt31_rxmonitorout_out,
        gt31_rxmonitorsel_in            =>      gt31_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt31_rxoutclk_out               =>      gt31_rxoutclk_i,
        gt31_rxoutclkfabric_out         =>      gt31_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt31_gtrxreset_in               =>      gt31_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt31_rxcharisk_out              =>      gt31_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt31_gthrxp_in                  =>      gt31_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt31_rxresetdone_out            =>      gt31_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt31_gttxreset_in               =>      gt31_gttxreset_i,
        gt31_txuserrdy_in               =>      gt31_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt31_txusrclk_in                =>      gt31_txusrclk_in,
        gt31_txusrclk2_in               =>      gt31_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt31_txdlyen_in                 =>      gt31_txdlyen_i,
        gt31_txdlysreset_in             =>      gt31_txdlysreset_i,
        gt31_txdlysresetdone_out        =>      gt31_txdlysresetdone_i,
        gt31_txphalign_in               =>      gt31_txphalign_i,
        gt31_txphaligndone_out          =>      gt31_txphaligndone_i,
        gt31_txphalignen_in             =>      gt31_txphalignen_i,
        gt31_txphdlyreset_in            =>      gt31_txphdlyreset_i,
        gt31_txphinit_in                =>      gt31_txphinit_i,
        gt31_txphinitdone_out           =>      gt31_txphinitdone_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt31_txdata_in                  =>      gt31_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt31_gthtxn_out                 =>      gt31_gthtxn_out,
        gt31_gthtxp_out                 =>      gt31_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt31_txoutclk_out               =>      gt31_txoutclk_i,
        gt31_txoutclkfabric_out         =>      gt31_txoutclkfabric_out,
        gt31_txoutclkpcs_out            =>      gt31_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt31_txresetdone_out            =>      gt31_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt31_txcharisk_in               =>      gt31_txcharisk_in,




    --____________________________COMMON PORTS________________________________
        gt0_qpllreset_in                =>      gt0_qpllreset_t,
        gt0_qplloutclk_in               =>      gt0_qplloutclk_in,
        gt0_qplloutrefclk_in            =>      gt0_qplloutrefclk_in,

    --____________________________COMMON PORTS________________________________
        gt1_qpllreset_in                =>      gt1_qpllreset_t,
        gt1_qplloutclk_in               =>      gt1_qplloutclk_in,
        gt1_qplloutrefclk_in            =>      gt1_qplloutrefclk_in,

    --____________________________COMMON PORTS________________________________
        gt2_qpllreset_in                =>      gt2_qpllreset_t,
        gt2_qplloutclk_in               =>      gt2_qplloutclk_in,
        gt2_qplloutrefclk_in            =>      gt2_qplloutrefclk_in,

    --____________________________COMMON PORTS________________________________
        gt3_qpllreset_in                =>      gt3_qpllreset_t,
        gt3_qplloutclk_in               =>      gt3_qplloutclk_in,
        gt3_qplloutrefclk_in            =>      gt3_qplloutrefclk_in,

    --____________________________COMMON PORTS________________________________
        gt4_qpllreset_in                =>      gt4_qpllreset_t,
        gt4_qplloutclk_in               =>      gt4_qplloutclk_in,
        gt4_qplloutrefclk_in            =>      gt4_qplloutrefclk_in,

    --____________________________COMMON PORTS________________________________
        gt5_qpllreset_in                =>      gt5_qpllreset_t,
        gt5_qplloutclk_in               =>      gt5_qplloutclk_in,
        gt5_qplloutrefclk_in            =>      gt5_qplloutrefclk_in,

    --____________________________COMMON PORTS________________________________
        gt6_qpllreset_in                =>      gt6_qpllreset_t,
        gt6_qplloutclk_in               =>      gt6_qplloutclk_in,
        gt6_qplloutrefclk_in            =>      gt6_qplloutrefclk_in,

    --____________________________COMMON PORTS________________________________
        gt7_qpllreset_in                =>      gt7_qpllreset_t,
        gt7_qplloutclk_in               =>      gt7_qplloutclk_in,
        gt7_qplloutrefclk_in            =>      gt7_qplloutrefclk_in
    );




GT0_TXRESETDONE_OUT                          <= gt0_txresetdone_i;
GT0_RXRESETDONE_OUT                          <= gt0_rxresetdone_i;
GT0_RXOUTCLK_OUT                             <= gt0_rxoutclk_i;
GT0_TXOUTCLK_OUT                             <= gt0_txoutclk_i;
GT1_TXRESETDONE_OUT                          <= gt1_txresetdone_i;
GT1_RXRESETDONE_OUT                          <= gt1_rxresetdone_i;
GT1_RXOUTCLK_OUT                             <= gt1_rxoutclk_i;
GT1_TXOUTCLK_OUT                             <= gt1_txoutclk_i;
GT2_TXRESETDONE_OUT                          <= gt2_txresetdone_i;
GT2_RXRESETDONE_OUT                          <= gt2_rxresetdone_i;
GT2_RXOUTCLK_OUT                             <= gt2_rxoutclk_i;
GT2_TXOUTCLK_OUT                             <= gt2_txoutclk_i;
GT3_TXRESETDONE_OUT                          <= gt3_txresetdone_i;
GT3_RXRESETDONE_OUT                          <= gt3_rxresetdone_i;
GT3_RXOUTCLK_OUT                             <= gt3_rxoutclk_i;
GT3_TXOUTCLK_OUT                             <= gt3_txoutclk_i;
GT4_TXRESETDONE_OUT                          <= gt4_txresetdone_i;
GT4_RXRESETDONE_OUT                          <= gt4_rxresetdone_i;
GT4_RXOUTCLK_OUT                             <= gt4_rxoutclk_i;
GT4_TXOUTCLK_OUT                             <= gt4_txoutclk_i;
GT5_TXRESETDONE_OUT                          <= gt5_txresetdone_i;
GT5_RXRESETDONE_OUT                          <= gt5_rxresetdone_i;
GT5_RXOUTCLK_OUT                             <= gt5_rxoutclk_i;
GT5_TXOUTCLK_OUT                             <= gt5_txoutclk_i;
GT6_TXRESETDONE_OUT                          <= gt6_txresetdone_i;
GT6_RXRESETDONE_OUT                          <= gt6_rxresetdone_i;
GT6_RXOUTCLK_OUT                             <= gt6_rxoutclk_i;
GT6_TXOUTCLK_OUT                             <= gt6_txoutclk_i;
GT7_TXRESETDONE_OUT                          <= gt7_txresetdone_i;
GT7_RXRESETDONE_OUT                          <= gt7_rxresetdone_i;
GT7_RXOUTCLK_OUT                             <= gt7_rxoutclk_i;
GT7_TXOUTCLK_OUT                             <= gt7_txoutclk_i;
GT8_TXRESETDONE_OUT                          <= gt8_txresetdone_i;
GT8_RXRESETDONE_OUT                          <= gt8_rxresetdone_i;
GT8_RXOUTCLK_OUT                             <= gt8_rxoutclk_i;
GT8_TXOUTCLK_OUT                             <= gt8_txoutclk_i;
GT9_TXRESETDONE_OUT                          <= gt9_txresetdone_i;
GT9_RXRESETDONE_OUT                          <= gt9_rxresetdone_i;
GT9_RXOUTCLK_OUT                             <= gt9_rxoutclk_i;
GT9_TXOUTCLK_OUT                             <= gt9_txoutclk_i;
GT10_TXRESETDONE_OUT                         <= gt10_txresetdone_i;
GT10_RXRESETDONE_OUT                         <= gt10_rxresetdone_i;
GT10_RXOUTCLK_OUT                            <= gt10_rxoutclk_i;
GT10_TXOUTCLK_OUT                            <= gt10_txoutclk_i;
GT11_TXRESETDONE_OUT                         <= gt11_txresetdone_i;
GT11_RXRESETDONE_OUT                         <= gt11_rxresetdone_i;
GT11_RXOUTCLK_OUT                            <= gt11_rxoutclk_i;
GT11_TXOUTCLK_OUT                            <= gt11_txoutclk_i;
GT12_TXRESETDONE_OUT                         <= gt12_txresetdone_i;
GT12_RXRESETDONE_OUT                         <= gt12_rxresetdone_i;
GT12_RXOUTCLK_OUT                            <= gt12_rxoutclk_i;
GT12_TXOUTCLK_OUT                            <= gt12_txoutclk_i;
GT13_TXRESETDONE_OUT                         <= gt13_txresetdone_i;
GT13_RXRESETDONE_OUT                         <= gt13_rxresetdone_i;
GT13_RXOUTCLK_OUT                            <= gt13_rxoutclk_i;
GT13_TXOUTCLK_OUT                            <= gt13_txoutclk_i;
GT14_TXRESETDONE_OUT                         <= gt14_txresetdone_i;
GT14_RXRESETDONE_OUT                         <= gt14_rxresetdone_i;
GT14_RXOUTCLK_OUT                            <= gt14_rxoutclk_i;
GT14_TXOUTCLK_OUT                            <= gt14_txoutclk_i;
GT15_TXRESETDONE_OUT                         <= gt15_txresetdone_i;
GT15_RXRESETDONE_OUT                         <= gt15_rxresetdone_i;
GT15_RXOUTCLK_OUT                            <= gt15_rxoutclk_i;
GT15_TXOUTCLK_OUT                            <= gt15_txoutclk_i;
GT16_TXRESETDONE_OUT                         <= gt16_txresetdone_i;
GT16_RXRESETDONE_OUT                         <= gt16_rxresetdone_i;
GT16_RXOUTCLK_OUT                            <= gt16_rxoutclk_i;
GT16_TXOUTCLK_OUT                            <= gt16_txoutclk_i;
GT17_TXRESETDONE_OUT                         <= gt17_txresetdone_i;
GT17_RXRESETDONE_OUT                         <= gt17_rxresetdone_i;
GT17_RXOUTCLK_OUT                            <= gt17_rxoutclk_i;
GT17_TXOUTCLK_OUT                            <= gt17_txoutclk_i;
GT18_TXRESETDONE_OUT                         <= gt18_txresetdone_i;
GT18_RXRESETDONE_OUT                         <= gt18_rxresetdone_i;
GT18_RXOUTCLK_OUT                            <= gt18_rxoutclk_i;
GT18_TXOUTCLK_OUT                            <= gt18_txoutclk_i;
GT19_TXRESETDONE_OUT                         <= gt19_txresetdone_i;
GT19_RXRESETDONE_OUT                         <= gt19_rxresetdone_i;
GT19_RXOUTCLK_OUT                            <= gt19_rxoutclk_i;
GT19_TXOUTCLK_OUT                            <= gt19_txoutclk_i;
GT20_TXRESETDONE_OUT                         <= gt20_txresetdone_i;
GT20_RXRESETDONE_OUT                         <= gt20_rxresetdone_i;
GT20_RXOUTCLK_OUT                            <= gt20_rxoutclk_i;
GT20_TXOUTCLK_OUT                            <= gt20_txoutclk_i;
GT21_TXRESETDONE_OUT                         <= gt21_txresetdone_i;
GT21_RXRESETDONE_OUT                         <= gt21_rxresetdone_i;
GT21_RXOUTCLK_OUT                            <= gt21_rxoutclk_i;
GT21_TXOUTCLK_OUT                            <= gt21_txoutclk_i;
GT22_TXRESETDONE_OUT                         <= gt22_txresetdone_i;
GT22_RXRESETDONE_OUT                         <= gt22_rxresetdone_i;
GT22_RXOUTCLK_OUT                            <= gt22_rxoutclk_i;
GT22_TXOUTCLK_OUT                            <= gt22_txoutclk_i;
GT23_TXRESETDONE_OUT                         <= gt23_txresetdone_i;
GT23_RXRESETDONE_OUT                         <= gt23_rxresetdone_i;
GT23_RXOUTCLK_OUT                            <= gt23_rxoutclk_i;
GT23_TXOUTCLK_OUT                            <= gt23_txoutclk_i;
GT24_TXRESETDONE_OUT                         <= gt24_txresetdone_i;
GT24_RXRESETDONE_OUT                         <= gt24_rxresetdone_i;
GT24_RXOUTCLK_OUT                            <= gt24_rxoutclk_i;
GT24_TXOUTCLK_OUT                            <= gt24_txoutclk_i;
GT25_TXRESETDONE_OUT                         <= gt25_txresetdone_i;
GT25_RXRESETDONE_OUT                         <= gt25_rxresetdone_i;
GT25_RXOUTCLK_OUT                            <= gt25_rxoutclk_i;
GT25_TXOUTCLK_OUT                            <= gt25_txoutclk_i;
GT26_TXRESETDONE_OUT                         <= gt26_txresetdone_i;
GT26_RXRESETDONE_OUT                         <= gt26_rxresetdone_i;
GT26_RXOUTCLK_OUT                            <= gt26_rxoutclk_i;
GT26_TXOUTCLK_OUT                            <= gt26_txoutclk_i;
GT27_TXRESETDONE_OUT                         <= gt27_txresetdone_i;
GT27_RXRESETDONE_OUT                         <= gt27_rxresetdone_i;
GT27_RXOUTCLK_OUT                            <= gt27_rxoutclk_i;
GT27_TXOUTCLK_OUT                            <= gt27_txoutclk_i;
GT28_TXRESETDONE_OUT                         <= gt28_txresetdone_i;
GT28_RXRESETDONE_OUT                         <= gt28_rxresetdone_i;
GT28_RXOUTCLK_OUT                            <= gt28_rxoutclk_i;
GT28_TXOUTCLK_OUT                            <= gt28_txoutclk_i;
GT29_TXRESETDONE_OUT                         <= gt29_txresetdone_i;
GT29_RXRESETDONE_OUT                         <= gt29_rxresetdone_i;
GT29_RXOUTCLK_OUT                            <= gt29_rxoutclk_i;
GT29_TXOUTCLK_OUT                            <= gt29_txoutclk_i;
GT30_TXRESETDONE_OUT                         <= gt30_txresetdone_i;
GT30_RXRESETDONE_OUT                         <= gt30_rxresetdone_i;
GT30_RXOUTCLK_OUT                            <= gt30_rxoutclk_i;
GT30_TXOUTCLK_OUT                            <= gt30_txoutclk_i;
GT31_TXRESETDONE_OUT                         <= gt31_txresetdone_i;
GT31_RXRESETDONE_OUT                         <= gt31_rxresetdone_i;
GT31_RXOUTCLK_OUT                            <= gt31_rxoutclk_i;
GT31_TXOUTCLK_OUT                            <= gt31_txoutclk_i;
    GT0_QPLLRESET_OUT                            <= gt0_qpllreset_t;
    GT1_QPLLRESET_OUT                            <= gt1_qpllreset_t;
    GT2_QPLLRESET_OUT                            <= gt2_qpllreset_t;
    GT3_QPLLRESET_OUT                            <= gt3_qpllreset_t;
    GT4_QPLLRESET_OUT                            <= gt4_qpllreset_t;
    GT5_QPLLRESET_OUT                            <= gt5_qpllreset_t;
    GT6_QPLLRESET_OUT                            <= gt6_qpllreset_t;
    GT7_QPLLRESET_OUT                            <= gt7_qpllreset_t;

chipscope : if EXAMPLE_USE_CHIPSCOPE = 1 generate
    gt0_gttxreset_i                              <= GT0_GTTXRESET_IN or gt0_gttxreset_t;
    gt0_gtrxreset_i                              <= GT0_GTRXRESET_IN or gt0_gtrxreset_t;
    gt0_txuserrdy_i                              <= GT0_TXUSERRDY_IN and gt0_txuserrdy_t;
    gt0_rxuserrdy_i                              <= GT0_RXUSERRDY_IN and gt0_rxuserrdy_t;
    gt1_gttxreset_i                              <= GT1_GTTXRESET_IN or gt1_gttxreset_t;
    gt1_gtrxreset_i                              <= GT1_GTRXRESET_IN or gt1_gtrxreset_t;
    gt1_txuserrdy_i                              <= GT1_TXUSERRDY_IN and gt1_txuserrdy_t;
    gt1_rxuserrdy_i                              <= GT1_RXUSERRDY_IN and gt1_rxuserrdy_t;
    gt2_gttxreset_i                              <= GT2_GTTXRESET_IN or gt2_gttxreset_t;
    gt2_gtrxreset_i                              <= GT2_GTRXRESET_IN or gt2_gtrxreset_t;
    gt2_txuserrdy_i                              <= GT2_TXUSERRDY_IN and gt2_txuserrdy_t;
    gt2_rxuserrdy_i                              <= GT2_RXUSERRDY_IN and gt2_rxuserrdy_t;
    gt3_gttxreset_i                              <= GT3_GTTXRESET_IN or gt3_gttxreset_t;
    gt3_gtrxreset_i                              <= GT3_GTRXRESET_IN or gt3_gtrxreset_t;
    gt3_txuserrdy_i                              <= GT3_TXUSERRDY_IN and gt3_txuserrdy_t;
    gt3_rxuserrdy_i                              <= GT3_RXUSERRDY_IN and gt3_rxuserrdy_t;
    gt4_gttxreset_i                              <= GT4_GTTXRESET_IN or gt4_gttxreset_t;
    gt4_gtrxreset_i                              <= GT4_GTRXRESET_IN or gt4_gtrxreset_t;
    gt4_txuserrdy_i                              <= GT4_TXUSERRDY_IN and gt4_txuserrdy_t;
    gt4_rxuserrdy_i                              <= GT4_RXUSERRDY_IN and gt4_rxuserrdy_t;
    gt5_gttxreset_i                              <= GT5_GTTXRESET_IN or gt5_gttxreset_t;
    gt5_gtrxreset_i                              <= GT5_GTRXRESET_IN or gt5_gtrxreset_t;
    gt5_txuserrdy_i                              <= GT5_TXUSERRDY_IN and gt5_txuserrdy_t;
    gt5_rxuserrdy_i                              <= GT5_RXUSERRDY_IN and gt5_rxuserrdy_t;
    gt6_gttxreset_i                              <= GT6_GTTXRESET_IN or gt6_gttxreset_t;
    gt6_gtrxreset_i                              <= GT6_GTRXRESET_IN or gt6_gtrxreset_t;
    gt6_txuserrdy_i                              <= GT6_TXUSERRDY_IN and gt6_txuserrdy_t;
    gt6_rxuserrdy_i                              <= GT6_RXUSERRDY_IN and gt6_rxuserrdy_t;
    gt7_gttxreset_i                              <= GT7_GTTXRESET_IN or gt7_gttxreset_t;
    gt7_gtrxreset_i                              <= GT7_GTRXRESET_IN or gt7_gtrxreset_t;
    gt7_txuserrdy_i                              <= GT7_TXUSERRDY_IN and gt7_txuserrdy_t;
    gt7_rxuserrdy_i                              <= GT7_RXUSERRDY_IN and gt7_rxuserrdy_t;
    gt8_gttxreset_i                              <= GT8_GTTXRESET_IN or gt8_gttxreset_t;
    gt8_gtrxreset_i                              <= GT8_GTRXRESET_IN or gt8_gtrxreset_t;
    gt8_txuserrdy_i                              <= GT8_TXUSERRDY_IN and gt8_txuserrdy_t;
    gt8_rxuserrdy_i                              <= GT8_RXUSERRDY_IN and gt8_rxuserrdy_t;
    gt9_gttxreset_i                              <= GT9_GTTXRESET_IN or gt9_gttxreset_t;
    gt9_gtrxreset_i                              <= GT9_GTRXRESET_IN or gt9_gtrxreset_t;
    gt9_txuserrdy_i                              <= GT9_TXUSERRDY_IN and gt9_txuserrdy_t;
    gt9_rxuserrdy_i                              <= GT9_RXUSERRDY_IN and gt9_rxuserrdy_t;
    gt10_gttxreset_i                             <= GT10_GTTXRESET_IN or gt10_gttxreset_t;
    gt10_gtrxreset_i                             <= GT10_GTRXRESET_IN or gt10_gtrxreset_t;
    gt10_txuserrdy_i                             <= GT10_TXUSERRDY_IN and gt10_txuserrdy_t;
    gt10_rxuserrdy_i                             <= GT10_RXUSERRDY_IN and gt10_rxuserrdy_t;
    gt11_gttxreset_i                             <= GT11_GTTXRESET_IN or gt11_gttxreset_t;
    gt11_gtrxreset_i                             <= GT11_GTRXRESET_IN or gt11_gtrxreset_t;
    gt11_txuserrdy_i                             <= GT11_TXUSERRDY_IN and gt11_txuserrdy_t;
    gt11_rxuserrdy_i                             <= GT11_RXUSERRDY_IN and gt11_rxuserrdy_t;
    gt12_gttxreset_i                             <= GT12_GTTXRESET_IN or gt12_gttxreset_t;
    gt12_gtrxreset_i                             <= GT12_GTRXRESET_IN or gt12_gtrxreset_t;
    gt12_txuserrdy_i                             <= GT12_TXUSERRDY_IN and gt12_txuserrdy_t;
    gt12_rxuserrdy_i                             <= GT12_RXUSERRDY_IN and gt12_rxuserrdy_t;
    gt13_gttxreset_i                             <= GT13_GTTXRESET_IN or gt13_gttxreset_t;
    gt13_gtrxreset_i                             <= GT13_GTRXRESET_IN or gt13_gtrxreset_t;
    gt13_txuserrdy_i                             <= GT13_TXUSERRDY_IN and gt13_txuserrdy_t;
    gt13_rxuserrdy_i                             <= GT13_RXUSERRDY_IN and gt13_rxuserrdy_t;
    gt14_gttxreset_i                             <= GT14_GTTXRESET_IN or gt14_gttxreset_t;
    gt14_gtrxreset_i                             <= GT14_GTRXRESET_IN or gt14_gtrxreset_t;
    gt14_txuserrdy_i                             <= GT14_TXUSERRDY_IN and gt14_txuserrdy_t;
    gt14_rxuserrdy_i                             <= GT14_RXUSERRDY_IN and gt14_rxuserrdy_t;
    gt15_gttxreset_i                             <= GT15_GTTXRESET_IN or gt15_gttxreset_t;
    gt15_gtrxreset_i                             <= GT15_GTRXRESET_IN or gt15_gtrxreset_t;
    gt15_txuserrdy_i                             <= GT15_TXUSERRDY_IN and gt15_txuserrdy_t;
    gt15_rxuserrdy_i                             <= GT15_RXUSERRDY_IN and gt15_rxuserrdy_t;
    gt16_gttxreset_i                             <= GT16_GTTXRESET_IN or gt16_gttxreset_t;
    gt16_gtrxreset_i                             <= GT16_GTRXRESET_IN or gt16_gtrxreset_t;
    gt16_txuserrdy_i                             <= GT16_TXUSERRDY_IN and gt16_txuserrdy_t;
    gt16_rxuserrdy_i                             <= GT16_RXUSERRDY_IN and gt16_rxuserrdy_t;
    gt17_gttxreset_i                             <= GT17_GTTXRESET_IN or gt17_gttxreset_t;
    gt17_gtrxreset_i                             <= GT17_GTRXRESET_IN or gt17_gtrxreset_t;
    gt17_txuserrdy_i                             <= GT17_TXUSERRDY_IN and gt17_txuserrdy_t;
    gt17_rxuserrdy_i                             <= GT17_RXUSERRDY_IN and gt17_rxuserrdy_t;
    gt18_gttxreset_i                             <= GT18_GTTXRESET_IN or gt18_gttxreset_t;
    gt18_gtrxreset_i                             <= GT18_GTRXRESET_IN or gt18_gtrxreset_t;
    gt18_txuserrdy_i                             <= GT18_TXUSERRDY_IN and gt18_txuserrdy_t;
    gt18_rxuserrdy_i                             <= GT18_RXUSERRDY_IN and gt18_rxuserrdy_t;
    gt19_gttxreset_i                             <= GT19_GTTXRESET_IN or gt19_gttxreset_t;
    gt19_gtrxreset_i                             <= GT19_GTRXRESET_IN or gt19_gtrxreset_t;
    gt19_txuserrdy_i                             <= GT19_TXUSERRDY_IN and gt19_txuserrdy_t;
    gt19_rxuserrdy_i                             <= GT19_RXUSERRDY_IN and gt19_rxuserrdy_t;
    gt20_gttxreset_i                             <= GT20_GTTXRESET_IN or gt20_gttxreset_t;
    gt20_gtrxreset_i                             <= GT20_GTRXRESET_IN or gt20_gtrxreset_t;
    gt20_txuserrdy_i                             <= GT20_TXUSERRDY_IN and gt20_txuserrdy_t;
    gt20_rxuserrdy_i                             <= GT20_RXUSERRDY_IN and gt20_rxuserrdy_t;
    gt21_gttxreset_i                             <= GT21_GTTXRESET_IN or gt21_gttxreset_t;
    gt21_gtrxreset_i                             <= GT21_GTRXRESET_IN or gt21_gtrxreset_t;
    gt21_txuserrdy_i                             <= GT21_TXUSERRDY_IN and gt21_txuserrdy_t;
    gt21_rxuserrdy_i                             <= GT21_RXUSERRDY_IN and gt21_rxuserrdy_t;
    gt22_gttxreset_i                             <= GT22_GTTXRESET_IN or gt22_gttxreset_t;
    gt22_gtrxreset_i                             <= GT22_GTRXRESET_IN or gt22_gtrxreset_t;
    gt22_txuserrdy_i                             <= GT22_TXUSERRDY_IN and gt22_txuserrdy_t;
    gt22_rxuserrdy_i                             <= GT22_RXUSERRDY_IN and gt22_rxuserrdy_t;
    gt23_gttxreset_i                             <= GT23_GTTXRESET_IN or gt23_gttxreset_t;
    gt23_gtrxreset_i                             <= GT23_GTRXRESET_IN or gt23_gtrxreset_t;
    gt23_txuserrdy_i                             <= GT23_TXUSERRDY_IN and gt23_txuserrdy_t;
    gt23_rxuserrdy_i                             <= GT23_RXUSERRDY_IN and gt23_rxuserrdy_t;
    gt24_gttxreset_i                             <= GT24_GTTXRESET_IN or gt24_gttxreset_t;
    gt24_gtrxreset_i                             <= GT24_GTRXRESET_IN or gt24_gtrxreset_t;
    gt24_txuserrdy_i                             <= GT24_TXUSERRDY_IN and gt24_txuserrdy_t;
    gt24_rxuserrdy_i                             <= GT24_RXUSERRDY_IN and gt24_rxuserrdy_t;
    gt25_gttxreset_i                             <= GT25_GTTXRESET_IN or gt25_gttxreset_t;
    gt25_gtrxreset_i                             <= GT25_GTRXRESET_IN or gt25_gtrxreset_t;
    gt25_txuserrdy_i                             <= GT25_TXUSERRDY_IN and gt25_txuserrdy_t;
    gt25_rxuserrdy_i                             <= GT25_RXUSERRDY_IN and gt25_rxuserrdy_t;
    gt26_gttxreset_i                             <= GT26_GTTXRESET_IN or gt26_gttxreset_t;
    gt26_gtrxreset_i                             <= GT26_GTRXRESET_IN or gt26_gtrxreset_t;
    gt26_txuserrdy_i                             <= GT26_TXUSERRDY_IN and gt26_txuserrdy_t;
    gt26_rxuserrdy_i                             <= GT26_RXUSERRDY_IN and gt26_rxuserrdy_t;
    gt27_gttxreset_i                             <= GT27_GTTXRESET_IN or gt27_gttxreset_t;
    gt27_gtrxreset_i                             <= GT27_GTRXRESET_IN or gt27_gtrxreset_t;
    gt27_txuserrdy_i                             <= GT27_TXUSERRDY_IN and gt27_txuserrdy_t;
    gt27_rxuserrdy_i                             <= GT27_RXUSERRDY_IN and gt27_rxuserrdy_t;
    gt28_gttxreset_i                             <= GT28_GTTXRESET_IN or gt28_gttxreset_t;
    gt28_gtrxreset_i                             <= GT28_GTRXRESET_IN or gt28_gtrxreset_t;
    gt28_txuserrdy_i                             <= GT28_TXUSERRDY_IN and gt28_txuserrdy_t;
    gt28_rxuserrdy_i                             <= GT28_RXUSERRDY_IN and gt28_rxuserrdy_t;
    gt29_gttxreset_i                             <= GT29_GTTXRESET_IN or gt29_gttxreset_t;
    gt29_gtrxreset_i                             <= GT29_GTRXRESET_IN or gt29_gtrxreset_t;
    gt29_txuserrdy_i                             <= GT29_TXUSERRDY_IN and gt29_txuserrdy_t;
    gt29_rxuserrdy_i                             <= GT29_RXUSERRDY_IN and gt29_rxuserrdy_t;
    gt30_gttxreset_i                             <= GT30_GTTXRESET_IN or gt30_gttxreset_t;
    gt30_gtrxreset_i                             <= GT30_GTRXRESET_IN or gt30_gtrxreset_t;
    gt30_txuserrdy_i                             <= GT30_TXUSERRDY_IN and gt30_txuserrdy_t;
    gt30_rxuserrdy_i                             <= GT30_RXUSERRDY_IN and gt30_rxuserrdy_t;
    gt31_gttxreset_i                             <= GT31_GTTXRESET_IN or gt31_gttxreset_t;
    gt31_gtrxreset_i                             <= GT31_GTRXRESET_IN or gt31_gtrxreset_t;
    gt31_txuserrdy_i                             <= GT31_TXUSERRDY_IN and gt31_txuserrdy_t;
    gt31_rxuserrdy_i                             <= GT31_RXUSERRDY_IN and gt31_rxuserrdy_t;
end generate chipscope;

no_chipscope : if EXAMPLE_USE_CHIPSCOPE = 0 generate
gt0_gttxreset_i                              <= gt0_gttxreset_t;
gt0_gtrxreset_i                              <= gt0_gtrxreset_t;
gt0_txuserrdy_i                              <= gt0_txuserrdy_t;
gt0_rxuserrdy_i                              <= gt0_rxuserrdy_t;
gt1_gttxreset_i                              <= gt1_gttxreset_t;
gt1_gtrxreset_i                              <= gt1_gtrxreset_t;
gt1_txuserrdy_i                              <= gt1_txuserrdy_t;
gt1_rxuserrdy_i                              <= gt1_rxuserrdy_t;
gt2_gttxreset_i                              <= gt2_gttxreset_t;
gt2_gtrxreset_i                              <= gt2_gtrxreset_t;
gt2_txuserrdy_i                              <= gt2_txuserrdy_t;
gt2_rxuserrdy_i                              <= gt2_rxuserrdy_t;
gt3_gttxreset_i                              <= gt3_gttxreset_t;
gt3_gtrxreset_i                              <= gt3_gtrxreset_t;
gt3_txuserrdy_i                              <= gt3_txuserrdy_t;
gt3_rxuserrdy_i                              <= gt3_rxuserrdy_t;
gt4_gttxreset_i                              <= gt4_gttxreset_t;
gt4_gtrxreset_i                              <= gt4_gtrxreset_t;
gt4_txuserrdy_i                              <= gt4_txuserrdy_t;
gt4_rxuserrdy_i                              <= gt4_rxuserrdy_t;
gt5_gttxreset_i                              <= gt5_gttxreset_t;
gt5_gtrxreset_i                              <= gt5_gtrxreset_t;
gt5_txuserrdy_i                              <= gt5_txuserrdy_t;
gt5_rxuserrdy_i                              <= gt5_rxuserrdy_t;
gt6_gttxreset_i                              <= gt6_gttxreset_t;
gt6_gtrxreset_i                              <= gt6_gtrxreset_t;
gt6_txuserrdy_i                              <= gt6_txuserrdy_t;
gt6_rxuserrdy_i                              <= gt6_rxuserrdy_t;
gt7_gttxreset_i                              <= gt7_gttxreset_t;
gt7_gtrxreset_i                              <= gt7_gtrxreset_t;
gt7_txuserrdy_i                              <= gt7_txuserrdy_t;
gt7_rxuserrdy_i                              <= gt7_rxuserrdy_t;
gt8_gttxreset_i                              <= gt8_gttxreset_t;
gt8_gtrxreset_i                              <= gt8_gtrxreset_t;
gt8_txuserrdy_i                              <= gt8_txuserrdy_t;
gt8_rxuserrdy_i                              <= gt8_rxuserrdy_t;
gt9_gttxreset_i                              <= gt9_gttxreset_t;
gt9_gtrxreset_i                              <= gt9_gtrxreset_t;
gt9_txuserrdy_i                              <= gt9_txuserrdy_t;
gt9_rxuserrdy_i                              <= gt9_rxuserrdy_t;
gt10_gttxreset_i                             <= gt10_gttxreset_t;
gt10_gtrxreset_i                             <= gt10_gtrxreset_t;
gt10_txuserrdy_i                             <= gt10_txuserrdy_t;
gt10_rxuserrdy_i                             <= gt10_rxuserrdy_t;
gt11_gttxreset_i                             <= gt11_gttxreset_t;
gt11_gtrxreset_i                             <= gt11_gtrxreset_t;
gt11_txuserrdy_i                             <= gt11_txuserrdy_t;
gt11_rxuserrdy_i                             <= gt11_rxuserrdy_t;
gt12_gttxreset_i                             <= gt12_gttxreset_t;
gt12_gtrxreset_i                             <= gt12_gtrxreset_t;
gt12_txuserrdy_i                             <= gt12_txuserrdy_t;
gt12_rxuserrdy_i                             <= gt12_rxuserrdy_t;
gt13_gttxreset_i                             <= gt13_gttxreset_t;
gt13_gtrxreset_i                             <= gt13_gtrxreset_t;
gt13_txuserrdy_i                             <= gt13_txuserrdy_t;
gt13_rxuserrdy_i                             <= gt13_rxuserrdy_t;
gt14_gttxreset_i                             <= gt14_gttxreset_t;
gt14_gtrxreset_i                             <= gt14_gtrxreset_t;
gt14_txuserrdy_i                             <= gt14_txuserrdy_t;
gt14_rxuserrdy_i                             <= gt14_rxuserrdy_t;
gt15_gttxreset_i                             <= gt15_gttxreset_t;
gt15_gtrxreset_i                             <= gt15_gtrxreset_t;
gt15_txuserrdy_i                             <= gt15_txuserrdy_t;
gt15_rxuserrdy_i                             <= gt15_rxuserrdy_t;
gt16_gttxreset_i                             <= gt16_gttxreset_t;
gt16_gtrxreset_i                             <= gt16_gtrxreset_t;
gt16_txuserrdy_i                             <= gt16_txuserrdy_t;
gt16_rxuserrdy_i                             <= gt16_rxuserrdy_t;
gt17_gttxreset_i                             <= gt17_gttxreset_t;
gt17_gtrxreset_i                             <= gt17_gtrxreset_t;
gt17_txuserrdy_i                             <= gt17_txuserrdy_t;
gt17_rxuserrdy_i                             <= gt17_rxuserrdy_t;
gt18_gttxreset_i                             <= gt18_gttxreset_t;
gt18_gtrxreset_i                             <= gt18_gtrxreset_t;
gt18_txuserrdy_i                             <= gt18_txuserrdy_t;
gt18_rxuserrdy_i                             <= gt18_rxuserrdy_t;
gt19_gttxreset_i                             <= gt19_gttxreset_t;
gt19_gtrxreset_i                             <= gt19_gtrxreset_t;
gt19_txuserrdy_i                             <= gt19_txuserrdy_t;
gt19_rxuserrdy_i                             <= gt19_rxuserrdy_t;
gt20_gttxreset_i                             <= gt20_gttxreset_t;
gt20_gtrxreset_i                             <= gt20_gtrxreset_t;
gt20_txuserrdy_i                             <= gt20_txuserrdy_t;
gt20_rxuserrdy_i                             <= gt20_rxuserrdy_t;
gt21_gttxreset_i                             <= gt21_gttxreset_t;
gt21_gtrxreset_i                             <= gt21_gtrxreset_t;
gt21_txuserrdy_i                             <= gt21_txuserrdy_t;
gt21_rxuserrdy_i                             <= gt21_rxuserrdy_t;
gt22_gttxreset_i                             <= gt22_gttxreset_t;
gt22_gtrxreset_i                             <= gt22_gtrxreset_t;
gt22_txuserrdy_i                             <= gt22_txuserrdy_t;
gt22_rxuserrdy_i                             <= gt22_rxuserrdy_t;
gt23_gttxreset_i                             <= gt23_gttxreset_t;
gt23_gtrxreset_i                             <= gt23_gtrxreset_t;
gt23_txuserrdy_i                             <= gt23_txuserrdy_t;
gt23_rxuserrdy_i                             <= gt23_rxuserrdy_t;
gt24_gttxreset_i                             <= gt24_gttxreset_t;
gt24_gtrxreset_i                             <= gt24_gtrxreset_t;
gt24_txuserrdy_i                             <= gt24_txuserrdy_t;
gt24_rxuserrdy_i                             <= gt24_rxuserrdy_t;
gt25_gttxreset_i                             <= gt25_gttxreset_t;
gt25_gtrxreset_i                             <= gt25_gtrxreset_t;
gt25_txuserrdy_i                             <= gt25_txuserrdy_t;
gt25_rxuserrdy_i                             <= gt25_rxuserrdy_t;
gt26_gttxreset_i                             <= gt26_gttxreset_t;
gt26_gtrxreset_i                             <= gt26_gtrxreset_t;
gt26_txuserrdy_i                             <= gt26_txuserrdy_t;
gt26_rxuserrdy_i                             <= gt26_rxuserrdy_t;
gt27_gttxreset_i                             <= gt27_gttxreset_t;
gt27_gtrxreset_i                             <= gt27_gtrxreset_t;
gt27_txuserrdy_i                             <= gt27_txuserrdy_t;
gt27_rxuserrdy_i                             <= gt27_rxuserrdy_t;
gt28_gttxreset_i                             <= gt28_gttxreset_t;
gt28_gtrxreset_i                             <= gt28_gtrxreset_t;
gt28_txuserrdy_i                             <= gt28_txuserrdy_t;
gt28_rxuserrdy_i                             <= gt28_rxuserrdy_t;
gt29_gttxreset_i                             <= gt29_gttxreset_t;
gt29_gtrxreset_i                             <= gt29_gtrxreset_t;
gt29_txuserrdy_i                             <= gt29_txuserrdy_t;
gt29_rxuserrdy_i                             <= gt29_rxuserrdy_t;
gt30_gttxreset_i                             <= gt30_gttxreset_t;
gt30_gtrxreset_i                             <= gt30_gtrxreset_t;
gt30_txuserrdy_i                             <= gt30_txuserrdy_t;
gt30_rxuserrdy_i                             <= gt30_rxuserrdy_t;
gt31_gttxreset_i                             <= gt31_gttxreset_t;
gt31_gtrxreset_i                             <= gt31_gtrxreset_t;
gt31_txuserrdy_i                             <= gt31_txuserrdy_t;
gt31_rxuserrdy_i                             <= gt31_rxuserrdy_t;
end generate no_chipscope;


gt0_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT0_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT0_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT0_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt0_txresetdone_i,
        MMCM_LOCK                       =>      GT0_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt0_gttxreset_t,
        MMCM_RESET                      =>      GT0_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      gt0_qpllreset_t,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT0_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt0_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt0_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt0_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt1_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT1_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT0_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT0_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt1_txresetdone_i,
        MMCM_LOCK                       =>      GT1_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt1_gttxreset_t,
        MMCM_RESET                      =>      GT1_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT1_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt1_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt1_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt1_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt2_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT2_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT0_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT0_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt2_txresetdone_i,
        MMCM_LOCK                       =>      GT2_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt2_gttxreset_t,
        MMCM_RESET                      =>      GT2_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT2_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt2_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt2_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt2_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt3_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT3_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT0_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT0_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt3_txresetdone_i,
        MMCM_LOCK                       =>      GT3_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt3_gttxreset_t,
        MMCM_RESET                      =>      GT3_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT3_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt3_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt3_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt3_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt4_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT4_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT1_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT1_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt4_txresetdone_i,
        MMCM_LOCK                       =>      GT4_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt4_gttxreset_t,
        MMCM_RESET                      =>      GT4_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      gt1_qpllreset_t,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT4_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt4_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt4_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt4_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt5_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT5_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT1_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT1_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt5_txresetdone_i,
        MMCM_LOCK                       =>      GT5_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt5_gttxreset_t,
        MMCM_RESET                      =>      GT5_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT5_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt5_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt5_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt5_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt6_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT6_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT1_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT1_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt6_txresetdone_i,
        MMCM_LOCK                       =>      GT6_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt6_gttxreset_t,
        MMCM_RESET                      =>      GT6_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT6_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt6_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt6_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt6_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt7_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT7_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT1_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT1_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt7_txresetdone_i,
        MMCM_LOCK                       =>      GT7_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt7_gttxreset_t,
        MMCM_RESET                      =>      GT7_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT7_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt7_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt7_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt7_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt8_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT8_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT2_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT2_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt8_txresetdone_i,
        MMCM_LOCK                       =>      GT8_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt8_gttxreset_t,
        MMCM_RESET                      =>      GT8_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      gt2_qpllreset_t,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT8_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt8_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt8_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt8_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt9_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT9_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT2_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT2_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt9_txresetdone_i,
        MMCM_LOCK                       =>      GT9_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt9_gttxreset_t,
        MMCM_RESET                      =>      GT9_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT9_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt9_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt9_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt9_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt10_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT10_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT2_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT2_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt10_txresetdone_i,
        MMCM_LOCK                       =>      GT10_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt10_gttxreset_t,
        MMCM_RESET                      =>      GT10_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT10_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt10_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt10_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt10_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt11_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT11_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT2_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT2_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt11_txresetdone_i,
        MMCM_LOCK                       =>      GT11_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt11_gttxreset_t,
        MMCM_RESET                      =>      GT11_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT11_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt11_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt11_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt11_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt12_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT12_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT3_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT3_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt12_txresetdone_i,
        MMCM_LOCK                       =>      GT12_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt12_gttxreset_t,
        MMCM_RESET                      =>      GT12_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      gt3_qpllreset_t,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT12_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt12_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt12_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt12_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt12_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt13_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT13_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT3_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT3_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt13_txresetdone_i,
        MMCM_LOCK                       =>      GT13_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt13_gttxreset_t,
        MMCM_RESET                      =>      GT13_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT13_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt13_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt13_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt13_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt12_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt14_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT14_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT3_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT3_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt14_txresetdone_i,
        MMCM_LOCK                       =>      GT14_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt14_gttxreset_t,
        MMCM_RESET                      =>      GT14_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT14_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt14_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt14_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt14_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt12_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt15_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT15_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT3_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT3_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt15_txresetdone_i,
        MMCM_LOCK                       =>      GT15_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt15_gttxreset_t,
        MMCM_RESET                      =>      GT15_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT15_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt15_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt15_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt15_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt12_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt16_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT16_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT4_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT4_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt16_txresetdone_i,
        MMCM_LOCK                       =>      GT16_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt16_gttxreset_t,
        MMCM_RESET                      =>      GT16_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      gt4_qpllreset_t,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT16_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt16_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt16_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt16_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt12_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt17_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT17_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT4_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT4_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt17_txresetdone_i,
        MMCM_LOCK                       =>      GT17_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt17_gttxreset_t,
        MMCM_RESET                      =>      GT17_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT17_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt17_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt17_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt17_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt12_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt18_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT18_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT4_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT4_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt18_txresetdone_i,
        MMCM_LOCK                       =>      GT18_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt18_gttxreset_t,
        MMCM_RESET                      =>      GT18_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT18_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt18_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt18_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt18_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt12_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt19_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT19_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT4_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT4_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt19_txresetdone_i,
        MMCM_LOCK                       =>      GT19_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt19_gttxreset_t,
        MMCM_RESET                      =>      GT19_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT19_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt19_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt19_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt19_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt12_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt20_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT20_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT5_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT5_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt20_txresetdone_i,
        MMCM_LOCK                       =>      GT20_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt20_gttxreset_t,
        MMCM_RESET                      =>      GT20_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      gt5_qpllreset_t,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT20_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt20_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt20_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt20_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt12_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt21_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT21_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT5_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT5_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt21_txresetdone_i,
        MMCM_LOCK                       =>      GT21_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt21_gttxreset_t,
        MMCM_RESET                      =>      GT21_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT21_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt21_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt21_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt21_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt12_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt22_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT22_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT5_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT5_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt22_txresetdone_i,
        MMCM_LOCK                       =>      GT22_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt22_gttxreset_t,
        MMCM_RESET                      =>      GT22_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT22_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt22_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt22_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt22_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt12_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt23_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT23_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT5_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT5_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt23_txresetdone_i,
        MMCM_LOCK                       =>      GT23_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt23_gttxreset_t,
        MMCM_RESET                      =>      GT23_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT23_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt23_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt23_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt23_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt12_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt24_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT24_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT6_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT6_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt24_txresetdone_i,
        MMCM_LOCK                       =>      GT24_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt24_gttxreset_t,
        MMCM_RESET                      =>      GT24_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      gt6_qpllreset_t,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT24_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt24_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt24_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt24_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt24_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt25_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT25_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT6_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT6_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt25_txresetdone_i,
        MMCM_LOCK                       =>      GT25_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt25_gttxreset_t,
        MMCM_RESET                      =>      GT25_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT25_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt25_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt25_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt25_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt24_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt26_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT26_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT6_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT6_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt26_txresetdone_i,
        MMCM_LOCK                       =>      GT26_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt26_gttxreset_t,
        MMCM_RESET                      =>      GT26_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT26_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt26_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt26_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt26_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt24_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt27_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT27_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT6_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT6_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt27_txresetdone_i,
        MMCM_LOCK                       =>      GT27_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt27_gttxreset_t,
        MMCM_RESET                      =>      GT27_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT27_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt27_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt27_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt27_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt24_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt28_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT28_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT7_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT7_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt28_txresetdone_i,
        MMCM_LOCK                       =>      GT28_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt28_gttxreset_t,
        MMCM_RESET                      =>      GT28_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      gt7_qpllreset_t,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT28_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt28_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt28_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt28_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt24_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt29_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT29_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT7_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT7_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt29_txresetdone_i,
        MMCM_LOCK                       =>      GT29_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt29_gttxreset_t,
        MMCM_RESET                      =>      GT29_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT29_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt29_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt29_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt29_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt24_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt30_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT30_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT7_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT7_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt30_txresetdone_i,
        MMCM_LOCK                       =>      GT30_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt30_gttxreset_t,
        MMCM_RESET                      =>      GT30_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT30_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt30_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt30_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt30_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt24_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt31_txresetfsm_i:  gtwizard_0_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT31_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_TX_IN,
        QPLLREFCLKLOST                  =>      GT7_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT7_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt31_txresetdone_i,
        MMCM_LOCK                       =>      GT31_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt31_gttxreset_t,
        MMCM_RESET                      =>      GT31_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT31_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt31_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt31_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt31_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt24_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );






    rxout0_i : BUFG
    port map
    (
        I                               =>      gt0_rxoutclk_i,
        O                               =>      gt0_rxoutclk_i2
    );
    rxout12_i : BUFG
    port map
    (
        I                               =>      gt12_rxoutclk_i,
        O                               =>      gt12_rxoutclk_i2
    );
    rxout24_i : BUFG
    port map
    (
        I                               =>      gt24_rxoutclk_i,
        O                               =>      gt24_rxoutclk_i2
    );
   gt0_txoutclk_i2 <='0';
   gt12_txoutclk_i2 <='0';
   gt24_txoutclk_i2 <='0';


gt0_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT0_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT0_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT0_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt0_rxresetdone_i,
        MMCM_LOCK                       =>      GT0_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT0_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt0_gtrxreset_t,
        MMCM_RESET                      =>      GT0_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT0_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt0_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt0_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt0_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt0_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt0_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt0_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt0_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt1_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT1_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT0_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT0_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt1_rxresetdone_i,
        MMCM_LOCK                       =>      GT1_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT1_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt1_gtrxreset_t,
        MMCM_RESET                      =>      GT1_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT1_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt1_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt1_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt1_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt1_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt1_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt1_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt1_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt2_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT2_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT0_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT0_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt2_rxresetdone_i,
        MMCM_LOCK                       =>      GT2_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT2_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt2_gtrxreset_t,
        MMCM_RESET                      =>      GT2_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT2_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt2_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt2_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt2_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt2_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt2_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt2_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt2_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt3_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT3_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT0_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT0_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt3_rxresetdone_i,
        MMCM_LOCK                       =>      GT3_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT3_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt3_gtrxreset_t,
        MMCM_RESET                      =>      GT3_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT3_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt3_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt3_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt3_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt3_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt3_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt3_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt3_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt4_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT4_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT1_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT1_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt4_rxresetdone_i,
        MMCM_LOCK                       =>      GT4_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT4_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt4_gtrxreset_t,
        MMCM_RESET                      =>      GT4_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT4_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt4_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt4_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt4_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt4_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt4_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt4_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt4_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt5_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT5_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT1_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT1_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt5_rxresetdone_i,
        MMCM_LOCK                       =>      GT5_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT5_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt5_gtrxreset_t,
        MMCM_RESET                      =>      GT5_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT5_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt5_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt5_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt5_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt5_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt5_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt5_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt5_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt6_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT6_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT1_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT1_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt6_rxresetdone_i,
        MMCM_LOCK                       =>      GT6_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT6_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt6_gtrxreset_t,
        MMCM_RESET                      =>      GT6_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT6_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt6_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt6_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt6_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt6_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt6_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt6_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt6_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt7_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT7_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT1_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT1_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt7_rxresetdone_i,
        MMCM_LOCK                       =>      GT7_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT7_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt7_gtrxreset_t,
        MMCM_RESET                      =>      GT7_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT7_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt7_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt7_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt7_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt7_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt7_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt7_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt7_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt8_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT8_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT2_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT2_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt8_rxresetdone_i,
        MMCM_LOCK                       =>      GT8_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT8_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt8_gtrxreset_t,
        MMCM_RESET                      =>      GT8_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT8_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt8_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt8_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt8_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt8_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt8_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt8_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt8_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt9_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT9_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT2_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT2_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt9_rxresetdone_i,
        MMCM_LOCK                       =>      GT9_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT9_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt9_gtrxreset_t,
        MMCM_RESET                      =>      GT9_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT9_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt9_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt9_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt9_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt9_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt9_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt9_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt9_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt10_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT10_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT2_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT2_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt10_rxresetdone_i,
        MMCM_LOCK                       =>      GT10_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT10_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt10_gtrxreset_t,
        MMCM_RESET                      =>      GT10_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT10_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt10_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt10_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt10_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt10_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt10_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt10_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt10_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt11_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT11_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT2_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT2_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt11_rxresetdone_i,
        MMCM_LOCK                       =>      GT11_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT11_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt11_gtrxreset_t,
        MMCM_RESET                      =>      GT11_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT11_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt11_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt11_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt11_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt11_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt11_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt11_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt11_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt12_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT12_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT3_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT3_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt12_rxresetdone_i,
        MMCM_LOCK                       =>      GT12_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT12_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt12_gtrxreset_t,
        MMCM_RESET                      =>      GT12_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT12_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt12_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt12_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt12_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt12_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt12_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt12_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt12_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt13_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT13_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT3_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT3_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt13_rxresetdone_i,
        MMCM_LOCK                       =>      GT13_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT13_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt13_gtrxreset_t,
        MMCM_RESET                      =>      GT13_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT13_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt13_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt13_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt13_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt13_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt13_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt13_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt13_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt14_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT14_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT3_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT3_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt14_rxresetdone_i,
        MMCM_LOCK                       =>      GT14_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT14_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt14_gtrxreset_t,
        MMCM_RESET                      =>      GT14_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT14_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt14_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt14_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt14_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt14_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt14_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt14_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt14_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt15_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT15_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT3_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT3_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt15_rxresetdone_i,
        MMCM_LOCK                       =>      GT15_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT15_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt15_gtrxreset_t,
        MMCM_RESET                      =>      GT15_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT15_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt15_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt15_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt15_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt15_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt15_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt15_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt15_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt16_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT16_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT4_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT4_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt16_rxresetdone_i,
        MMCM_LOCK                       =>      GT16_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT16_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt16_gtrxreset_t,
        MMCM_RESET                      =>      GT16_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT16_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt16_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt16_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt16_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt16_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt16_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt16_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt16_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt17_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT17_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT4_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT4_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt17_rxresetdone_i,
        MMCM_LOCK                       =>      GT17_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT17_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt17_gtrxreset_t,
        MMCM_RESET                      =>      GT17_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT17_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt17_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt17_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt17_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt17_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt17_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt17_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt17_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt18_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT18_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT4_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT4_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt18_rxresetdone_i,
        MMCM_LOCK                       =>      GT18_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT18_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt18_gtrxreset_t,
        MMCM_RESET                      =>      GT18_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT18_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt18_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt18_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt18_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt18_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt18_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt18_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt18_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt19_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT19_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT4_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT4_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt19_rxresetdone_i,
        MMCM_LOCK                       =>      GT19_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT19_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt19_gtrxreset_t,
        MMCM_RESET                      =>      GT19_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT19_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt19_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt19_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt19_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt19_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt19_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt19_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt19_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt20_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT20_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT5_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT5_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt20_rxresetdone_i,
        MMCM_LOCK                       =>      GT20_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT20_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt20_gtrxreset_t,
        MMCM_RESET                      =>      GT20_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT20_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt20_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt20_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt20_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt20_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt20_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt20_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt20_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt21_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT21_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT5_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT5_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt21_rxresetdone_i,
        MMCM_LOCK                       =>      GT21_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT21_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt21_gtrxreset_t,
        MMCM_RESET                      =>      GT21_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT21_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt21_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt21_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt21_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt21_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt21_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt21_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt21_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt22_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT22_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT5_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT5_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt22_rxresetdone_i,
        MMCM_LOCK                       =>      GT22_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT22_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt22_gtrxreset_t,
        MMCM_RESET                      =>      GT22_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT22_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt22_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt22_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt22_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt22_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt22_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt22_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt22_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt23_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT23_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT5_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT5_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt23_rxresetdone_i,
        MMCM_LOCK                       =>      GT23_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT23_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt23_gtrxreset_t,
        MMCM_RESET                      =>      GT23_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT23_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt23_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt23_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt23_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt23_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt23_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt23_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt23_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt24_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT24_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT6_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT6_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt24_rxresetdone_i,
        MMCM_LOCK                       =>      GT24_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT24_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt24_gtrxreset_t,
        MMCM_RESET                      =>      GT24_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT24_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt24_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt24_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt24_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt24_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt24_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt24_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt24_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt25_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT25_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT6_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT6_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt25_rxresetdone_i,
        MMCM_LOCK                       =>      GT25_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT25_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt25_gtrxreset_t,
        MMCM_RESET                      =>      GT25_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT25_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt25_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt25_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt25_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt25_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt25_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt25_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt25_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt26_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT26_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT6_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT6_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt26_rxresetdone_i,
        MMCM_LOCK                       =>      GT26_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT26_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt26_gtrxreset_t,
        MMCM_RESET                      =>      GT26_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT26_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt26_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt26_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt26_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt26_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt26_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt26_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt26_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt27_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT27_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT6_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT6_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt27_rxresetdone_i,
        MMCM_LOCK                       =>      GT27_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT27_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt27_gtrxreset_t,
        MMCM_RESET                      =>      GT27_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT27_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt27_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt27_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt27_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt27_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt27_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt27_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt27_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt28_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT28_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT7_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT7_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt28_rxresetdone_i,
        MMCM_LOCK                       =>      GT28_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT28_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt28_gtrxreset_t,
        MMCM_RESET                      =>      GT28_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT28_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt28_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt28_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt28_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt28_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt28_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt28_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt28_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt29_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT29_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT7_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT7_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt29_rxresetdone_i,
        MMCM_LOCK                       =>      GT29_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT29_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt29_gtrxreset_t,
        MMCM_RESET                      =>      GT29_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT29_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt29_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt29_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt29_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt29_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt29_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt29_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt29_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt30_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT30_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT7_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT7_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt30_rxresetdone_i,
        MMCM_LOCK                       =>      GT30_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT30_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt30_gtrxreset_t,
        MMCM_RESET                      =>      GT30_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT30_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt30_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt30_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt30_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt30_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt30_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt30_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt30_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );


gt31_rxresetfsm_i:  gtwizard_0_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT31_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_RX_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxoutclk_i2,
        QPLLREFCLKLOST                  =>      GT7_QPLLREFCLKLOST_IN,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      GT7_QPLLLOCK_IN,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt31_rxresetdone_i,
        MMCM_LOCK                       =>      GT31_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT31_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt31_gtrxreset_t,
        MMCM_RESET                      =>      GT31_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT31_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt31_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt31_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt31_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt31_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt31_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt31_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt31_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );



  gt0_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt0_gtrxreset_i = '1') then
          gt0_rx_cdrlocked       <= '0';
          gt0_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt0_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt0_rx_cdrlocked       <= '1';
          gt0_rx_cdrlock_counter <= gt0_rx_cdrlock_counter        after DLY;
        else
          gt0_rx_cdrlock_counter <= gt0_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt1_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt1_gtrxreset_i = '1') then
          gt1_rx_cdrlocked       <= '0';
          gt1_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt1_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt1_rx_cdrlocked       <= '1';
          gt1_rx_cdrlock_counter <= gt1_rx_cdrlock_counter        after DLY;
        else
          gt1_rx_cdrlock_counter <= gt1_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt2_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt2_gtrxreset_i = '1') then
          gt2_rx_cdrlocked       <= '0';
          gt2_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt2_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt2_rx_cdrlocked       <= '1';
          gt2_rx_cdrlock_counter <= gt2_rx_cdrlock_counter        after DLY;
        else
          gt2_rx_cdrlock_counter <= gt2_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt3_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt3_gtrxreset_i = '1') then
          gt3_rx_cdrlocked       <= '0';
          gt3_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt3_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt3_rx_cdrlocked       <= '1';
          gt3_rx_cdrlock_counter <= gt3_rx_cdrlock_counter        after DLY;
        else
          gt3_rx_cdrlock_counter <= gt3_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt4_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt4_gtrxreset_i = '1') then
          gt4_rx_cdrlocked       <= '0';
          gt4_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt4_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt4_rx_cdrlocked       <= '1';
          gt4_rx_cdrlock_counter <= gt4_rx_cdrlock_counter        after DLY;
        else
          gt4_rx_cdrlock_counter <= gt4_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt5_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt5_gtrxreset_i = '1') then
          gt5_rx_cdrlocked       <= '0';
          gt5_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt5_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt5_rx_cdrlocked       <= '1';
          gt5_rx_cdrlock_counter <= gt5_rx_cdrlock_counter        after DLY;
        else
          gt5_rx_cdrlock_counter <= gt5_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt6_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt6_gtrxreset_i = '1') then
          gt6_rx_cdrlocked       <= '0';
          gt6_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt6_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt6_rx_cdrlocked       <= '1';
          gt6_rx_cdrlock_counter <= gt6_rx_cdrlock_counter        after DLY;
        else
          gt6_rx_cdrlock_counter <= gt6_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt7_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt7_gtrxreset_i = '1') then
          gt7_rx_cdrlocked       <= '0';
          gt7_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt7_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt7_rx_cdrlocked       <= '1';
          gt7_rx_cdrlock_counter <= gt7_rx_cdrlock_counter        after DLY;
        else
          gt7_rx_cdrlock_counter <= gt7_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt8_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt8_gtrxreset_i = '1') then
          gt8_rx_cdrlocked       <= '0';
          gt8_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt8_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt8_rx_cdrlocked       <= '1';
          gt8_rx_cdrlock_counter <= gt8_rx_cdrlock_counter        after DLY;
        else
          gt8_rx_cdrlock_counter <= gt8_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt9_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt9_gtrxreset_i = '1') then
          gt9_rx_cdrlocked       <= '0';
          gt9_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt9_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt9_rx_cdrlocked       <= '1';
          gt9_rx_cdrlock_counter <= gt9_rx_cdrlock_counter        after DLY;
        else
          gt9_rx_cdrlock_counter <= gt9_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt10_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt10_gtrxreset_i = '1') then
          gt10_rx_cdrlocked       <= '0';
          gt10_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt10_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt10_rx_cdrlocked       <= '1';
          gt10_rx_cdrlock_counter <= gt10_rx_cdrlock_counter        after DLY;
        else
          gt10_rx_cdrlock_counter <= gt10_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt11_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt11_gtrxreset_i = '1') then
          gt11_rx_cdrlocked       <= '0';
          gt11_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt11_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt11_rx_cdrlocked       <= '1';
          gt11_rx_cdrlock_counter <= gt11_rx_cdrlock_counter        after DLY;
        else
          gt11_rx_cdrlock_counter <= gt11_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt12_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt12_gtrxreset_i = '1') then
          gt12_rx_cdrlocked       <= '0';
          gt12_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt12_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt12_rx_cdrlocked       <= '1';
          gt12_rx_cdrlock_counter <= gt12_rx_cdrlock_counter        after DLY;
        else
          gt12_rx_cdrlock_counter <= gt12_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt13_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt13_gtrxreset_i = '1') then
          gt13_rx_cdrlocked       <= '0';
          gt13_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt13_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt13_rx_cdrlocked       <= '1';
          gt13_rx_cdrlock_counter <= gt13_rx_cdrlock_counter        after DLY;
        else
          gt13_rx_cdrlock_counter <= gt13_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt14_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt14_gtrxreset_i = '1') then
          gt14_rx_cdrlocked       <= '0';
          gt14_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt14_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt14_rx_cdrlocked       <= '1';
          gt14_rx_cdrlock_counter <= gt14_rx_cdrlock_counter        after DLY;
        else
          gt14_rx_cdrlock_counter <= gt14_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt15_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt15_gtrxreset_i = '1') then
          gt15_rx_cdrlocked       <= '0';
          gt15_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt15_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt15_rx_cdrlocked       <= '1';
          gt15_rx_cdrlock_counter <= gt15_rx_cdrlock_counter        after DLY;
        else
          gt15_rx_cdrlock_counter <= gt15_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt16_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt16_gtrxreset_i = '1') then
          gt16_rx_cdrlocked       <= '0';
          gt16_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt16_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt16_rx_cdrlocked       <= '1';
          gt16_rx_cdrlock_counter <= gt16_rx_cdrlock_counter        after DLY;
        else
          gt16_rx_cdrlock_counter <= gt16_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt17_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt17_gtrxreset_i = '1') then
          gt17_rx_cdrlocked       <= '0';
          gt17_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt17_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt17_rx_cdrlocked       <= '1';
          gt17_rx_cdrlock_counter <= gt17_rx_cdrlock_counter        after DLY;
        else
          gt17_rx_cdrlock_counter <= gt17_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt18_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt18_gtrxreset_i = '1') then
          gt18_rx_cdrlocked       <= '0';
          gt18_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt18_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt18_rx_cdrlocked       <= '1';
          gt18_rx_cdrlock_counter <= gt18_rx_cdrlock_counter        after DLY;
        else
          gt18_rx_cdrlock_counter <= gt18_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt19_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt19_gtrxreset_i = '1') then
          gt19_rx_cdrlocked       <= '0';
          gt19_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt19_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt19_rx_cdrlocked       <= '1';
          gt19_rx_cdrlock_counter <= gt19_rx_cdrlock_counter        after DLY;
        else
          gt19_rx_cdrlock_counter <= gt19_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt20_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt20_gtrxreset_i = '1') then
          gt20_rx_cdrlocked       <= '0';
          gt20_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt20_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt20_rx_cdrlocked       <= '1';
          gt20_rx_cdrlock_counter <= gt20_rx_cdrlock_counter        after DLY;
        else
          gt20_rx_cdrlock_counter <= gt20_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt21_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt21_gtrxreset_i = '1') then
          gt21_rx_cdrlocked       <= '0';
          gt21_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt21_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt21_rx_cdrlocked       <= '1';
          gt21_rx_cdrlock_counter <= gt21_rx_cdrlock_counter        after DLY;
        else
          gt21_rx_cdrlock_counter <= gt21_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt22_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt22_gtrxreset_i = '1') then
          gt22_rx_cdrlocked       <= '0';
          gt22_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt22_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt22_rx_cdrlocked       <= '1';
          gt22_rx_cdrlock_counter <= gt22_rx_cdrlock_counter        after DLY;
        else
          gt22_rx_cdrlock_counter <= gt22_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt23_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt23_gtrxreset_i = '1') then
          gt23_rx_cdrlocked       <= '0';
          gt23_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt23_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt23_rx_cdrlocked       <= '1';
          gt23_rx_cdrlock_counter <= gt23_rx_cdrlock_counter        after DLY;
        else
          gt23_rx_cdrlock_counter <= gt23_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt24_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt24_gtrxreset_i = '1') then
          gt24_rx_cdrlocked       <= '0';
          gt24_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt24_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt24_rx_cdrlocked       <= '1';
          gt24_rx_cdrlock_counter <= gt24_rx_cdrlock_counter        after DLY;
        else
          gt24_rx_cdrlock_counter <= gt24_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt25_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt25_gtrxreset_i = '1') then
          gt25_rx_cdrlocked       <= '0';
          gt25_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt25_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt25_rx_cdrlocked       <= '1';
          gt25_rx_cdrlock_counter <= gt25_rx_cdrlock_counter        after DLY;
        else
          gt25_rx_cdrlock_counter <= gt25_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt26_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt26_gtrxreset_i = '1') then
          gt26_rx_cdrlocked       <= '0';
          gt26_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt26_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt26_rx_cdrlocked       <= '1';
          gt26_rx_cdrlock_counter <= gt26_rx_cdrlock_counter        after DLY;
        else
          gt26_rx_cdrlock_counter <= gt26_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt27_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt27_gtrxreset_i = '1') then
          gt27_rx_cdrlocked       <= '0';
          gt27_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt27_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt27_rx_cdrlocked       <= '1';
          gt27_rx_cdrlock_counter <= gt27_rx_cdrlock_counter        after DLY;
        else
          gt27_rx_cdrlock_counter <= gt27_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt28_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt28_gtrxreset_i = '1') then
          gt28_rx_cdrlocked       <= '0';
          gt28_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt28_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt28_rx_cdrlocked       <= '1';
          gt28_rx_cdrlock_counter <= gt28_rx_cdrlock_counter        after DLY;
        else
          gt28_rx_cdrlock_counter <= gt28_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt29_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt29_gtrxreset_i = '1') then
          gt29_rx_cdrlocked       <= '0';
          gt29_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt29_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt29_rx_cdrlocked       <= '1';
          gt29_rx_cdrlock_counter <= gt29_rx_cdrlock_counter        after DLY;
        else
          gt29_rx_cdrlock_counter <= gt29_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt30_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt30_gtrxreset_i = '1') then
          gt30_rx_cdrlocked       <= '0';
          gt30_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt30_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt30_rx_cdrlocked       <= '1';
          gt30_rx_cdrlock_counter <= gt30_rx_cdrlock_counter        after DLY;
        else
          gt30_rx_cdrlock_counter <= gt30_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt31_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt31_gtrxreset_i = '1') then
          gt31_rx_cdrlocked       <= '0';
          gt31_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt31_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt31_rx_cdrlocked       <= '1';
          gt31_rx_cdrlock_counter <= gt31_rx_cdrlock_counter        after DLY;
        else
          gt31_rx_cdrlock_counter <= gt31_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

gt0_recclk_stable_i                          <= gt0_rx_cdrlocked;
gt1_recclk_stable_i                          <= gt1_rx_cdrlocked;
gt2_recclk_stable_i                          <= gt2_rx_cdrlocked;
gt3_recclk_stable_i                          <= gt3_rx_cdrlocked;
gt4_recclk_stable_i                          <= gt4_rx_cdrlocked;
gt5_recclk_stable_i                          <= gt5_rx_cdrlocked;
gt6_recclk_stable_i                          <= gt6_rx_cdrlocked;
gt7_recclk_stable_i                          <= gt7_rx_cdrlocked;
gt8_recclk_stable_i                          <= gt8_rx_cdrlocked;
gt9_recclk_stable_i                          <= gt9_rx_cdrlocked;
gt10_recclk_stable_i                         <= gt10_rx_cdrlocked;
gt11_recclk_stable_i                         <= gt11_rx_cdrlocked;
gt12_recclk_stable_i                         <= gt12_rx_cdrlocked;
gt13_recclk_stable_i                         <= gt13_rx_cdrlocked;
gt14_recclk_stable_i                         <= gt14_rx_cdrlocked;
gt15_recclk_stable_i                         <= gt15_rx_cdrlocked;
gt16_recclk_stable_i                         <= gt16_rx_cdrlocked;
gt17_recclk_stable_i                         <= gt17_rx_cdrlocked;
gt18_recclk_stable_i                         <= gt18_rx_cdrlocked;
gt19_recclk_stable_i                         <= gt19_rx_cdrlocked;
gt20_recclk_stable_i                         <= gt20_rx_cdrlocked;
gt21_recclk_stable_i                         <= gt21_rx_cdrlocked;
gt22_recclk_stable_i                         <= gt22_rx_cdrlocked;
gt23_recclk_stable_i                         <= gt23_rx_cdrlocked;
gt24_recclk_stable_i                         <= gt24_rx_cdrlocked;
gt25_recclk_stable_i                         <= gt25_rx_cdrlocked;
gt26_recclk_stable_i                         <= gt26_rx_cdrlocked;
gt27_recclk_stable_i                         <= gt27_rx_cdrlocked;
gt28_recclk_stable_i                         <= gt28_rx_cdrlocked;
gt29_recclk_stable_i                         <= gt29_rx_cdrlocked;
gt30_recclk_stable_i                         <= gt30_rx_cdrlocked;
gt31_recclk_stable_i                         <= gt31_rx_cdrlocked;



    --------------------------- TX Buffer Bypass Logic --------------------
    -- The TX SYNC Module drives the ports needed to Bypass the TX Buffer.
    -- Include the TX SYNC module in your own design if TX Buffer is bypassed.

--Manual
   gt0_tx_manual_phase_i : gtwizard_0_TX_MANUAL_PHASE_ALIGN
   generic map
   ( NUMBER_OF_LANES	  => 12,
     MASTER_LANE_ID       =>  0
   )
   port map
   (
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RESET_PHALIGNMENT               =>      U0_rst_tx_phalignment_i,   --TODO
        RUN_PHALIGNMENT                 =>      U0_run_tx_phalignment_i,      --TODO
        PHASE_ALIGNMENT_DONE            =>      gt0_tx_phalignment_done_i,
        TXDLYSRESET                     =>      U0_TXDLYSRESET,
        TXDLYSRESETDONE                 =>      U0_TXDLYSRESETDONE,
        TXPHINIT                        =>      U0_TXPHINIT,
        TXPHINITDONE                    =>      U0_TXPHINITDONE,
        TXPHALIGN                       =>      U0_TXPHALIGN,
        TXPHALIGNDONE                   =>      U0_TXPHALIGNDONE,
        TXDLYEN                         =>      U0_TXDLYEN
   );

gt0_txphdlyreset_i                           <= tied_to_ground_i;
gt0_txphalignen_i                            <= tied_to_vcc_i;
gt0_txdlysreset_i                            <= U0_TXDLYSRESET(0);
gt0_txphinit_i                               <= U0_TXPHINIT(0);
gt0_txphalign_i                              <= U0_TXPHALIGN(0);
gt0_txdlyen_i                                <= U0_TXDLYEN(0);
U0_TXDLYSRESETDONE(0)                        <= gt0_txdlysresetdone_i;
U0_TXPHINITDONE(0)                           <= gt0_txphinitdone_i;
U0_TXPHALIGNDONE(0)                          <= gt0_txphaligndone_i;

gt0_txsyncallin_i                            <= gt0_txphaligndone_i;
gt0_txsyncin_i                               <= gt0_txsyncout_i;
gt0_txsyncmode_i                             <= tied_to_vcc_i;

 
gt1_txdlysreset_i                            <= U0_TXDLYSRESET(1);
gt1_txphinit_i                               <= U0_TXPHINIT(1);
gt1_txphalign_i                              <= U0_TXPHALIGN(1);
gt1_txphalignen_i                            <= tied_to_vcc_i;
gt1_txphdlyreset_i                           <= tied_to_ground_i;
gt1_txdlyen_i                                <= tied_to_ground_i;
U0_TXDLYSRESETDONE(1)                        <= gt1_txdlysresetdone_i;
U0_TXPHINITDONE(1)                           <= gt1_txphinitdone_i;
U0_TXPHALIGNDONE(1)                          <= gt1_txphaligndone_i;

gt1_txsyncallin_i                            <= tied_to_ground_i;
gt1_txsyncin_i                               <= tied_to_ground_i;
gt1_txsyncmode_i                             <= tied_to_ground_i;
 
gt2_txdlysreset_i                            <= U0_TXDLYSRESET(2);
gt2_txphinit_i                               <= U0_TXPHINIT(2);
gt2_txphalign_i                              <= U0_TXPHALIGN(2);
gt2_txphalignen_i                            <= tied_to_vcc_i;
gt2_txphdlyreset_i                           <= tied_to_ground_i;
gt2_txdlyen_i                                <= tied_to_ground_i;
U0_TXDLYSRESETDONE(2)                        <= gt2_txdlysresetdone_i;
U0_TXPHINITDONE(2)                           <= gt2_txphinitdone_i;
U0_TXPHALIGNDONE(2)                          <= gt2_txphaligndone_i;

gt2_txsyncallin_i                            <= tied_to_ground_i;
gt2_txsyncin_i                               <= tied_to_ground_i;
gt2_txsyncmode_i                             <= tied_to_ground_i;
 
gt3_txdlysreset_i                            <= U0_TXDLYSRESET(3);
gt3_txphinit_i                               <= U0_TXPHINIT(3);
gt3_txphalign_i                              <= U0_TXPHALIGN(3);
gt3_txphalignen_i                            <= tied_to_vcc_i;
gt3_txphdlyreset_i                           <= tied_to_ground_i;
gt3_txdlyen_i                                <= tied_to_ground_i;
U0_TXDLYSRESETDONE(3)                        <= gt3_txdlysresetdone_i;
U0_TXPHINITDONE(3)                           <= gt3_txphinitdone_i;
U0_TXPHALIGNDONE(3)                          <= gt3_txphaligndone_i;

gt3_txsyncallin_i                            <= tied_to_ground_i;
gt3_txsyncin_i                               <= tied_to_ground_i;
gt3_txsyncmode_i                             <= tied_to_ground_i;
 
gt4_txdlysreset_i                            <= U0_TXDLYSRESET(4);
gt4_txphinit_i                               <= U0_TXPHINIT(4);
gt4_txphalign_i                              <= U0_TXPHALIGN(4);
gt4_txphalignen_i                            <= tied_to_vcc_i;
gt4_txphdlyreset_i                           <= tied_to_ground_i;
gt4_txdlyen_i                                <= tied_to_ground_i;
U0_TXDLYSRESETDONE(4)                        <= gt4_txdlysresetdone_i;
U0_TXPHINITDONE(4)                           <= gt4_txphinitdone_i;
U0_TXPHALIGNDONE(4)                          <= gt4_txphaligndone_i;

gt4_txsyncallin_i                            <= tied_to_ground_i;
gt4_txsyncin_i                               <= tied_to_ground_i;
gt4_txsyncmode_i                             <= tied_to_ground_i;
 
gt5_txdlysreset_i                            <= U0_TXDLYSRESET(5);
gt5_txphinit_i                               <= U0_TXPHINIT(5);
gt5_txphalign_i                              <= U0_TXPHALIGN(5);
gt5_txphalignen_i                            <= tied_to_vcc_i;
gt5_txphdlyreset_i                           <= tied_to_ground_i;
gt5_txdlyen_i                                <= tied_to_ground_i;
U0_TXDLYSRESETDONE(5)                        <= gt5_txdlysresetdone_i;
U0_TXPHINITDONE(5)                           <= gt5_txphinitdone_i;
U0_TXPHALIGNDONE(5)                          <= gt5_txphaligndone_i;

gt5_txsyncallin_i                            <= tied_to_ground_i;
gt5_txsyncin_i                               <= tied_to_ground_i;
gt5_txsyncmode_i                             <= tied_to_ground_i;
 
gt6_txdlysreset_i                            <= U0_TXDLYSRESET(6);
gt6_txphinit_i                               <= U0_TXPHINIT(6);
gt6_txphalign_i                              <= U0_TXPHALIGN(6);
gt6_txphalignen_i                            <= tied_to_vcc_i;
gt6_txphdlyreset_i                           <= tied_to_ground_i;
gt6_txdlyen_i                                <= tied_to_ground_i;
U0_TXDLYSRESETDONE(6)                        <= gt6_txdlysresetdone_i;
U0_TXPHINITDONE(6)                           <= gt6_txphinitdone_i;
U0_TXPHALIGNDONE(6)                          <= gt6_txphaligndone_i;

gt6_txsyncallin_i                            <= tied_to_ground_i;
gt6_txsyncin_i                               <= tied_to_ground_i;
gt6_txsyncmode_i                             <= tied_to_ground_i;
 
gt7_txdlysreset_i                            <= U0_TXDLYSRESET(7);
gt7_txphinit_i                               <= U0_TXPHINIT(7);
gt7_txphalign_i                              <= U0_TXPHALIGN(7);
gt7_txphalignen_i                            <= tied_to_vcc_i;
gt7_txphdlyreset_i                           <= tied_to_ground_i;
gt7_txdlyen_i                                <= tied_to_ground_i;
U0_TXDLYSRESETDONE(7)                        <= gt7_txdlysresetdone_i;
U0_TXPHINITDONE(7)                           <= gt7_txphinitdone_i;
U0_TXPHALIGNDONE(7)                          <= gt7_txphaligndone_i;

gt7_txsyncallin_i                            <= tied_to_ground_i;
gt7_txsyncin_i                               <= tied_to_ground_i;
gt7_txsyncmode_i                             <= tied_to_ground_i;
 
gt8_txdlysreset_i                            <= U0_TXDLYSRESET(8);
gt8_txphinit_i                               <= U0_TXPHINIT(8);
gt8_txphalign_i                              <= U0_TXPHALIGN(8);
gt8_txphalignen_i                            <= tied_to_vcc_i;
gt8_txphdlyreset_i                           <= tied_to_ground_i;
gt8_txdlyen_i                                <= tied_to_ground_i;
U0_TXDLYSRESETDONE(8)                        <= gt8_txdlysresetdone_i;
U0_TXPHINITDONE(8)                           <= gt8_txphinitdone_i;
U0_TXPHALIGNDONE(8)                          <= gt8_txphaligndone_i;

gt8_txsyncallin_i                            <= tied_to_ground_i;
gt8_txsyncin_i                               <= tied_to_ground_i;
gt8_txsyncmode_i                             <= tied_to_ground_i;
 
gt9_txdlysreset_i                            <= U0_TXDLYSRESET(9);
gt9_txphinit_i                               <= U0_TXPHINIT(9);
gt9_txphalign_i                              <= U0_TXPHALIGN(9);
gt9_txphalignen_i                            <= tied_to_vcc_i;
gt9_txphdlyreset_i                           <= tied_to_ground_i;
gt9_txdlyen_i                                <= tied_to_ground_i;
U0_TXDLYSRESETDONE(9)                        <= gt9_txdlysresetdone_i;
U0_TXPHINITDONE(9)                           <= gt9_txphinitdone_i;
U0_TXPHALIGNDONE(9)                          <= gt9_txphaligndone_i;

gt9_txsyncallin_i                            <= tied_to_ground_i;
gt9_txsyncin_i                               <= tied_to_ground_i;
gt9_txsyncmode_i                             <= tied_to_ground_i;
 
gt10_txdlysreset_i                           <= U0_TXDLYSRESET(10);
gt10_txphinit_i                              <= U0_TXPHINIT(10);
gt10_txphalign_i                             <= U0_TXPHALIGN(10);
gt10_txphalignen_i                           <= tied_to_vcc_i;
gt10_txphdlyreset_i                          <= tied_to_ground_i;
gt10_txdlyen_i                               <= tied_to_ground_i;
U0_TXDLYSRESETDONE(10)                       <= gt10_txdlysresetdone_i;
U0_TXPHINITDONE(10)                          <= gt10_txphinitdone_i;
U0_TXPHALIGNDONE(10)                         <= gt10_txphaligndone_i;

gt10_txsyncallin_i                           <= tied_to_ground_i;
gt10_txsyncin_i                              <= tied_to_ground_i;
gt10_txsyncmode_i                            <= tied_to_ground_i;
 
gt11_txdlysreset_i                           <= U0_TXDLYSRESET(11);
gt11_txphinit_i                              <= U0_TXPHINIT(11);
gt11_txphalign_i                             <= U0_TXPHALIGN(11);
gt11_txphalignen_i                           <= tied_to_vcc_i;
gt11_txphdlyreset_i                          <= tied_to_ground_i;
gt11_txdlyen_i                               <= tied_to_ground_i;
U0_TXDLYSRESETDONE(11)                       <= gt11_txdlysresetdone_i;
U0_TXPHINITDONE(11)                          <= gt11_txphinitdone_i;
U0_TXPHALIGNDONE(11)                         <= gt11_txphaligndone_i;

gt11_txsyncallin_i                           <= tied_to_ground_i;
gt11_txsyncin_i                              <= tied_to_ground_i;
gt11_txsyncmode_i                            <= tied_to_ground_i;

    U0_run_tx_phalignment_i    <=  gt0_run_tx_phalignment_i 
 
                                             and gt1_run_tx_phalignment_i
 
                                             and gt2_run_tx_phalignment_i
 
                                             and gt3_run_tx_phalignment_i
 
                                             and gt4_run_tx_phalignment_i
 
                                             and gt5_run_tx_phalignment_i
 
                                             and gt6_run_tx_phalignment_i
 
                                             and gt7_run_tx_phalignment_i
 
                                             and gt8_run_tx_phalignment_i
 
                                             and gt9_run_tx_phalignment_i
 
                                             and gt10_run_tx_phalignment_i
 
                                             and gt11_run_tx_phalignment_i
                                             ;

    U0_rst_tx_phalignment_i    <=  gt0_rst_tx_phalignment_i 
 
                                             or gt1_rst_tx_phalignment_i
 
                                             or gt2_rst_tx_phalignment_i
 
                                             or gt3_rst_tx_phalignment_i
 
                                             or gt4_rst_tx_phalignment_i
 
                                             or gt5_rst_tx_phalignment_i
 
                                             or gt6_rst_tx_phalignment_i
 
                                             or gt7_rst_tx_phalignment_i
 
                                             or gt8_rst_tx_phalignment_i
 
                                             or gt9_rst_tx_phalignment_i
 
                                             or gt10_rst_tx_phalignment_i
 
                                             or gt11_rst_tx_phalignment_i
                                             ;

--Manual
   gt12_tx_manual_phase_i : gtwizard_0_TX_MANUAL_PHASE_ALIGN
   generic map
   ( NUMBER_OF_LANES	  => 12,
     MASTER_LANE_ID       =>  0
   )
   port map
   (
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RESET_PHALIGNMENT               =>      U12_rst_tx_phalignment_i,   --TODO
        RUN_PHALIGNMENT                 =>      U12_run_tx_phalignment_i,      --TODO
        PHASE_ALIGNMENT_DONE            =>      gt12_tx_phalignment_done_i,
        TXDLYSRESET                     =>      U12_TXDLYSRESET,
        TXDLYSRESETDONE                 =>      U12_TXDLYSRESETDONE,
        TXPHINIT                        =>      U12_TXPHINIT,
        TXPHINITDONE                    =>      U12_TXPHINITDONE,
        TXPHALIGN                       =>      U12_TXPHALIGN,
        TXPHALIGNDONE                   =>      U12_TXPHALIGNDONE,
        TXDLYEN                         =>      U12_TXDLYEN
   );

gt12_txphdlyreset_i                          <= tied_to_ground_i;
gt12_txphalignen_i                           <= tied_to_vcc_i;
gt12_txdlysreset_i                           <= U12_TXDLYSRESET(0);
gt12_txphinit_i                              <= U12_TXPHINIT(0);
gt12_txphalign_i                             <= U12_TXPHALIGN(0);
gt12_txdlyen_i                               <= U12_TXDLYEN(0);
U12_TXDLYSRESETDONE(0)                       <= gt12_txdlysresetdone_i;
U12_TXPHINITDONE(0)                          <= gt12_txphinitdone_i;
U12_TXPHALIGNDONE(0)                         <= gt12_txphaligndone_i;

gt12_txsyncallin_i                           <= gt12_txphaligndone_i;
gt12_txsyncin_i                              <= gt12_txsyncout_i;
gt12_txsyncmode_i                            <= tied_to_vcc_i;

 
gt13_txdlysreset_i                           <= U12_TXDLYSRESET(1);
gt13_txphinit_i                              <= U12_TXPHINIT(1);
gt13_txphalign_i                             <= U12_TXPHALIGN(1);
gt13_txphalignen_i                           <= tied_to_vcc_i;
gt13_txphdlyreset_i                          <= tied_to_ground_i;
gt13_txdlyen_i                               <= tied_to_ground_i;
U12_TXDLYSRESETDONE(1)                       <= gt13_txdlysresetdone_i;
U12_TXPHINITDONE(1)                          <= gt13_txphinitdone_i;
U12_TXPHALIGNDONE(1)                         <= gt13_txphaligndone_i;

gt13_txsyncallin_i                           <= tied_to_ground_i;
gt13_txsyncin_i                              <= tied_to_ground_i;
gt13_txsyncmode_i                            <= tied_to_ground_i;
 
gt14_txdlysreset_i                           <= U12_TXDLYSRESET(2);
gt14_txphinit_i                              <= U12_TXPHINIT(2);
gt14_txphalign_i                             <= U12_TXPHALIGN(2);
gt14_txphalignen_i                           <= tied_to_vcc_i;
gt14_txphdlyreset_i                          <= tied_to_ground_i;
gt14_txdlyen_i                               <= tied_to_ground_i;
U12_TXDLYSRESETDONE(2)                       <= gt14_txdlysresetdone_i;
U12_TXPHINITDONE(2)                          <= gt14_txphinitdone_i;
U12_TXPHALIGNDONE(2)                         <= gt14_txphaligndone_i;

gt14_txsyncallin_i                           <= tied_to_ground_i;
gt14_txsyncin_i                              <= tied_to_ground_i;
gt14_txsyncmode_i                            <= tied_to_ground_i;
 
gt15_txdlysreset_i                           <= U12_TXDLYSRESET(3);
gt15_txphinit_i                              <= U12_TXPHINIT(3);
gt15_txphalign_i                             <= U12_TXPHALIGN(3);
gt15_txphalignen_i                           <= tied_to_vcc_i;
gt15_txphdlyreset_i                          <= tied_to_ground_i;
gt15_txdlyen_i                               <= tied_to_ground_i;
U12_TXDLYSRESETDONE(3)                       <= gt15_txdlysresetdone_i;
U12_TXPHINITDONE(3)                          <= gt15_txphinitdone_i;
U12_TXPHALIGNDONE(3)                         <= gt15_txphaligndone_i;

gt15_txsyncallin_i                           <= tied_to_ground_i;
gt15_txsyncin_i                              <= tied_to_ground_i;
gt15_txsyncmode_i                            <= tied_to_ground_i;
 
gt16_txdlysreset_i                           <= U12_TXDLYSRESET(4);
gt16_txphinit_i                              <= U12_TXPHINIT(4);
gt16_txphalign_i                             <= U12_TXPHALIGN(4);
gt16_txphalignen_i                           <= tied_to_vcc_i;
gt16_txphdlyreset_i                          <= tied_to_ground_i;
gt16_txdlyen_i                               <= tied_to_ground_i;
U12_TXDLYSRESETDONE(4)                       <= gt16_txdlysresetdone_i;
U12_TXPHINITDONE(4)                          <= gt16_txphinitdone_i;
U12_TXPHALIGNDONE(4)                         <= gt16_txphaligndone_i;

gt16_txsyncallin_i                           <= tied_to_ground_i;
gt16_txsyncin_i                              <= tied_to_ground_i;
gt16_txsyncmode_i                            <= tied_to_ground_i;
 
gt17_txdlysreset_i                           <= U12_TXDLYSRESET(5);
gt17_txphinit_i                              <= U12_TXPHINIT(5);
gt17_txphalign_i                             <= U12_TXPHALIGN(5);
gt17_txphalignen_i                           <= tied_to_vcc_i;
gt17_txphdlyreset_i                          <= tied_to_ground_i;
gt17_txdlyen_i                               <= tied_to_ground_i;
U12_TXDLYSRESETDONE(5)                       <= gt17_txdlysresetdone_i;
U12_TXPHINITDONE(5)                          <= gt17_txphinitdone_i;
U12_TXPHALIGNDONE(5)                         <= gt17_txphaligndone_i;

gt17_txsyncallin_i                           <= tied_to_ground_i;
gt17_txsyncin_i                              <= tied_to_ground_i;
gt17_txsyncmode_i                            <= tied_to_ground_i;
 
gt18_txdlysreset_i                           <= U12_TXDLYSRESET(6);
gt18_txphinit_i                              <= U12_TXPHINIT(6);
gt18_txphalign_i                             <= U12_TXPHALIGN(6);
gt18_txphalignen_i                           <= tied_to_vcc_i;
gt18_txphdlyreset_i                          <= tied_to_ground_i;
gt18_txdlyen_i                               <= tied_to_ground_i;
U12_TXDLYSRESETDONE(6)                       <= gt18_txdlysresetdone_i;
U12_TXPHINITDONE(6)                          <= gt18_txphinitdone_i;
U12_TXPHALIGNDONE(6)                         <= gt18_txphaligndone_i;

gt18_txsyncallin_i                           <= tied_to_ground_i;
gt18_txsyncin_i                              <= tied_to_ground_i;
gt18_txsyncmode_i                            <= tied_to_ground_i;
 
gt19_txdlysreset_i                           <= U12_TXDLYSRESET(7);
gt19_txphinit_i                              <= U12_TXPHINIT(7);
gt19_txphalign_i                             <= U12_TXPHALIGN(7);
gt19_txphalignen_i                           <= tied_to_vcc_i;
gt19_txphdlyreset_i                          <= tied_to_ground_i;
gt19_txdlyen_i                               <= tied_to_ground_i;
U12_TXDLYSRESETDONE(7)                       <= gt19_txdlysresetdone_i;
U12_TXPHINITDONE(7)                          <= gt19_txphinitdone_i;
U12_TXPHALIGNDONE(7)                         <= gt19_txphaligndone_i;

gt19_txsyncallin_i                           <= tied_to_ground_i;
gt19_txsyncin_i                              <= tied_to_ground_i;
gt19_txsyncmode_i                            <= tied_to_ground_i;
 
gt20_txdlysreset_i                           <= U12_TXDLYSRESET(8);
gt20_txphinit_i                              <= U12_TXPHINIT(8);
gt20_txphalign_i                             <= U12_TXPHALIGN(8);
gt20_txphalignen_i                           <= tied_to_vcc_i;
gt20_txphdlyreset_i                          <= tied_to_ground_i;
gt20_txdlyen_i                               <= tied_to_ground_i;
U12_TXDLYSRESETDONE(8)                       <= gt20_txdlysresetdone_i;
U12_TXPHINITDONE(8)                          <= gt20_txphinitdone_i;
U12_TXPHALIGNDONE(8)                         <= gt20_txphaligndone_i;

gt20_txsyncallin_i                           <= tied_to_ground_i;
gt20_txsyncin_i                              <= tied_to_ground_i;
gt20_txsyncmode_i                            <= tied_to_ground_i;
 
gt21_txdlysreset_i                           <= U12_TXDLYSRESET(9);
gt21_txphinit_i                              <= U12_TXPHINIT(9);
gt21_txphalign_i                             <= U12_TXPHALIGN(9);
gt21_txphalignen_i                           <= tied_to_vcc_i;
gt21_txphdlyreset_i                          <= tied_to_ground_i;
gt21_txdlyen_i                               <= tied_to_ground_i;
U12_TXDLYSRESETDONE(9)                       <= gt21_txdlysresetdone_i;
U12_TXPHINITDONE(9)                          <= gt21_txphinitdone_i;
U12_TXPHALIGNDONE(9)                         <= gt21_txphaligndone_i;

gt21_txsyncallin_i                           <= tied_to_ground_i;
gt21_txsyncin_i                              <= tied_to_ground_i;
gt21_txsyncmode_i                            <= tied_to_ground_i;
 
gt22_txdlysreset_i                           <= U12_TXDLYSRESET(10);
gt22_txphinit_i                              <= U12_TXPHINIT(10);
gt22_txphalign_i                             <= U12_TXPHALIGN(10);
gt22_txphalignen_i                           <= tied_to_vcc_i;
gt22_txphdlyreset_i                          <= tied_to_ground_i;
gt22_txdlyen_i                               <= tied_to_ground_i;
U12_TXDLYSRESETDONE(10)                      <= gt22_txdlysresetdone_i;
U12_TXPHINITDONE(10)                         <= gt22_txphinitdone_i;
U12_TXPHALIGNDONE(10)                        <= gt22_txphaligndone_i;

gt22_txsyncallin_i                           <= tied_to_ground_i;
gt22_txsyncin_i                              <= tied_to_ground_i;
gt22_txsyncmode_i                            <= tied_to_ground_i;
 
gt23_txdlysreset_i                           <= U12_TXDLYSRESET(11);
gt23_txphinit_i                              <= U12_TXPHINIT(11);
gt23_txphalign_i                             <= U12_TXPHALIGN(11);
gt23_txphalignen_i                           <= tied_to_vcc_i;
gt23_txphdlyreset_i                          <= tied_to_ground_i;
gt23_txdlyen_i                               <= tied_to_ground_i;
U12_TXDLYSRESETDONE(11)                      <= gt23_txdlysresetdone_i;
U12_TXPHINITDONE(11)                         <= gt23_txphinitdone_i;
U12_TXPHALIGNDONE(11)                        <= gt23_txphaligndone_i;

gt23_txsyncallin_i                           <= tied_to_ground_i;
gt23_txsyncin_i                              <= tied_to_ground_i;
gt23_txsyncmode_i                            <= tied_to_ground_i;

    U12_run_tx_phalignment_i    <=  gt12_run_tx_phalignment_i 
 
                                             and gt13_run_tx_phalignment_i
 
                                             and gt14_run_tx_phalignment_i
 
                                             and gt15_run_tx_phalignment_i
 
                                             and gt16_run_tx_phalignment_i
 
                                             and gt17_run_tx_phalignment_i
 
                                             and gt18_run_tx_phalignment_i
 
                                             and gt19_run_tx_phalignment_i
 
                                             and gt20_run_tx_phalignment_i
 
                                             and gt21_run_tx_phalignment_i
 
                                             and gt22_run_tx_phalignment_i
 
                                             and gt23_run_tx_phalignment_i
                                             ;

    U12_rst_tx_phalignment_i    <=  gt12_rst_tx_phalignment_i 
 
                                             or gt13_rst_tx_phalignment_i
 
                                             or gt14_rst_tx_phalignment_i
 
                                             or gt15_rst_tx_phalignment_i
 
                                             or gt16_rst_tx_phalignment_i
 
                                             or gt17_rst_tx_phalignment_i
 
                                             or gt18_rst_tx_phalignment_i
 
                                             or gt19_rst_tx_phalignment_i
 
                                             or gt20_rst_tx_phalignment_i
 
                                             or gt21_rst_tx_phalignment_i
 
                                             or gt22_rst_tx_phalignment_i
 
                                             or gt23_rst_tx_phalignment_i
                                             ;

--Manual
   gt24_tx_manual_phase_i : gtwizard_0_TX_MANUAL_PHASE_ALIGN
   generic map
   ( NUMBER_OF_LANES	  => 8,
     MASTER_LANE_ID       =>  0
   )
   port map
   (
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RESET_PHALIGNMENT               =>      U24_rst_tx_phalignment_i,   --TODO
        RUN_PHALIGNMENT                 =>      U24_run_tx_phalignment_i,      --TODO
        PHASE_ALIGNMENT_DONE            =>      gt24_tx_phalignment_done_i,
        TXDLYSRESET                     =>      U24_TXDLYSRESET,
        TXDLYSRESETDONE                 =>      U24_TXDLYSRESETDONE,
        TXPHINIT                        =>      U24_TXPHINIT,
        TXPHINITDONE                    =>      U24_TXPHINITDONE,
        TXPHALIGN                       =>      U24_TXPHALIGN,
        TXPHALIGNDONE                   =>      U24_TXPHALIGNDONE,
        TXDLYEN                         =>      U24_TXDLYEN
   );

gt24_txphdlyreset_i                          <= tied_to_ground_i;
gt24_txphalignen_i                           <= tied_to_vcc_i;
gt24_txdlysreset_i                           <= U24_TXDLYSRESET(0);
gt24_txphinit_i                              <= U24_TXPHINIT(0);
gt24_txphalign_i                             <= U24_TXPHALIGN(0);
gt24_txdlyen_i                               <= U24_TXDLYEN(0);
U24_TXDLYSRESETDONE(0)                       <= gt24_txdlysresetdone_i;
U24_TXPHINITDONE(0)                          <= gt24_txphinitdone_i;
U24_TXPHALIGNDONE(0)                         <= gt24_txphaligndone_i;

gt24_txsyncallin_i                           <= gt24_txphaligndone_i;
gt24_txsyncin_i                              <= gt24_txsyncout_i;
gt24_txsyncmode_i                            <= tied_to_vcc_i;

 
gt25_txdlysreset_i                           <= U24_TXDLYSRESET(1);
gt25_txphinit_i                              <= U24_TXPHINIT(1);
gt25_txphalign_i                             <= U24_TXPHALIGN(1);
gt25_txphalignen_i                           <= tied_to_vcc_i;
gt25_txphdlyreset_i                          <= tied_to_ground_i;
gt25_txdlyen_i                               <= tied_to_ground_i;
U24_TXDLYSRESETDONE(1)                       <= gt25_txdlysresetdone_i;
U24_TXPHINITDONE(1)                          <= gt25_txphinitdone_i;
U24_TXPHALIGNDONE(1)                         <= gt25_txphaligndone_i;

gt25_txsyncallin_i                           <= tied_to_ground_i;
gt25_txsyncin_i                              <= tied_to_ground_i;
gt25_txsyncmode_i                            <= tied_to_ground_i;
 
gt26_txdlysreset_i                           <= U24_TXDLYSRESET(2);
gt26_txphinit_i                              <= U24_TXPHINIT(2);
gt26_txphalign_i                             <= U24_TXPHALIGN(2);
gt26_txphalignen_i                           <= tied_to_vcc_i;
gt26_txphdlyreset_i                          <= tied_to_ground_i;
gt26_txdlyen_i                               <= tied_to_ground_i;
U24_TXDLYSRESETDONE(2)                       <= gt26_txdlysresetdone_i;
U24_TXPHINITDONE(2)                          <= gt26_txphinitdone_i;
U24_TXPHALIGNDONE(2)                         <= gt26_txphaligndone_i;

gt26_txsyncallin_i                           <= tied_to_ground_i;
gt26_txsyncin_i                              <= tied_to_ground_i;
gt26_txsyncmode_i                            <= tied_to_ground_i;
 
gt27_txdlysreset_i                           <= U24_TXDLYSRESET(3);
gt27_txphinit_i                              <= U24_TXPHINIT(3);
gt27_txphalign_i                             <= U24_TXPHALIGN(3);
gt27_txphalignen_i                           <= tied_to_vcc_i;
gt27_txphdlyreset_i                          <= tied_to_ground_i;
gt27_txdlyen_i                               <= tied_to_ground_i;
U24_TXDLYSRESETDONE(3)                       <= gt27_txdlysresetdone_i;
U24_TXPHINITDONE(3)                          <= gt27_txphinitdone_i;
U24_TXPHALIGNDONE(3)                         <= gt27_txphaligndone_i;

gt27_txsyncallin_i                           <= tied_to_ground_i;
gt27_txsyncin_i                              <= tied_to_ground_i;
gt27_txsyncmode_i                            <= tied_to_ground_i;
 
gt28_txdlysreset_i                           <= U24_TXDLYSRESET(4);
gt28_txphinit_i                              <= U24_TXPHINIT(4);
gt28_txphalign_i                             <= U24_TXPHALIGN(4);
gt28_txphalignen_i                           <= tied_to_vcc_i;
gt28_txphdlyreset_i                          <= tied_to_ground_i;
gt28_txdlyen_i                               <= tied_to_ground_i;
U24_TXDLYSRESETDONE(4)                       <= gt28_txdlysresetdone_i;
U24_TXPHINITDONE(4)                          <= gt28_txphinitdone_i;
U24_TXPHALIGNDONE(4)                         <= gt28_txphaligndone_i;

gt28_txsyncallin_i                           <= tied_to_ground_i;
gt28_txsyncin_i                              <= tied_to_ground_i;
gt28_txsyncmode_i                            <= tied_to_ground_i;
 
gt29_txdlysreset_i                           <= U24_TXDLYSRESET(5);
gt29_txphinit_i                              <= U24_TXPHINIT(5);
gt29_txphalign_i                             <= U24_TXPHALIGN(5);
gt29_txphalignen_i                           <= tied_to_vcc_i;
gt29_txphdlyreset_i                          <= tied_to_ground_i;
gt29_txdlyen_i                               <= tied_to_ground_i;
U24_TXDLYSRESETDONE(5)                       <= gt29_txdlysresetdone_i;
U24_TXPHINITDONE(5)                          <= gt29_txphinitdone_i;
U24_TXPHALIGNDONE(5)                         <= gt29_txphaligndone_i;

gt29_txsyncallin_i                           <= tied_to_ground_i;
gt29_txsyncin_i                              <= tied_to_ground_i;
gt29_txsyncmode_i                            <= tied_to_ground_i;
 
gt30_txdlysreset_i                           <= U24_TXDLYSRESET(6);
gt30_txphinit_i                              <= U24_TXPHINIT(6);
gt30_txphalign_i                             <= U24_TXPHALIGN(6);
gt30_txphalignen_i                           <= tied_to_vcc_i;
gt30_txphdlyreset_i                          <= tied_to_ground_i;
gt30_txdlyen_i                               <= tied_to_ground_i;
U24_TXDLYSRESETDONE(6)                       <= gt30_txdlysresetdone_i;
U24_TXPHINITDONE(6)                          <= gt30_txphinitdone_i;
U24_TXPHALIGNDONE(6)                         <= gt30_txphaligndone_i;

gt30_txsyncallin_i                           <= tied_to_ground_i;
gt30_txsyncin_i                              <= tied_to_ground_i;
gt30_txsyncmode_i                            <= tied_to_ground_i;
 
gt31_txdlysreset_i                           <= U24_TXDLYSRESET(7);
gt31_txphinit_i                              <= U24_TXPHINIT(7);
gt31_txphalign_i                             <= U24_TXPHALIGN(7);
gt31_txphalignen_i                           <= tied_to_vcc_i;
gt31_txphdlyreset_i                          <= tied_to_ground_i;
gt31_txdlyen_i                               <= tied_to_ground_i;
U24_TXDLYSRESETDONE(7)                       <= gt31_txdlysresetdone_i;
U24_TXPHINITDONE(7)                          <= gt31_txphinitdone_i;
U24_TXPHALIGNDONE(7)                         <= gt31_txphaligndone_i;

gt31_txsyncallin_i                           <= tied_to_ground_i;
gt31_txsyncin_i                              <= tied_to_ground_i;
gt31_txsyncmode_i                            <= tied_to_ground_i;

    U24_run_tx_phalignment_i    <=  gt24_run_tx_phalignment_i 
 
                                             and gt25_run_tx_phalignment_i
 
                                             and gt26_run_tx_phalignment_i
 
                                             and gt27_run_tx_phalignment_i
 
                                             and gt28_run_tx_phalignment_i
 
                                             and gt29_run_tx_phalignment_i
 
                                             and gt30_run_tx_phalignment_i
 
                                             and gt31_run_tx_phalignment_i
                                             ;

    U24_rst_tx_phalignment_i    <=  gt24_rst_tx_phalignment_i 
 
                                             or gt25_rst_tx_phalignment_i
 
                                             or gt26_rst_tx_phalignment_i
 
                                             or gt27_rst_tx_phalignment_i
 
                                             or gt28_rst_tx_phalignment_i
 
                                             or gt29_rst_tx_phalignment_i
 
                                             or gt30_rst_tx_phalignment_i
 
                                             or gt31_rst_tx_phalignment_i
                                             ;



   --------------------------- RX Buffer Bypass Logic --------------------
--   The RX SYNC Module drives the ports needed to Bypass the RX Buffer.
--   Include the RX SYNC module in your own design if RX Buffer is bypassed.


--Auto
--Master

gt0_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt0_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt0_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt0_rxsyncdone_i,
        DLYSRESET                       =>      gt0_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt0_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );

gt0_rxphdlyreset_i                           <= tied_to_ground_i;
gt0_rxphalignen_i                            <= tied_to_ground_i;
gt0_rxdlyen_i                                <= tied_to_ground_i;
gt0_rxphalign_i                              <= tied_to_ground_i;
gt0_rxsyncallin_i                            <= rxmstr0_rxsyncallin_i;
gt0_rxsyncmode_i                             <= tied_to_vcc_i;
gt0_rxsyncin_i                               <= gt0_rxsyncout_i;


gt1_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt1_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt1_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt1_rxphaligndone_i,
        DLYSRESET                       =>      gt1_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt1_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );
gt1_rxphdlyreset_i                           <= tied_to_ground_i;
gt1_rxphalignen_i                            <= tied_to_ground_i;
gt1_rxdlyen_i                                <= tied_to_ground_i;
gt1_rxphalign_i                              <= tied_to_ground_i;
gt1_rxsyncallin_i                            <= rxmstr0_rxsyncallin_i;
gt1_rxsyncmode_i                             <= tied_to_ground_i;
gt1_rxsyncin_i                               <= gt0_rxsyncout_i;
gt2_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt2_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt2_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt2_rxphaligndone_i,
        DLYSRESET                       =>      gt2_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt2_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );
gt2_rxphdlyreset_i                           <= tied_to_ground_i;
gt2_rxphalignen_i                            <= tied_to_ground_i;
gt2_rxdlyen_i                                <= tied_to_ground_i;
gt2_rxphalign_i                              <= tied_to_ground_i;
gt2_rxsyncallin_i                            <= rxmstr0_rxsyncallin_i;
gt2_rxsyncmode_i                             <= tied_to_ground_i;
gt2_rxsyncin_i                               <= gt0_rxsyncout_i;
gt3_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt3_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt3_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt3_rxphaligndone_i,
        DLYSRESET                       =>      gt3_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt3_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );
gt3_rxphdlyreset_i                           <= tied_to_ground_i;
gt3_rxphalignen_i                            <= tied_to_ground_i;
gt3_rxdlyen_i                                <= tied_to_ground_i;
gt3_rxphalign_i                              <= tied_to_ground_i;
gt3_rxsyncallin_i                            <= rxmstr0_rxsyncallin_i;
gt3_rxsyncmode_i                             <= tied_to_ground_i;
gt3_rxsyncin_i                               <= gt0_rxsyncout_i;
gt4_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt4_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt4_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt4_rxphaligndone_i,
        DLYSRESET                       =>      gt4_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt4_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );
gt4_rxphdlyreset_i                           <= tied_to_ground_i;
gt4_rxphalignen_i                            <= tied_to_ground_i;
gt4_rxdlyen_i                                <= tied_to_ground_i;
gt4_rxphalign_i                              <= tied_to_ground_i;
gt4_rxsyncallin_i                            <= rxmstr0_rxsyncallin_i;
gt4_rxsyncmode_i                             <= tied_to_ground_i;
gt4_rxsyncin_i                               <= gt0_rxsyncout_i;
gt5_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt5_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt5_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt5_rxphaligndone_i,
        DLYSRESET                       =>      gt5_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt5_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );
gt5_rxphdlyreset_i                           <= tied_to_ground_i;
gt5_rxphalignen_i                            <= tied_to_ground_i;
gt5_rxdlyen_i                                <= tied_to_ground_i;
gt5_rxphalign_i                              <= tied_to_ground_i;
gt5_rxsyncallin_i                            <= rxmstr0_rxsyncallin_i;
gt5_rxsyncmode_i                             <= tied_to_ground_i;
gt5_rxsyncin_i                               <= gt0_rxsyncout_i;
gt6_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt6_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt6_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt6_rxphaligndone_i,
        DLYSRESET                       =>      gt6_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt6_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );
gt6_rxphdlyreset_i                           <= tied_to_ground_i;
gt6_rxphalignen_i                            <= tied_to_ground_i;
gt6_rxdlyen_i                                <= tied_to_ground_i;
gt6_rxphalign_i                              <= tied_to_ground_i;
gt6_rxsyncallin_i                            <= rxmstr0_rxsyncallin_i;
gt6_rxsyncmode_i                             <= tied_to_ground_i;
gt6_rxsyncin_i                               <= gt0_rxsyncout_i;
gt7_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt7_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt7_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt7_rxphaligndone_i,
        DLYSRESET                       =>      gt7_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt7_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );
gt7_rxphdlyreset_i                           <= tied_to_ground_i;
gt7_rxphalignen_i                            <= tied_to_ground_i;
gt7_rxdlyen_i                                <= tied_to_ground_i;
gt7_rxphalign_i                              <= tied_to_ground_i;
gt7_rxsyncallin_i                            <= rxmstr0_rxsyncallin_i;
gt7_rxsyncmode_i                             <= tied_to_ground_i;
gt7_rxsyncin_i                               <= gt0_rxsyncout_i;
gt8_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt8_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt8_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt8_rxphaligndone_i,
        DLYSRESET                       =>      gt8_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt8_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );
gt8_rxphdlyreset_i                           <= tied_to_ground_i;
gt8_rxphalignen_i                            <= tied_to_ground_i;
gt8_rxdlyen_i                                <= tied_to_ground_i;
gt8_rxphalign_i                              <= tied_to_ground_i;
gt8_rxsyncallin_i                            <= rxmstr0_rxsyncallin_i;
gt8_rxsyncmode_i                             <= tied_to_ground_i;
gt8_rxsyncin_i                               <= gt0_rxsyncout_i;
gt9_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt9_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt9_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt9_rxphaligndone_i,
        DLYSRESET                       =>      gt9_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt9_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );
gt9_rxphdlyreset_i                           <= tied_to_ground_i;
gt9_rxphalignen_i                            <= tied_to_ground_i;
gt9_rxdlyen_i                                <= tied_to_ground_i;
gt9_rxphalign_i                              <= tied_to_ground_i;
gt9_rxsyncallin_i                            <= rxmstr0_rxsyncallin_i;
gt9_rxsyncmode_i                             <= tied_to_ground_i;
gt9_rxsyncin_i                               <= gt0_rxsyncout_i;
gt10_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt10_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt10_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt10_rxphaligndone_i,
        DLYSRESET                       =>      gt10_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt10_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );
gt10_rxphdlyreset_i                          <= tied_to_ground_i;
gt10_rxphalignen_i                           <= tied_to_ground_i;
gt10_rxdlyen_i                               <= tied_to_ground_i;
gt10_rxphalign_i                             <= tied_to_ground_i;
gt10_rxsyncallin_i                           <= rxmstr0_rxsyncallin_i;
gt10_rxsyncmode_i                            <= tied_to_ground_i;
gt10_rxsyncin_i                              <= gt0_rxsyncout_i;
gt11_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt11_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt11_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt11_rxphaligndone_i,
        DLYSRESET                       =>      gt11_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt11_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );
gt11_rxphdlyreset_i                          <= tied_to_ground_i;
gt11_rxphalignen_i                           <= tied_to_ground_i;
gt11_rxdlyen_i                               <= tied_to_ground_i;
gt11_rxphalign_i                             <= tied_to_ground_i;
gt11_rxsyncallin_i                           <= rxmstr0_rxsyncallin_i;
gt11_rxsyncmode_i                            <= tied_to_ground_i;
gt11_rxsyncin_i                              <= gt0_rxsyncout_i;
gt12_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt12_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt12_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt12_rxphaligndone_i,
        DLYSRESET                       =>      gt12_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt12_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );
gt12_rxphdlyreset_i                          <= tied_to_ground_i;
gt12_rxphalignen_i                           <= tied_to_ground_i;
gt12_rxdlyen_i                               <= tied_to_ground_i;
gt12_rxphalign_i                             <= tied_to_ground_i;
gt12_rxsyncallin_i                           <= rxmstr0_rxsyncallin_i;
gt12_rxsyncmode_i                            <= tied_to_ground_i;
gt12_rxsyncin_i                              <= gt0_rxsyncout_i;
gt13_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt13_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt13_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt13_rxphaligndone_i,
        DLYSRESET                       =>      gt13_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt13_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );
gt13_rxphdlyreset_i                          <= tied_to_ground_i;
gt13_rxphalignen_i                           <= tied_to_ground_i;
gt13_rxdlyen_i                               <= tied_to_ground_i;
gt13_rxphalign_i                             <= tied_to_ground_i;
gt13_rxsyncallin_i                           <= rxmstr0_rxsyncallin_i;
gt13_rxsyncmode_i                            <= tied_to_ground_i;
gt13_rxsyncin_i                              <= gt0_rxsyncout_i;
gt14_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt14_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt14_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt14_rxphaligndone_i,
        DLYSRESET                       =>      gt14_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt14_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );
gt14_rxphdlyreset_i                          <= tied_to_ground_i;
gt14_rxphalignen_i                           <= tied_to_ground_i;
gt14_rxdlyen_i                               <= tied_to_ground_i;
gt14_rxphalign_i                             <= tied_to_ground_i;
gt14_rxsyncallin_i                           <= rxmstr0_rxsyncallin_i;
gt14_rxsyncmode_i                            <= tied_to_ground_i;
gt14_rxsyncin_i                              <= gt0_rxsyncout_i;
gt15_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt15_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt15_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt15_rxphaligndone_i,
        DLYSRESET                       =>      gt15_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt15_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );
gt15_rxphdlyreset_i                          <= tied_to_ground_i;
gt15_rxphalignen_i                           <= tied_to_ground_i;
gt15_rxdlyen_i                               <= tied_to_ground_i;
gt15_rxphalign_i                             <= tied_to_ground_i;
gt15_rxsyncallin_i                           <= rxmstr0_rxsyncallin_i;
gt15_rxsyncmode_i                            <= tied_to_ground_i;
gt15_rxsyncin_i                              <= gt0_rxsyncout_i;
gt16_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt16_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt16_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt16_rxphaligndone_i,
        DLYSRESET                       =>      gt16_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt16_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );
gt16_rxphdlyreset_i                          <= tied_to_ground_i;
gt16_rxphalignen_i                           <= tied_to_ground_i;
gt16_rxdlyen_i                               <= tied_to_ground_i;
gt16_rxphalign_i                             <= tied_to_ground_i;
gt16_rxsyncallin_i                           <= rxmstr0_rxsyncallin_i;
gt16_rxsyncmode_i                            <= tied_to_ground_i;
gt16_rxsyncin_i                              <= gt0_rxsyncout_i;
gt17_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt17_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt17_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt17_rxphaligndone_i,
        DLYSRESET                       =>      gt17_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt17_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );
gt17_rxphdlyreset_i                          <= tied_to_ground_i;
gt17_rxphalignen_i                           <= tied_to_ground_i;
gt17_rxdlyen_i                               <= tied_to_ground_i;
gt17_rxphalign_i                             <= tied_to_ground_i;
gt17_rxsyncallin_i                           <= rxmstr0_rxsyncallin_i;
gt17_rxsyncmode_i                            <= tied_to_ground_i;
gt17_rxsyncin_i                              <= gt0_rxsyncout_i;
gt18_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt18_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt18_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt18_rxphaligndone_i,
        DLYSRESET                       =>      gt18_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt18_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );
gt18_rxphdlyreset_i                          <= tied_to_ground_i;
gt18_rxphalignen_i                           <= tied_to_ground_i;
gt18_rxdlyen_i                               <= tied_to_ground_i;
gt18_rxphalign_i                             <= tied_to_ground_i;
gt18_rxsyncallin_i                           <= rxmstr0_rxsyncallin_i;
gt18_rxsyncmode_i                            <= tied_to_ground_i;
gt18_rxsyncin_i                              <= gt0_rxsyncout_i;
gt19_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt19_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt19_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt19_rxphaligndone_i,
        DLYSRESET                       =>      gt19_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt19_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );
gt19_rxphdlyreset_i                          <= tied_to_ground_i;
gt19_rxphalignen_i                           <= tied_to_ground_i;
gt19_rxdlyen_i                               <= tied_to_ground_i;
gt19_rxphalign_i                             <= tied_to_ground_i;
gt19_rxsyncallin_i                           <= rxmstr0_rxsyncallin_i;
gt19_rxsyncmode_i                            <= tied_to_ground_i;
gt19_rxsyncin_i                              <= gt0_rxsyncout_i;
gt20_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt20_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt20_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt20_rxphaligndone_i,
        DLYSRESET                       =>      gt20_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt20_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );
gt20_rxphdlyreset_i                          <= tied_to_ground_i;
gt20_rxphalignen_i                           <= tied_to_ground_i;
gt20_rxdlyen_i                               <= tied_to_ground_i;
gt20_rxphalign_i                             <= tied_to_ground_i;
gt20_rxsyncallin_i                           <= rxmstr0_rxsyncallin_i;
gt20_rxsyncmode_i                            <= tied_to_ground_i;
gt20_rxsyncin_i                              <= gt0_rxsyncout_i;
gt21_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt21_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt21_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt21_rxphaligndone_i,
        DLYSRESET                       =>      gt21_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt21_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );
gt21_rxphdlyreset_i                          <= tied_to_ground_i;
gt21_rxphalignen_i                           <= tied_to_ground_i;
gt21_rxdlyen_i                               <= tied_to_ground_i;
gt21_rxphalign_i                             <= tied_to_ground_i;
gt21_rxsyncallin_i                           <= rxmstr0_rxsyncallin_i;
gt21_rxsyncmode_i                            <= tied_to_ground_i;
gt21_rxsyncin_i                              <= gt0_rxsyncout_i;
gt22_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt22_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt22_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt22_rxphaligndone_i,
        DLYSRESET                       =>      gt22_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt22_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );
gt22_rxphdlyreset_i                          <= tied_to_ground_i;
gt22_rxphalignen_i                           <= tied_to_ground_i;
gt22_rxdlyen_i                               <= tied_to_ground_i;
gt22_rxphalign_i                             <= tied_to_ground_i;
gt22_rxsyncallin_i                           <= rxmstr0_rxsyncallin_i;
gt22_rxsyncmode_i                            <= tied_to_ground_i;
gt22_rxsyncin_i                              <= gt0_rxsyncout_i;
gt23_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt23_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt23_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt23_rxphaligndone_i,
        DLYSRESET                       =>      gt23_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt23_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );
gt23_rxphdlyreset_i                          <= tied_to_ground_i;
gt23_rxphalignen_i                           <= tied_to_ground_i;
gt23_rxdlyen_i                               <= tied_to_ground_i;
gt23_rxphalign_i                             <= tied_to_ground_i;
gt23_rxsyncallin_i                           <= rxmstr0_rxsyncallin_i;
gt23_rxsyncmode_i                            <= tied_to_ground_i;
gt23_rxsyncin_i                              <= gt0_rxsyncout_i;
gt24_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt24_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt24_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt24_rxphaligndone_i,
        DLYSRESET                       =>      gt24_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt24_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );
gt24_rxphdlyreset_i                          <= tied_to_ground_i;
gt24_rxphalignen_i                           <= tied_to_ground_i;
gt24_rxdlyen_i                               <= tied_to_ground_i;
gt24_rxphalign_i                             <= tied_to_ground_i;
gt24_rxsyncallin_i                           <= rxmstr0_rxsyncallin_i;
gt24_rxsyncmode_i                            <= tied_to_ground_i;
gt24_rxsyncin_i                              <= gt0_rxsyncout_i;
gt25_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt25_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt25_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt25_rxphaligndone_i,
        DLYSRESET                       =>      gt25_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt25_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );
gt25_rxphdlyreset_i                          <= tied_to_ground_i;
gt25_rxphalignen_i                           <= tied_to_ground_i;
gt25_rxdlyen_i                               <= tied_to_ground_i;
gt25_rxphalign_i                             <= tied_to_ground_i;
gt25_rxsyncallin_i                           <= rxmstr0_rxsyncallin_i;
gt25_rxsyncmode_i                            <= tied_to_ground_i;
gt25_rxsyncin_i                              <= gt0_rxsyncout_i;
gt26_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt26_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt26_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt26_rxphaligndone_i,
        DLYSRESET                       =>      gt26_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt26_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );
gt26_rxphdlyreset_i                          <= tied_to_ground_i;
gt26_rxphalignen_i                           <= tied_to_ground_i;
gt26_rxdlyen_i                               <= tied_to_ground_i;
gt26_rxphalign_i                             <= tied_to_ground_i;
gt26_rxsyncallin_i                           <= rxmstr0_rxsyncallin_i;
gt26_rxsyncmode_i                            <= tied_to_ground_i;
gt26_rxsyncin_i                              <= gt0_rxsyncout_i;
gt27_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt27_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt27_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt27_rxphaligndone_i,
        DLYSRESET                       =>      gt27_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt27_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );
gt27_rxphdlyreset_i                          <= tied_to_ground_i;
gt27_rxphalignen_i                           <= tied_to_ground_i;
gt27_rxdlyen_i                               <= tied_to_ground_i;
gt27_rxphalign_i                             <= tied_to_ground_i;
gt27_rxsyncallin_i                           <= rxmstr0_rxsyncallin_i;
gt27_rxsyncmode_i                            <= tied_to_ground_i;
gt27_rxsyncin_i                              <= gt0_rxsyncout_i;
gt28_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt28_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt28_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt28_rxphaligndone_i,
        DLYSRESET                       =>      gt28_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt28_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );
gt28_rxphdlyreset_i                          <= tied_to_ground_i;
gt28_rxphalignen_i                           <= tied_to_ground_i;
gt28_rxdlyen_i                               <= tied_to_ground_i;
gt28_rxphalign_i                             <= tied_to_ground_i;
gt28_rxsyncallin_i                           <= rxmstr0_rxsyncallin_i;
gt28_rxsyncmode_i                            <= tied_to_ground_i;
gt28_rxsyncin_i                              <= gt0_rxsyncout_i;
gt29_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt29_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt29_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt29_rxphaligndone_i,
        DLYSRESET                       =>      gt29_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt29_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );
gt29_rxphdlyreset_i                          <= tied_to_ground_i;
gt29_rxphalignen_i                           <= tied_to_ground_i;
gt29_rxdlyen_i                               <= tied_to_ground_i;
gt29_rxphalign_i                             <= tied_to_ground_i;
gt29_rxsyncallin_i                           <= rxmstr0_rxsyncallin_i;
gt29_rxsyncmode_i                            <= tied_to_ground_i;
gt29_rxsyncin_i                              <= gt0_rxsyncout_i;
gt30_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt30_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt30_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt30_rxphaligndone_i,
        DLYSRESET                       =>      gt30_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt30_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );
gt30_rxphdlyreset_i                          <= tied_to_ground_i;
gt30_rxphalignen_i                           <= tied_to_ground_i;
gt30_rxdlyen_i                               <= tied_to_ground_i;
gt30_rxphalign_i                             <= tied_to_ground_i;
gt30_rxsyncallin_i                           <= rxmstr0_rxsyncallin_i;
gt30_rxsyncmode_i                            <= tied_to_ground_i;
gt30_rxsyncin_i                              <= gt0_rxsyncout_i;
gt31_rx_auto_phase_align_i : gtwizard_0_AUTO_PHASE_ALIGN    
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt31_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt31_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt31_rxphaligndone_i,
        DLYSRESET                       =>      gt31_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt31_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
           );
gt31_rxphdlyreset_i                          <= tied_to_ground_i;
gt31_rxphalignen_i                           <= tied_to_ground_i;
gt31_rxdlyen_i                               <= tied_to_ground_i;
gt31_rxphalign_i                             <= tied_to_ground_i;
gt31_rxsyncallin_i                           <= rxmstr0_rxsyncallin_i;
gt31_rxsyncmode_i                            <= tied_to_ground_i;
gt31_rxsyncin_i                              <= gt0_rxsyncout_i;

    rxmstr0_rxsyncallin_i   <= (gt0_rxphaligndone_i 
                                          and gt1_rxphaligndone_i
                                          and gt2_rxphaligndone_i
                                          and gt3_rxphaligndone_i
                                          and gt4_rxphaligndone_i
                                          and gt5_rxphaligndone_i
                                          and gt6_rxphaligndone_i
                                          and gt7_rxphaligndone_i
                                          and gt8_rxphaligndone_i
                                          and gt9_rxphaligndone_i
                                          and gt10_rxphaligndone_i
                                          and gt11_rxphaligndone_i
                                          and gt12_rxphaligndone_i
                                          and gt13_rxphaligndone_i
                                          and gt14_rxphaligndone_i
                                          and gt15_rxphaligndone_i
                                          and gt16_rxphaligndone_i
                                          and gt17_rxphaligndone_i
                                          and gt18_rxphaligndone_i
                                          and gt19_rxphaligndone_i
                                          and gt20_rxphaligndone_i
                                          and gt21_rxphaligndone_i
                                          and gt22_rxphaligndone_i
                                          and gt23_rxphaligndone_i
                                          and gt24_rxphaligndone_i
                                          and gt25_rxphaligndone_i
                                          and gt26_rxphaligndone_i
                                          and gt27_rxphaligndone_i
                                          and gt28_rxphaligndone_i
                                          and gt29_rxphaligndone_i
                                          and gt30_rxphaligndone_i
                                          and gt31_rxphaligndone_i
                                    );

end RTL;


