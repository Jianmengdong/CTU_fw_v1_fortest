

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
RyffiulBG9yray92XSWIlgI2WAetX/UVC+q0Z7efs5TjeyYMALW4MUyGitOBiAYlCSTOM1vVAHPW
Dyw82okGLQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
rimQZJKtQGQJzltFhJXAQIKTKEPCr0gmY8hUnpX7foRCR3gurN5OGiG2zPFxPkvg7BDCy3mbele6
Xt6kIVrlKZ4dJ41V49F7Wd0tgbjqJ4yZGzrKV9H/LfuMDgukGDBTwP8pmUBpqAt5LhElrr7DvLd5
DJ6THnbvDKdUBOxbUJs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hKY0JBzbgea8xWVR3hiXbbfwid6oBYVk1H6bQjlx2c/4Igf19PYjaI2u4rwfGsxORD6rR+CKl5sV
nPqykldAQz4eBJ9HC4cRHG5+TE3tA6PJatXqkWsUfOg7DASqjGxJQm+nUcdbaJocCoQQ6aFn7dTM
uoh4DGLg3SfaDQ6A4m8Ykcl7qdAJMhV8LgYbwKVE84BRieVyPNL2kjlSXhMAq9wJqt3aTFpbjAi3
cri4+eL//e4NxqoIM24Im7QkUCkt5LNGP62V4HYf/K1ZcR8Pd0YE/OsGW5Mww4xgW62NgpWn0cwK
IJo9x/J6vCMukKeLZTXsjyLsOPvckv59xk69jw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Br6ZvKm4NdT2KtaRiamSTouR9wa1QvLdMENyXsKqZTUYQ1NpYAREbFc/p0DTCJ6ZIVDwzvFERR9F
uBqjQznay5KRzam7DXASIunRpreYPFSI8lweGk0i5aehcu4sANrxGO0nhhMFz17XAK4eFuLLuIcb
tZVI40jAT/WnNUp7/0mk3Pqzn6Rptt6OYMdtQ3rV0zJhWyGWBxYKKWDGaz+bdf67UYutsrLwRyOe
+nSz1iBQDsZkHOfk/OZzUgPfwU+XaE47O0j+dcCHD8HGNZ5+rSyIjDaz6jICuM8LROQnEqMjrNqE
8PMJJln8b/v5LiPve2M1AAGUPAcu1J3N9PWzvQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GuHEPjnAcllqBAw9XE0/C9vDbSQfiKB7BuymJyg9A62rWf77qd/mZohqEvbem3QrLXwjOoWnMEJZ
6esdv+RuxDyNjIvX+5zcKtM3tg/YelhyW5Yrs3erpq7/+3wE36q4KohHlk8NBUHD99Drl6DCl/+v
tfP1tCSgJtRa8ap4Cstxhjzn5HK3frc/YrST5QSRjwjCmlih0zwAEmbom7XmxAdI0AW1cotQCkoN
VXWJ9d7uvDTGLsvN+cxzH5xh5kiyIfwp6SXB0VK2HmiMSOACKKlNg/FAQs2jMLZjgyEznB+QkBpQ
8fL0EeFT/cgXquJJ5t8uN4xWp1CCWsMm3CpRyA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VNIVki8CRk9kWGG4smtEjl4elbfSt2tJqXpkbDnTTkhlJw5SQufV0hJtqG3ygtXATOrMwTtwlJcw
wBW/gSpWV0rnBKfcLzSBLmKm38GFHG+K+cEcY0fuyfm7bp0DP1Mn5AgsttDG9Jg4wUwPiXCVa0Kb
BRqKewRQbIIPXNdYuQg=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
d8lIT6H7Vyn4rBnYvZVeSmqj/ZK923mpNqmvpP5ASvOloylHeh2+kEoElQkZiNxU07Q84uZerDNy
wWriOG+DDFNx5KvUWWR7CbUJoYuE4npSGYK/rlPA7NkaBe+QeM2qGwTfJB3xl0LehoIuswHavS9B
562mduZP7nhcXIK7mIdTsN9bhOUsi5W8ZRMKmRvLAxqwbAFK6m6yx8CoUkVdIQ0gnBvTAAFTPFuG
ariOqh83aKdsZn17Q+xW9k4sdvddp3DVuo8woscCM6ERlIcvcJiAw+gqBNdgGd3hs0m0eNgk2l+j
wrEJN533dkz1/3kxa+HAlZIWmPC+3IYXHbhMjw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74224)
`protect data_block
r4Dwo6nL2e5tjgrph2ZPYQznWTDEr9AFhBSOHMyMLbYuDKYVcqikJY4N8Rq4xZTzFm/5TqQx5DTO
R+28YaEVE/4odx3juFUAPU6rjQJbllmkig6dkltq0zSLHYo3DDmPFfEDiDW2vGItgoQ3/xxmPxsH
2j1gT4DK3RpU9KONc2EsWjrAm14hSuN3TKBimmveIL3MldI+OWDYeo+VW/wnhYFR5dpNoF2oL1Qc
dz1JL01UrKHODeZSlR36B1ceyXA1OiCNsPjRuiC//NR/39tVA9e8gCRYT2Xc/88XMk+ReI7S00ug
li0lUxcK5YiLOKfj00o8GSS1C59YuGvxwONGGeYUpFqPCpxsmKNwZDv5poD55zkuX9tVFfza56zr
QmF5vQopN7HC6LCiC6nlVE5IJ+NclknOPDGB5WizhEhFvjRF7uKGOzjOwjFY85xlKFeWAaSJV9vs
/BJ25YvgOHAbTEcLl4W+hZZivyLBbyZFTrywHfSiZ4g0leMwP7pI3cllEN3vWH7Ydpc5n4nyEGHG
y7qL23Je5yeIpr2KiKoidgPEkyTl2z3vUezG0e1zTlmlq2MPumNY6YSWAyLRaatYtBJ6XKc+WIBk
pSRJ1RMUAYs7EJkSCL4qS93BLLyrYRT/11KTJ3de/rjuacsrHmLqzbMtED21ME/iFS0cX/tEjp/1
dKlzNVU6IBEoIiBL0MA3RkPumf5Y4iSvjlXr3g+1xRPaTR538288Ixi7Y6cIux678JRloRBshK7H
0uXMmMDj1wnotY9gQ009uEv6v/DTOzyc+ARVZEJDVDAqVDNwY7nvHQYjnr17zB+DL0JCpJE0hpgD
w1x+hRgghMMQsY+LQ7b94PhBkMsNcKIa9yS8UDlBEliUpeCT5AnPqWGbFxUrfOxMmBWRYX3uWSTu
7WjL8fnX1RYH4aYJugPQp68GQSoW5MIY5y/r+vADjYOFF748xwQ/rpXtbdV8UKOMeHoIcqsUOYYI
vwygzu/coPar0NiB1ygjYU36TtKagyvdbgI81VR6z5R4mZ+Ns45zk/zS0WJ/wTqy992gxwsI9lls
SHpJCZ7V1YLx6OQYxgfuHyDqrmfCwWzc3bQ69fAt9kPw9K0RO9vxvAiXiK05R0XkX0ourq2NUo7a
7xnPP9o03gg16h6BwdD5Tdg8ymg6FWKSAVi87+2CF+kHP7BPpfhnksWyO7jvdI7dhCYtOK9irNMz
mXUub4eQ0qP1ZdVPGxuoEvrtS0xKQ4Uia1puYoVogBsXHWZt/40pP/8mdBEW7Y5ACBN4tGnux+MX
i29nB2Aej8IBrbZbd8Nhscg2dv/0bwYfe7vPWbCP2WJDGzYtA3lQgHhxKJ6zHSH8NCpHxSThzR/c
PRPzLxyLtDfzDoVTfc1R/uzm6JdvDoYMajlPwMB1JhK4olR3p6zpi+oBkuhnLnhASNGIlyEkYaWt
LRNhUxm6XSDFcP+qZG+TaMVGVmIR5wiGsRF8xpFSLXoNoZ6GrUj7iUBEa6ECQIpro0v4Jl3qprF1
0THt3jY82iuGW329+3y0WwrdHgnAbzm5HklkHm947wxXHPaTrTmMdHzPak9tJCE/3NRjY1WAfOgg
wTPdW8ljnHUPQeEuJLwwrp6FOivArkydoIBwW9kHxRrYP2YKOHoiqYd1vdVP1PGzSmSRk4WkNdqT
35VF2IHsQptFROdgCmTpOkAQswL3u8SGmlhEUhrm565dWYxEVnJEKExBXDYtU0zwk6GoqYqdKhO9
baxfohOGDqHpdqiEKzRWyQZIb+4WgKC5xYPeseA3UMqtc5y4B3dVIFKGdZouTyKe8TPLFlPV+Xvw
AAUVXPW4XwOxO+7vcU7b6+nJaU0K08LsIrj8IJD4mOMM1kuWvl4/ULobKqUKBo0NdqQiV4hxR1Vu
RMnZqH4kFQcaPfwq9u6x8QW5Qq1XLphWQiwVmRG7oy2ArI9BumiHFLAhMUqGhIZd5PKkDBJ6g0cs
cAul2/N6zxZIs6GSfF8OWrUy3oGqdKg/Lrz9F3JwzHjdUNnFg6oy7c50XXeYG3U3lRCUGRfNZoMo
ikimMTAUSyWNZEwqPHtrQKovDk5/f0dLJur8OVdXcafGYkFvPRiKsWHL7yxxMBV30pHE9UG6DKL+
c5+/7BUpwaP9hH+zQMJ3TFNl+16NkY9UKzsW3D6VcXelHbMAg14jqZx/smzTrd/8biI47ma1uAg1
AOCbvLPwroeMt9uVSlI9TtADhDyQURnSwqPR7Wmg6BPv195Ow9VEBLZxQAx0yP5vhFymKK6WFwHH
m3XiqBfBxbFFZ9jjZypRz4vtMSnZOUOYUu5Z2oDe3Dwq4RK6e7pk9hiWIfGICsiCm/3dvsj+0bND
0ltBk5TOtpAs6aFVgKQ//0lMe+Zk36z/AVHEEamhkQc9I9SGXxM9187gEpvdE94KYP7LxYMcO7uy
5tTIwDOYjr0CJhJDZtZ4nzKAM71sgxH1359fqw9WcXKkOCLklnc4OJ+oLtgkrU6WBw61WrroGdD3
QB94PRwWqs4ArNhEq79MIqe0l0BdA4xFNYogHQoWamRCdsPVKzhqu5ES/e0IxyuMvXuTK0+ZDmmU
nvi+yuqW2NbZV0TbYOvQuogxu4D4PmITLRQaU9XxgkEA801K1TG/Zy+CjbZv4otWU9oey72YqlOe
7QscS0mRLiVHatvBoJvTlzZDNLxDltnoJpBM10Klcfp4hp1/2X04vkLactLt1ohNvpGt30P+Ray/
xYcgbTbw6c2zjCyHrvjoLKcbJy+0i4+FJg9GQdeiRZscAUpXruj2NEG6y+UR/9EsDGIjFmMeSPSo
bDbHFYUjmDEkPbWW0LLSFcB5S8e5VGj4I7o/0Qw1a4W1bzHmfEpJZhNqv9TI8aHFaNEzxnXKZ1RX
BSaOAinA1LEOv0keblUAkO9YAHpF+mqwIu1oFsjhoKDOT0lwCxP8f7RxqlZJhLbEll2NGjzB/bxl
SIMFkfsIxn/fdPmM71mM4bv9+cp7XjerrpKVula8tk5hZfpoKcRhFVp8xa2q315FfKK5sH7hMXON
QVrncwoVM5Gs7ItIcZnsrl0r8ZxrSYEoaakf+8N8noqVkWQ0RJc14QySwhYoxO6SuO8v4l5zbyzf
G0/dhwRkHqWDp6XjRW85C/82hdko4l0LNXIvgV3JyLO/4f9MNUTf6W+4mlhHv/kBJILvFTXTGyVf
yBMWx4alQGuv3qjS5nnKUfu+ouHlvZTm5NfuMXQf4/qhR1Jas/6BKE8hZ+SaoXMWUwodHUWxGiyk
FdaL8oDk6OghM6lL+SNUvpfR4VSf9YL96fYgiZDr2QtSTp6Kfb3QZSm9nXl+ukEIzaLys8c1iCPT
yFQ7Qq8xPmX0vfkaoexdWdRxXrareOkjkeaBfSX5m8IPR8lss89tRatBAKfC+uzM80nmUtO39m0h
LJ34b90jHOhOq7L46UGACdBl3iTlxJJYAQRGDD94v/XbNla92SQmNRtK2ftoklFgxkNw6az5BTst
vZ336ZhTU4JG5rSmPYbMlHEq/GKD1NNuMQhGi1x+NtBv5GIwUAxIvuAuxBxN27SI9qPe3odUklbU
a+rZoeMrbrw1FsjGJ1QYvSxZPHgHtJ89j81tbQFD2FzNxNTlkIjTI2JUZI/pSc43ceZcb3F3ugRn
t7swQQMHb90Yf1MVlSKITneMsaHpMYhx33hgA35jeffBpnIiCYWJnA/C0lFgjGZtxKq7/WCPHYL2
rLOSN68R0yzno57IrtJJ20QA1op/BS9mRhDCR4jt+v7yX8lkVUMjJpxzE8JokmyLyxNYv/U+roYQ
b9HwvtmIrV+NUQi/SRfXN2gZzA3ezm+7Lcb53CorbgPlCwTC1ISw1kUiNqalGwWoBzSKqGJ3nRuP
lirp6b0e76kV55RQdHM1K/MqmQCaN1gddL1mkiqP7hnJaJm/bwNTxr+PhoEA1jU244Pd2YxQev3r
iIrRniXKw21JzXdS9Dbqv7fJ9XFjwuWh6yf/LbCpFcsrPsYFPkV4GDAfe2pea5F3G1sIquGRzSvE
eILRH69s7gwBhvzl/5sv3tSVxD+aTINk/q3aL7/ogG2FRMX1GTC7g/n+ux76HDYfuJusDcXLxILx
QgTfGd2n3g3yWtN7cMYj2kII/wAhqVaRSonP8byC3zO+tRwuHnoa4fFe1hCgxhlu8BPzqYhdni1O
9CpGXvXAPcT7htR6JnTS7CDvoufOyc+H/inwN6toCBXEA1ej3B/HnNv6xhL2hbL5i9zvyqEAjLA9
/ApBc3OPo1lnnomQH5WnuH4OfUHjjWwqVa+o387XFln3mVg9BTpwEsPTGi6AUd0O6TE+hLUd1dwP
8k5+a0deRpGiN07i9g2nNCkH/Nng8lTW0uN9idQbf6SPVm3tAz/5Utwu+8IrdOntI265s+vqrBme
KHwyIi5A7d/Xsw7x8r2zwP1tjr2SiWj3tsJVQiJ3ae/jO5f1uAMwBtRHv1so29JQID/BS1KhKfQ2
+N8JmHEuAba3p2GCDDvcUEvoqSI7rcmEXMeQ7goOU0SUV2JEiO76nO2VpciBqzfjFlbEV0/TiwyJ
vvUGFcIv1iti6FpGp2bjPuIdpB4H9P1RfnXmW5Ae5DF58Z8xUQMhtIEuBsv4SenAJNfxVO7Ukuax
eSRfaMhE8EBWtPdPjjvUKRLhQjitma9LRgykhJUfQASMkXo6ZqQnJW3w5BbJ6lD4ZnbnmoCJbWSi
hfcJSrAuzydhrPOB8Sh9PfGTwFNSOeNGq2HVlToYZwaO+KXvE00IJ0SYJCtXS2Dxh8cSVX3flEPG
usJkUUYaH//JclSXuwIxd+nLQiqnqy1O/qX5TaY1H59bE3aO2pFNS+M/VQiTa+5s6w0szgFByea6
Sal4oBv7zFDXYIFKeNGejbEmen0rL3tNr+k0nOdpsH39t0i6lSAg6FPiQLSy4AbFydZ0HiZq8xTm
S85OYUYDdmuzhzQZLDx4ce1rysO3E8dDUxMS2UKqWvHpzfUS6qOn55DzAN+Y23eBk6YSg8SQvzwL
YUkvAdCQvNfHjCvBdvVIxHk+h4RyU8LYD8fxvuTw548XDS8AGcxLS3eOz7UskBWPrV/sUHf50Oj3
kqQbvXjeatEkj11ikndaqSWVefsX9S7qycv2trF042fQPXqPGg7sv1ueKjxX3bTENBJk6dXFshZF
BVd3fPzuErCFZGPg6e+sdhAw/FsHctkE7PfLeMqebYFvuf+NtIcYQN9QfJcoJQcGCG3EpxFtphpz
daFQ1Q0Lr21Ql7/qlqVZIgcRhI+kSI4I+zP5MRN5n+HRG+2FeiH2Vp3fyoTlM0Kif5WEMLdkzFYS
UWYwaCulJVPkm1FUG0MleLlDR2wSOdwNzXxiAWuobVVJgHoVq/YxAHMpFS6+PmblJMfVTt+UZ/Au
QcBrQOMII9qug9F1xEM5fiDdh12J5rXSWUPRoX4VwVwNQiJWs9g8O3hmkkUWbqvTzDVNebVpRyf4
dXb1Jz9pRtBUc7S9EYXz6h5r/HDkaYfoHUxqC+7JopMQ0zSQjlRU1+LUEvlYtLHIWoAN3OLzW/G+
bXmeV6KhC3Rr/bUYMlOBxLMw6iRa+IQu/Zp8l6MWEaHg1ky9e4aFJTq/MaCHHHOunF6szyLH9IiI
e4BWYKUVWoos5UJYe4jtcO29CSRVDtKELvvGYCygRlsMY1VLrwpz5cnFeU7/hL4+AXDnl6IW1Req
wi6kNY6Z2ZAGFB+TtbYiBDnGSiAcNf3Eq1cNMZBt2nMAW9GaFWaatl/dGmrcCOxqsiVnAyFKIO2Z
j73O755CU970osYrl1utEBr+n6E3/yzULc0CxB3cAZ1S1c74MeVctheU1u1H+WxthiyKFOZE5BIV
QQj1cI3XX9u2JrR13eWzTK9J2ejzfggWu3vBM6eROvrv9lidYuOkq25YPwo08E/58MH4g8RN9pJC
r3e30rNi8gEMsv+srLyaTgsM2ItMxkF7C5wISD0MQArH4sP0IOeb+lopnJNC/k+8scT4Rt/Bryci
71dFck4A4zik3829hqSQn9bVuOHfaAcLwWgojO8YwghVaUjBZF3VpjKExhMoG9dLh2UuTCGkeMIr
nJkHItLRGQ8Tj6GbdTmDCSH7YutMsT7B2OjYKvedQ/z6MJVImismgpEks0EN8wAu8diVdwOHYGjM
dtrc11IEhfq4I/4GreQ986ZgyVveON98ikwrDaSgOh0MVaqVFyJVaBdbq0Gvv6Vf2ykRww1zrRpl
55MBbMEUv3Bdu1I9tx0xCwX2Tl4CgGI46UR5Vh/uW77KJce6p/bEaSCWTkZMOUD9pxFzCkR0xHeb
WwnlDoLTt8cWU1heqWDSe2Os2L2HonXHuepEOCivqrfD9bn1/aVqjyHxmAsQb6p+PYKTF+OhBHi1
El2gY39f4gB6+4KKuIXD9TTj9kcUVcTGi+zad2v8/09381/RCVagnsUulzGvLfkUkQ8zcsG43dfn
24XROZCQtHeOEUWv3YV8giE6tfZuUeSWUN5gLrL9Fdsih11NiIfiZF8H8UhJyQ1qaH+vTOHyvfCD
70AKqmAjPjQPbI8ciT8Ad2btJbyRE3SEyj+jdwJpNrmv1dxOgeozTLFHMShgjwp0nAi61RirxHfE
xQp2qzF+Q+GJHreVT2XlZrybJ7dX+cyGqbmcFTr3ij8oKHD4a8/ZDX10MfW54Xh0Rj1PNz+25FYw
k9GUMTd9xG1dmcnonRH9NSv++pYhF+d+7rwghTY51lip4h66Sq/ps24AxzY2Dw5H7Fho1HRKkY0F
BD6/5IcVlMUUu/7c3xo0FzXNr2hawuGnmoxxIwrpff5NuXg7hJtGxHIKrKopo2DqKrnZHnzloVas
FdeEI3v5uyX4fXNxhlssI4Sr3JVv+ZeDOoqWxKkuZ3QDzxBBxGYRBwjZTUQQVMFDppgl75BPYWMp
UxYS0ehhdD5EZmJEHBvheW+sllcs43reav/Pn68L3vKPFvvIYAzZm2GvvHK6DiNGJMUZ1ZvfYdID
HycV0yv0cEEXjAPh1Pl74+fp2Zrvg/cFk2svzxbpxirrH5UvBWy4uDXbJcuYxCd21temGtkp34FA
n6ipbOoSYdHQbOyOQUTIeaGMjJcH0nT0XQkhWor/O5UWwAE8WzCmK91N6KAsg4ZT8ZJYsmCCWsKC
W9VZdTruGqy+ISkaPk742u49vwRyzT9mw0ep7q8fwyKSu53wJ4ibFvyCyxbY4xbJQ3TdpabSx8WQ
bL2TuutBxx+roVIzwq51wIh3yCXCP+pwbImHLuKlX5zcJ7dpN6OQ0zbo9kYLwaFYlOVPlIeHHM7g
3Q4g03Fc4tcnEPXfmvBEjkFHzhxOuRyrAlkBY9mC2aneafyyG0lI7+cFxxRx0aR5zHbsxSIxFBG1
6+hk91lS6fzkL80rzUOLVOB2aZCJp0h4aRetC7FfDAWd4Sz3EtZjbUpvPykv2/ug5hPsXkbrmw7q
+nuVn4jWJsL5G9gtm2WgU/SOwGmObTT9aCSKpwC8yExyrXptYmAcPbbHdKohqYcmr+7QfBCSru5l
w9AFr3uPIESDh1LRaSAVquLePOjGIzzhaeo/FdnsZNUU0hcv9+V5ESxU7irR0LCQ2uJN/G1mzYYf
OpcNXzOmtt0xVGU41iic9KNEhgOumfqTtvkYbn6CEme72Ceq+o+lnsjgZQ1YAN4XEiEqUSYnEwzk
Ml0rrFD4Td8G/mjz1NkshkY8Uno3DwEwdeEp7QVtD36U3qObdeBXOT1SD5H2VTDm1YiVoapjWk6Y
n5TDB1F6W2l+butKFKf4zotGz2rWt8aCyUl7B1Zt7llQAxUoA3zgs5HPvVox4a9oMMdizaaKHsB1
OMD7d06EFottlHvUa1qTswnvGScl/Dy1j3K+NOYBKBJdcqnoBsJWTkqeLlZJJGff2rYN5/lkU31G
Wot+1MGfNdHusYjQf1pet1ntBPzsk+9deGkKWEkLwVgD+FyI/quTgyD6RJzDFPI3A41l9Ao1OEJx
glQq7z73t9fDPzP2fDfkmRBZUaOIpBSFvoi580/9bwW0SKX4+Q+62frklwY0Fb7ygUP7r73RvR2L
2hmKH9edq1Bv+BabH5QoMEvemDQBw6GEyPsvr97VW8JXPSEyiP6J9iCCUSpPo7/pMMUCywbr4JUs
L49s4pT97u9e+XS75EmX/EaNofSsfM+pHBTahU+OT/9/nHR6nrJCqxOmx95cMwS64sE3l0rOx7LO
H2M14MNMhEIttOVoMvIGGVubaEVwUzCoLMouCiDJ9yNrL03TXFIfyhSkXG4nMJSh4NDcg2qjEYEn
0uovlQKZbHQ8ecBi6Pm7ZLilg6fmSr3TIQ21Q4bMa/v1p43+AoFrY0Q0/da4FX3xBj6vwIwCTc9L
sMqn2WlXQ2iwh6jnApP/Rpkzn7FQlArP2byA7Aq42rehEEAwcUJc+FraSv0aYJ7i+HP9DKheDLqf
yVG5XWu9VYedD4yNvEnfC4LZSEh0/+cilVaXhe626JwSBQ2zb8i8eb6P6/7NQxqslCVq8zwvjRyH
UdBbVV3C4BCzyc2p0cJsvnklc/YiBpy9iEpydKbffPWwCExLM8WtYZ/MNCFv54jEOL1zX1fX8M7c
tmd/qqNwFaiAYN7/C9KYBZCBeg55xGz5pzplMqDsBMdnECRm9AKUcgBbz1SaCaRGiI1etqECAcTq
+uOHdpKvARmQZN1mM3L2u9+iGalfIY0+rv0Dyv67wOSfm80eFBw5uQXYL+b4Z1PS+ZP05+XYKFIw
I9JS0hwSBg2K33YCamlNJFd6N1o1qSPQJA3FwJMeMaCk1ad4c0ijPH6uWLXhXlnBVgB0KQQJ9p8l
ZCSuFu+M8OTDyJje+n6qHmw9KabaU0RFW33h9tssgODp4WSo7BqCoNS3BLu4T5/X3eI8EsK0gn2c
8tdJAiVFdLTI9+rw2xlvcBHrDlWHK8VG0Td9cCV8+Ew5kIQYaQ8znSUfwTPEc8nya6dp26Xz0pPm
8lmHW/LArBuul20RKj4DGcj1P8wh7/aOkQNuq2xiR3wP9gYUTpSX6mwogKL/Ym40kqdAr2Kf/and
cXe1Fyu/7opGDZyj0oZkReflhDqZ9EfaJCvlaoSdsduV7BWO0qxO0v7C6ym+Y+krW2IvO72soEgg
pxq3ovbDBS6KxFZYL2h0TnrjyKkEKfCgNt37COiLLODt4pojrpU6he9yv0FjSmJOBHJkw1dO/7Id
1t9AGRmnMjVz4BjGYAhT4+W7dBDpweoL74LPAlcJgrLcHpIAsbOTnB/UQFpAe7Z3d8i9LCxOH6hr
7NAF+StIxLdgsBw7JR8Anh3kTpQ10nMdYj9NAa+RDFSUTeZ8uOAKdl05NRPDOjV/tA+ly4xF9ITU
ulzWOe0aFxPZDtY/T+ohAvcCYnG0f7WLeZFZPYJF+dWK7eSvig2XQoirxXxKAEk+dv8f/oEJ33Hj
0DDo0+x0jpc6VC4yDWyqkTFGYRqbqQQXVCMOuozMc/JwxpyIZ5U+3RMATykz2pJQBm4ByMcM35qo
dtTavhPJkM7zTJkDc3s4csIPNFOxE0LTgXgtuLx2z0dZIuFKDOP6ON6yC6wJQ6RkCfuJHo92FWpY
30v/elPolgx03g7SitSKa/E9PTtRwFYuwQATC53RLrO5A2bjJ8PzNZb7qDr3OhQhwRxewFAfPk5E
Wu8UPi/UX5WR8o/eMVkSOQiDUNoVLiWGqoX7F+8Z8xcWkr9bqa3Lghc3uBCwory7GddAhOGRah3/
d0gUYoietM0Rra7J8xBQLkSwvGiZLyz6s5vNWRj8CLWCFL7HZ4Rgn/LNchZ4oeGncHaVHeVnw6w2
X+gsE3oomwxC44w+TpXBOsM17N++okn6MSPs6IN4Vd0b1WTRQlQTFB2WAjZpkwWNMIS2yrf+o787
jS1iKdOv+Doc98dJ8ABfnrMzLqc0QAwQpD2uNFYUyx8dGSVxWKKzGfxiU2X0r5SBtBbOFX+ccQJh
Ss0zGAo7moGS3EoKP745nywg2yHbH6mb2pr30d/nKSlYiEAplptnUmVAKWxAwA9Zo2s8MeV6yc3z
hAISdd/iC2kUhRNnjvwU0etTXb08KiGH+1yLENkqFF/1NgdIDV/XqNvo35lrALJrZIFkepTC/9wD
aJCs6yo4ZAZ3RMZCCho1LEDA3DHGZKzatdUnHvseIyfk25IUHFoo8Txj6ANvi/kHQuHKbYegxCLE
rh6RbUYzEdFVBwe/8HDN2FcPAHH03RWPR2MsXqs9xPMKlL0bvLpUP3lfA4bTQqUBgOH0pO6vYUSL
LCli1YJLaI3kkWzziWSMSNEHBqrFva/ZwWPZqhzXy4XSWYjBj1AH1SD5ru53sADXZlcGZbBel+kS
dZRB3CFimIMh52FWwNYW6nHkS3ZyCLpJ1pD/BKy+YvtXhBs6BRWkvuIEUHKQqZaA4dOZkmpPBvim
7vRkGjxvd7vJ9vdPZ155N9b3rKbuwWJj6PJ4ELLb4Xl9Rm+U1QFSQgZ13XvR+o/Py2aQLXfNKnHO
TZSn+KbBZMYdVb8FFal0VkxwyvrKu/IESFxI7J2ndTPA8abUkVKhMObnaTu7R5iHCKKRiaJlQE5v
TnXuoLObiDnGrJegqHprLmNqFc2jdkGTIf/qc8fGQMv/PN9fL3gnZfLngTouNl/Br9goaTL6VLO/
b971smIDAf6Alf3fla67raOvuZDU2rn8t5xpO+gEnKeZDeFhwwdoK6K58Di2m/3rdTGZkeBST9GH
BqNVtdBAoapQaBk62PmiMygyTqmZOy8xIcQOWmXGjEpQZO/v8jpSRK7KDMuKeT17ndR4rF/tQDpV
2Si/92a3zE9v02BcsWHtpq54AUTlMVS2zoBkSk6hUCvEAmUW/0a85yhAIThyv7rZroh4ZhRtPpZH
crhrIn+DfiGDS1YznwDLA2kEESoXviukCpkLQxE+6xAAPyI9NuB6wk9VJByye3vvDhbcX2oCqUMU
xg2mfRk5+EHURTakTwC3z6QnVhosKZcFQkahXOezJSHDMpuZQu5Uddl5WGiUPfSZBnOAH4LKlYGB
Hrn3Ylsrd/dWBL7Bwexml94WkjcQqRLD4a0zv0czW1aq9Lwy3fuj59JLT+ecn1IE5dmQB1NlwCG8
lLGzHsStodObiZfppjtUQhL4QqkHz5AvBJNGgbYlfg1k6C/FRk1QQavyDqz4MmnpHk97SzUA5xL/
AJ+VCf0FGV3Oz+PaJbMusrzNLsMoPzadinpr9xWn29jY3fAO1iLSJF6lE6zK0TchrRVdIhmA9d+F
SsmYzWurmQhuNUsCwbtOLJYKvkiVZp2/HyC3V6Iglsnbep0ZlAdGCuaNP3CLuhVNGE31rz6AOB1n
ZJNbR6qmpC2islC9CQv3n192SLrqUYjBVUZ+a+hSuMHsY3VbGED5vX/wLRGfgLRNU6KCF8scxXFO
hZrfSYWv6YeinImLL6QE/t6NTWAvZvBSmQg+eUJ/jBc7GGKYXLh3KQJ6SfJ1SIj2rhqTjZcZi6s2
yXjz+2+jjcASjJZB6a0I7r9OuYVJPAGC/lXzGDxaiINck9f+FcVwq9sRmQ0aJDbbG+Tl6DN5DKrI
9wiyoojEUYQPV68IJI6185FKLW13uQraab0qTm7wMnqCxVZYnsLQ0b7tDb8n1et+RuI5kRE0cLom
sv+MJegJon2I79J7wC8u1pt2yDdL5+ukQS/bwj5pASn/mrFA28t6cZG7C71Zyp+L0RHTQQcawpO9
RlX7Z91yoHRpqAAtz4lyroIQqh1kxjSTfaYHaWFrV+slFSEYBvV8mJEF2QP/zW4rH5YuLN6orh0Y
T7zcpjroZ4u2DIUklRoti6dHpfzjkBJ+DIU7jEnwj4ticUwQVp2mevLp+iQ/QWqXv6i5zNmQdivY
IIFp/GozfktJfZWMXJLSDXcTO08JKN7ROhb5oEFmKYhgMkJyRHq53N8+OMrJO/pFVC/YVtODGbry
eiE/y9AZYSTpy+s4yE7LIpEmLTmV3vh6iR3c6rvFOhjdXxy+mM4nSP0aUr/4VnGPKkq0mw06MQXE
+wp4J0l7jciyI0qTISj3dCsiQkXGhuNA8po48Znd/Ms7w94+DfovOGpRjHiojZgnTvRVBLjMbLOl
0vJgZL4zjD8JLoQS9+9rv+zcoxrexP8H3bbvKbLXxBUvyGykQPEg40vh7Qd/ozH9EAITaTVtwp+F
U3D6WAOrU8XPvUIQFJ/2pYSk0yfHpAV1wkrbixAke49uj98VUGFgWP/vcTM46jmez4WyrrUFMgX+
XJUCk+05IMM6etCQVXVuJosiYK3utEYNSqPHbbH385v3hxTsnLWKsz+1WI7jubY2Qo2iQo8+jOJK
DVuL1Ex/WXKXh9WZp2UUivyahQ5VjSiJ5YBE9WUb+NF2oq7IhTHXCDWJ2b6RmEvJgWrQAFJanC49
dm3E3yymbpBLZheF79bGFgSS26D8Zqxj/PIaHdi3BmVMNPjJqkSWZy3zt3HhZtbC6b94fru0J80f
Oj1p9eF6XtPJQGwLx6RmFMEH0xEQjMVmqP/u6OvgfU2Ah0whvwqf9rYbdmMEsO6QHQgBLFCV9QuK
xWdspIXlcGTkeE9JG56MwqyAHnb+iVEjaLlI5OyurHuUOSydm146d6gIm7xuZ790Map38KT0XZqw
FgteErZcfgCIkBRgJxi8jXtoTsSVI6MhAVynOjBf7qj2t1C2JBSGKsL9mvh/jcV1mhOwVIogjwgl
GFMLWPDx5nb3xGILL6tyVHl+1lbXnmnjkPrpkg6s2w028IqPNmQG+el2uASenMDAdivAdapOsXuV
3MhjmohUUV8As481rI0OQjo/vIKcyN5TEyvkIV5/8eWqrMFTZC+1B+kg4So77VUb+fnCSqzse67w
ZSHnq9FZRZW4SoTwzYGBFKeXgc1wk5jRGS/uMOVRm1YBzLLuJu03jQmLbJb/kLHOBSVxH8AnN6n3
OVPni83HgnoLKm+23B9qb6JjDeHzJQIWo6QcnhurefOcMy3vOU8TGADIEAKs9txHUVZsTBKEDbuN
tgNE+ourvIdOiryrLeMNP0qoqyRD80WJYZs6zXPCsTPS4OuY36H1lM8VJrgg46tjRE9jDtiSKpwR
hIOfulxXSsP1Yvq6WIRaZ1qHURYANLxYTj7hPATj2NGSp+owvVS/vKwYzIyfAjqzV3tFDMQ/mqUm
v2RsXpAuMBuY4Lqs0KaCobH05EwN0TrZMzdW5BL5Q3yQBeLdjeQbUhBXIZ/PxdSPHQikJDwFna1r
D8d80D28w1JB/U7Y2uGFXQ5ABqELYVJapshTtk5FXw+f/+FHfcMlo827Fakbhoegc/KexanJDcZu
84e2hgKw/nFXfxOJlO8ZHf0J/xWSrMo4fcr5oFMkp1Ox1SqQ0M4cpjsjTB2ZQq5g+aJnQsWOnyA2
IOvdtZ9soAgWyqOUbHFdxS/HZ9rIe71v21Z6PsvUAOdIF9OmkmO2tOA32nf7emYnaP13etGZuN5l
xSlWdwKt1U2h5dweBI9vAS4jbHftuGb/PJtdXgQCt3Mtb3RW+FZG1w2bKIksJHzaqYj6aUjqihJz
7JkPEGo6iGoADNfKpM9RIwcZx8ZjemdA3HvnZ6Mi/djlHkRI2R0p5Kk9vdslQcHgsCglBaCovXjd
JlIR7ekmTpzKqaCmLZ8qwdC4TuL4rLBBbUyb9m6affdHNh1SOtGy3fSUEh+B0ZMbyw1orwX96xWM
r9pQw6z74jJDGSCMzEpnoXhh70BLtvd3I30hlfJcpzMfaB98fIA3U+tqfLuQmMRj+TVyNQreSHT/
8NwVokoK92hS6WgLTxT2VzXqbK3HgAeJtCmrp0/klIDG69UB8GBefGZn6MXerT4H5vpv7C3rWKRu
9+1k9bXC2aEg4/bdIAyTWz6ITiv8yWTS0qkSCGsty7u7YzFOjT/6d2FtIWrHKTQgjUjiqbkbddnY
dKdmmXmTy/vM+GWV9LXBFiaqGadaIPkSae86bqSPazkW6qx+JE+FKhwg44VdFW2pG7Ch4vo3TC4j
qyVT0tcWsDYtl6CoA7u4N++FLz2uO6r5SKPjIX3rcD66PGoQrJHi0b3aFsPE890jtccINfQdRabA
J2QVF3aKDvuLPAeMy+1cnl57xIjOZGy7G3FelaviRan89Dac7LN1p8SNsIMGrO1l4+AHIfDnlqYm
NQ/iL00Y5Ig6cDaL7aZeZP0ud5iHQIW2ytS3Hn55fNUtPEreZT33hZYDzOZShjJt+ml+jtay8EB3
W6J/GTgQK63TFvVFoiA9QoKSfbVXvqkaIDBoDsom7nS/7B6CEI2lWE3wHlesa1wXO7plT2ipFBMx
dhNSbKLw+AG41GaZvI0jpycpTEubGZNYzN/gmvPxNwzfZjvs77yve1/zzDAf3rrFiBmLXIVqg/kW
m63xCFFzUgt6Jbrp44dTecJOR5KVwDr0luATh/pEpVVHCE3gnBNpmBw2tDd5CiFMwB3bamxLFMyu
GuA3FRuklqlIAPBUlQaRgPBfyUy05v1igTGw/09BPIFov1M00ZlS5nH5mUn0E7wTQdFDn07C1bQy
II53gHqHLWarmosOLhIfrCvL/AkWDffUqAqf1ZsMjCOE/fjLCaKjVvTMqgXXn/jkpRBULWIfxDzU
WKSI7aKC1NMjtNwf3dTq931b2TZvOasXfPa2Q5rGBci6XwbC2/TmtM3iWcw3D66MC3BOROgvr2i6
CfMkw/+eGuijbZMk/1PLaOneZIQnqCPoewJw2WSc48z1OPPcpprZfSmz1x/vo0GLp44fJ/bUPoMm
aNZhRGSN4IJV0uzoJJ1R81ZY32J2C+AWCrabmE0qWbsxyWYzINhD5VkWgtBZ1cjMW9YRwgbkf+oA
x1NhZL25NrL1t7PB54nixjDaDcS7M0wzTX+LtPSgHOob4d8Bt1E6fxJM5UcLasl0k0rWvfHzttSh
3jdExPOjF8EdTy5XxWXKtbU/Q++EMjuIx0MDfxATiZ3ohsZCJ3C92F57CQEzl5WXhuQKOvYyaJVw
Kf+/ehtaM1Tq1BOJF301wpeT+HRlCVDRFelV4Fgk7Y+pFy4MSIgti+ugf2+s1KXjzFgOftu2c5Dz
Xjx1VEZsFbKD4rqW3aDlK4sA3aZUva5zsHL1yxSyNOjG3dgGenuZiY8lF1Rp2m3FcCNgL1mVmTZ4
tzxHwtLgORicYx7tVbEUgmUfT3dHaP2ZpPVZ8qqtLlRhE/Cc1j49ZaW+toCRMnmACMGk7muuhU3Z
DOShhfhes5K2u5JFktuXrWQ9MvdSuewvPn9VhGe+QG3bgrCOSH7llyPtlRVpnkmVh4alDEs9UHF5
V27nAbW41FtujCcy34pBRMs0OjS49nQaTj1AXCl0x9O56MyVrZfvZmwIWEAZFr8LzrE8Hogt3MN5
JOs/C/UV4ELQEp2ly84EU9w8WAowBMS7DcXPIupa7BGndIxVMCQ0kiz5zZr1jfyeVVvXpR2phQBq
XlmK61AgvzoGig+7xfv6VOYzYgA2oeMZqUYC8ftCcZ8ckSI4qIdeqQIgDJkmiJjXy+kXbqJB5hI9
EjbmItJxi4lzZqEGKHl7aVujctlcWRbvIN2wTQHA1aqdcQXoZ27oimbZ3eAKByd/EB9EvQFO8iuR
d2oDtMeOQ8w4w1oIqG6WoJ8VI3rnIfoiVxqz+9EyTv60Cf9pVEvZh04nNAjYTnpnb8jDGOge8eSQ
RNpcUUaP+Az6494E5/ZXpduAzFIIOBfy01122Swx3BZyRGS0Mhn8z/cXPrMB6BWAYOlQ+J8lBYb1
7crt9+Kr85QGjw+hIJBGfxx0+uRGWmi/WhhHE6cd3Sq50H5XPkKMu5ZiwnuHYWGQkgV7VF+CVKt6
issGQxfSSZGnRvvwUw/1b4PvL1AyVOHHFh+fKSQuySiqgkDyCiW01ezN9OocXo81N4qrpq4rWFnc
NejbVeleEA1Ysm/fI8NK8nC0qOSu99UW+NwkRxKmwSGYrDut9kiOyr3WYfk283w0W+2nP9H7oKqQ
LrjMUzGHFY/DnsxaMS5EWNm6zW6J4U/ka9ATqQuEQ88DFiLolEgzyzdpBHqbMhNHlJMHxRbnsJwW
zta+tUsXIUSu8rUN3fDZ9jz9u2wzWfRQxJutxGCoih6Ys+Dl6HJNuBN18nQLQGsPZV3OAAK4E7Iq
QXSkGZrdVS5d/3rylvFYO0WB4UILgnKNVeZwGkEHXMy1GhMIM6CoDXRiaf8t4Qnb9EI1bRYOzFnN
guTcm0d/szN/JB3z2pbQ09fYoxZqrJlMvk8633J6Ya/Hr21ejM257+ObCEKQ0mccWtDsN3phgcK+
WNHiW7PGjf9vaxq4XAUB4MM4Z6oEW9PFZI992v+KlE4NvzU6N4eMrfE/zY/DqOL2HuPAA2eBzG85
nrWdvkrezCJRY8FK4Dz3o9QmuWd/RTW/YkiLdRq5yI2crCNV0+C/apX+fi3XYBeTsiq5QYqdrTeu
SLVkmtJhL46xyTm11PkLOH7DAMkTJ5ilnnz0w0rAhLFiiuraZDZpqHMQu0jB6tzj+RF2xlXCzJAw
f/8cOJXscvjazrnDyjfvvjk/zZTXJcGeZw+HIJZr6ytWdP0fuZxFA4kIqje2mAccBxEuRLh9BKCL
ViYUIwA4Xo/o81Cp3x47D/wj/KsE9gPM0c0uPWr5P7lOB//AitN1DOqBT4404nEpkmxYCd3BBLee
PGog996zQp9AKqMlhyatalXNZzKqL/iyvHd0VUZkH2mAcl+tnQrqzoZrkBUVuCR8PPz8tPudPdfY
H/uSYPiILZuBEtxHInlC0hh2pC52yV1tRrM7dc02vSijhTFFfSTQW8t8nr7OsAaCTKL0h18+qv48
FYyYB3/29pqEcvuF2LuGomlD+MnyAp1/HRbLoZNbftsNUrpBemdJ4UNKvoZhaHQ0MBY3ZXYpvvBA
TRw8k2ykSLlM9887VPj9lyhNRg1dW3bhK3Mtt+an4v8ZFGVMVxDmZ2A/II9sIP8CmeI+/dhlHwGn
VG94YYSJxKLwpPXlL5dI3Ans0k960MU5kr74jFU8nDN0kX7vObTveLNxmUsga9K29s1iEqulr8Xp
Sdt8YhIyPYpNSaPaLOQfJoKVOqiMkLgPcEVhNdwAc04Q+2nNaBJtcVqz1EI0gw4pxwcupXgzT3v1
uoNhnuordETbYd9XOoeBjefopQzRwyEicLaNJpdd7TiJfnfJ1/Q8QEr2AkRdRuBP/UcF8X6lsWBK
c8qILPrPA2Vi8KjcD7V9Cbf+BvLtnUEu73vB2ssogkW6jbTvds0VifJUv7XAeKB/jREBZXDfzNq0
Qo8aszhPGmjvA+7s+Cm2wqggtPkRGtMKlqievc/sYhnGgsyPWwY0xw/DqG+PSB5FtBc/IswLrFXG
mZXhR8UGYVjcpLSGGmSDn11f3xM3374Xnp/rr4j56C6suRG2zdx/cKsjxXbI4pRHxL0AeydG1y5c
YXKJ7/4JhUC12baok7XeN6QMkRwloxgdMZvyr8l7gl7ysS/NMH/LyZ/XUn4X7A+G0tyUlir+omQ/
/mOKbhj4sFFkNQlVBzUTlqOKft+JiLO4fwC45uK3KP2TSQnCLBGdi+Wk7nVD6zBEPbP6lU/RUDbZ
9qwZhpLGArgteCy9F76HONDKfrSOFaPlkHkmyg3qNddyBD2BugJf/ys8jnGhYXCV0z2SnBAATzni
i+zHkoImTjtXixktt0wtO7HQuShP2YbvVPqy5CNejqf3zzlpkrsOJklllfgFHluKsv7dG+qWSXXs
Ye/mO0q6g6FUE1yilZiek7ShSXywbhHvbqQq9j0Qc4w5/E8HtDU90ziYwKcKyt09L4N59KB7Gvz0
uKjD7uLuf1aJOEgjogGljfzlvcLnEPWs+mpSCw0yJAdGomx3iOb/kTQ3f6E9YgO7Yj3zI1r8gol1
p3jyx+dDnhEc07kNZLTjOWNeKacaurBawJZHcnvOit5vyl86rzo+AratpM+j8kT4DQ4g0fSg1yyl
pDzq5eHt71WcN7DRIh6Y+ZzJlOuFL9xNDNSQf8tf2NNoEdI3qfwYPsfdEIaBl3/i6RNAjAMNkNmh
AKBVGdly+ZBUPRbz2q0GwYNvEny2DFtrCs+T+NvZRDAgpkRn10Rwl7EUPKwgK6kJAYkE47cXzp/u
NfStd+IH3fofjVfEwrVb6+x2uqumPzc0V/NCNUIT+Tc8GNMp5kA9nnGCA8f1Usm/vqZ2bHvVxl5Q
xZWmW9413tLQ/fsSgVJovbOvQrXv86a6EGooaiNSaToNqA+tPM3BU5+HJbkgv/oKw9fKe8zaKDtS
KTydMvsjeYf9JM+cVIXbl/zsaj2a2ae89G0IqeCTbvPuk905MNEgy6kr245Incnb3TRqnGiOUG7H
Qgd9Y3vBJInjS5TQxqo8BmVomvL6DnFZ6GWgEf/XlTUkIwSeOrU8zQ245mMGiIF2DYBHeXc3YRvW
87PqmWhedpa9NUwSmgcgLrYdJlNVvX92xgbaoHPgWyOHMA0KUjzHvgDAr3e9QOtPtdcu1yPgcmbz
mfqkAN5UgsJJO5fHKMGLcvtQCMtbaSb+t/zKe3xRAxPePbpfgsMuwxWAUVGX7BoXC+3HQEXyKUCy
eWwbjrn2cVFTt+DhU+V5cK8/h3Lk5Ot052BhKON7CRRu03lXpPGNDzFVQaskpZc5d7S6KXHyOWf6
BLcXSLS/FPlXd6/lbHRQcMiyTa5mq3YZj0g8+R0efAueF+DEpTHviDFh/U7HA6tXfblrtRZ/WHiN
hC1g2oRXUrd9sYBJegsa9hoDvG8GKv/2NCUEpfKkLoWPhusdbyVdMg/X3a3JhmgnTVx+l27wGrOC
zhpjd5LZRb4GJHG24BHo5JbXpEjJDlp3WtqBNkfGZ/SHpEDZUn+xHPeU9BlBz38LqWCqU1j/RNAc
WDKI5UNKMc5j63Aeczsuak2aspV18dr7FthgucfFC1VXIBxe4yaGDAW1AOfnpV5Q9fGpHWspi49U
bZMtLY6OLV3j2vCojQGbYMmBgLo3G3BY+czhPMslWL62x4T7rSv+BhiQvBuKE8MY3tomtRt3c4rN
FmmytxbmOSwCHEa3S0EzZr7eD2gH9ln3X4Q5j1HiOzmX3SnHIzZwUnJeFsV4FKz71VtFAPCrdHzs
aGGKVbJbVrP4vRZ5MNTSResHPo62pSYzJIYkFWQ17wHjqNT4TZBvivudAc0xMSQl7SeztBwy/RBU
B1qGA44KHhVhjI2O3GYUuRLsLYa1SZ19HS77mFD4HiuC9rl0xuJ8CferiJt+Z0krOhCoATiAs7yB
kNYusmH9nyDYCQ17N0Q5g9q2bxpi/eyLjELOqeUHzZ/6yOVnISbInE5j34Y+vBpY9qzMtlg+0WzV
2Fk5jRwAeOeWoom00fPWrMvZrxplsG6K8phrLzP+wuK3gkOCBn9Rdvix3a5W08w57loO7O20zdK6
ckbKBx5Cf6VcrdkG3pfhyqG7TV7Nil9TvHnXKcOsthccfGsuTRdNxVQ+QgyG/p73BNEURMrw5Dun
jJkECHrGttibR6J44PN/U3wzeTqjWSod/aknocxEsHA941Mhf34VwwwYYvDFh+z9g6IgPQ3iyNjZ
ZD5IFEf98zdaZErzBZ5fX9Xk2Y0pLeaIRdwXJxgvoZeY7ToU8vyiYOiknLTUBvM+fnPnX7JUcSqi
7KBSewu5jlgGavciUQvnZvqVP2yCy2MZOlzavdM/XSAKLHXiqMirLgtSAJLAESFwrKNRKUdlUaST
Lwo0h6ll/YLJ5x5Jjxx7I1t4FLA5l0jtirYK+eb3+SyRJ0zxniAWM9nGG0f9Mn8Uew0aI7Sh+kvq
xbhrx3VsFOsnby3Tgq2LI78tShyA0fYW9A+RDuR/24vpLZeMXsCnizq2khgT1RuGIz6yB2zG+iVZ
GwYONGvr9WuPB51RgQSgC5iJSz7l+JtAIXqeBrPPiqi3YfQ7V45DB2ymgj/MjQVjKUTc0YuJw4G1
Brz3iO96YSmh3+qPYU74AJbwjJxECNqWr1Chz5zw89ONUvJABQ49GnJXZPxtrZEXL4T5z2z4Au/U
NUp/PJ2zgb0vCj8Spn6MdwzcnvepZOYR15D2cGwt9Lx1V7w8zVC2jywUcxIN10ez0i9Ah0gw5F9o
dOqlfDV5efMKyVOK7TzvlSXOKbkyDrs1YlQK51U1ldYnCyM75mWzEzqYemVs87HD5f3o1sjOsOHR
eA1K8BcgFljImeZmArvsje8gaongngmagemGEuHucnuUi11rEkeFmt6CEQAcZB3kASWfv4ADIFqQ
5eSB5NLNRCrD06aTseYIO+2HrrW7U2gnSwWBKvN/SdNf7TolKwKg7UQaP9dbBLkVqpEM4Q9DmxEW
hQ0pmcSff86AjpVxFpZ1U40j1HrvzFxTq7/j8SFfBk/0M/K8OXCcWqscZ/s60wc6Rjp1Z2X7Stnx
5645sRz/KTSGqoP/jeIZLmsek4wvMNIMjyxhycjpssq0PSg2Y9ByN9Zz5Grsu8bEs1ehlVP6GEbF
GIlh1iQgavwlh0p1ZM0dMV4Jdy55d4R/XmIvvn7qtg+cdkkLM5M+n5zkhanExXuFS2Qxesl33C8r
3gBNzW2fo7GzDhOoETBS3j4Nk2V0uBzCZG7GIDp0EwXFETMjn4LoqAtq8q2RdNBI81s0H7bSL8aj
l1FHjFFJ8E5VtigTeGvfHmsBrHF9BNREcZaidrJ10S/lIOK2CPOGTke1JHL1D6INgKh7Cgg8jjgZ
c/LG6Vjv9XMsPV5Zqadb0zMn0tkZU7fQ9VuhVNwjBtXx353ZqzDXE3wbmzZosmKfG+0c54n1Gbd8
mqiXEfAd+MY0aDPFz485Gj2lPA7/zNuSqUSpz5jyd4Ac62miqYQxtmyAkUoEN2zDt44ZLHt6hO9S
r70NkL/bcbF8iw6KRTbnEJksUasML3YGqNjVEphcl/Cu+Zd4+LhzDZblss1qe0LYxguvZLdtIJii
6qTLVCQa3zRtkcq/1jtXoxl6xvPyg5bchDJiWK/cGPi5abM4te6+qGWoZZtayepsSfTyj2Ujifp0
a7cMrQLPMnZNKa1n3EyEw5xkhDmvopokLmE/ugUOpCbPpxV6Je6HXRKe/1ITcNcPaZeDM3C9kvds
MShgDg3unBdhMk6PdQn3GYX7H0rg8W3+uEVAz9QtlMfkJkVRcWuLX+SOm8MM43wHAlvVL7SBgnkG
iwJr8mSkRgJMSElzGE/kTaSzD4hCNrjx1IbtRKtWsupjtUzqzIcQIBGRmcemgn2vEAeVBasRXDNU
W+XzcVPSh18X7cW1PbuP/MdONvsdZ9H3GFsvr8sEVXhDgeAR4UB7oue1CsbMBLE5CjcMt0tv/29u
2wwQGJcYWw+6fu71TTgwyKEtHXRUezxWot6M64pmDHGQDfd50zBmWH4MQM1NDAFLXykpotBfps+5
yE4724up4ZKNfIBmSNRKihTnCvvltUYfsYxQvda2z+VEktq8ZsVKYL+ufP1IemyFFjmqRprQoVDY
HB1D74mXmZ6kepTNTq65iT8tID2ek6Czbippe5itxIqgAaP9mCLYHzaAAkYlaeQH9+CXdI9+UAnJ
v5rvfOB+q7jue/uNr4a9NS30dRiWvBHihdhlTN4TcUlOIkRKr5HyBzZBBo6A8EpRX0hdOrmf+wXX
HIcWYPFQmBhysFDJszm1bF1hoTucakNS5owEdr67ngXise7ZqCT2PzVFdESp5IbWgK7h8aQ/sOvh
yCAM+4oJH+xOeFLXOjzUCVmzA6iYfkdl51/zesSQtTLPiGO40gpHASm0VF73gDSl5S8nAenKJ3kR
oVcW3dbSZpNx0Ob4NI14we2lFnzJI325X2YgAqqoDY5salhglRt79wLFucYxyxdSuQIu39S0Hl5p
crT3byUsHwzxXBpzLKDyvX67uwVlcYMM4+JuuuoUV6vccaNULKmTq8feNmCthkJvyV3YNi24ERzc
HrTYnR0tuZxMQwLWxQ4unkfQ+jUtbpMgTPXJw/gudC3BPAdiRZMCewERgNsIzeL2m9bq/3BrSbq3
L7MDBAL+GU0f0cjitWNUZQWDs4i1VJaS4/d15pfjNheDm0CxgRRBCnrm6CC5G8dt/PPUW7lY6fq5
tGFd4RRDMwv1IgyUssJSCPibT/G71WabUx2s1RHZMD2oennXEKd7Tzi6qrjjf/gnGyBivi1qGREE
fKzuC/Jt85n09o8aqaA9KBN5a9mj48IG4BOwKWeqA31Zjc7vBYJOHDL7uwa5yslbdRzh6EPkcK7T
YcxFimstrSyxOyye3tp6Fpgbs0qDDYv7va8XsHeeqXo5SjsNE8+41KFIXrvsKWiFyJRaw6UFSq1f
zMxLN5v9hMqqvJOAYrhdIuJzHAnA3kG+uHSCHsLS6P+PqAlZl30O7pPShzw43huHpAO4VTMSJvzY
zFnOsAsrsPobRGglW6m2HExUvp8i/xvjTXJ6biM+z/CNqfenF8CvL+CEwnGjf8R8rra/l7YZX1Uc
KYOKRwER6v+ZjWxAExW+Z4FL2yMHfMUIai3dDEw0Dg/T4zH+m6vlDAWckY7SP93puraZyAsu5Ovr
X67WZtowGT5R5is/9pvSXdhYgTB7tbUWMHM2OjqpYgR5kzeo0qqMuPQNbq5Cbw5qy4PNhe++cF0w
M8MdX81jz5aKluR2Cbaz+5MtFiNqoL7JCjdaSWhTPXVM6qUSeGX5sxB7FoukaXEs1VPE7Ht4lJ99
2+eKb6rzY+49GFfvLqS09BB3vYcRSrZ14JIg6KFGaPSitr2BpQMpjY864f7A/GqO7h93wl8gNPvZ
pBdjpyLx+u/8OmFmZeK7E07Xdvky4GhRHyGX5StK4pwb6jkTo01cQiCVVK5ULLiMeOnFHT6v7bcY
p1EYToQRj/1N8CQ188BP9Zb07l3pL1TM9VvOYasUh4h5TC/ymy5shnYYHUOaYtWubMvk0JaliKtO
iVAr/uar64iYA7KhucyV+T2PauNam9oGlKseFjx/jmWOfjgR/xrzbCVda9bExBmCGImdFF84wuGX
MEBDj9JcPdSUv8Wcw2Kh2p3JbgI+SxyHiSI0g2XnM/17GoBCCNtr6jJYq/klKhk+tSd92NQ/IckF
I9+Pb+Gwtd9UwrCuvpy5IWWCEJOwcMmU8j7UTqKQhdwbNTM+7FvsZkcSD1z35iKJ2r4aIyPwzQ+M
s0DjiswIobdtUO+RVc7FWtrjtuRl7P2UxfDmEAldsIAshdeYSxOzJwC0+3fM+JzIGJ7/74z87Chy
LpKzWU3mWGLBi4ZKWNDKtD9CZMd50S4AqEan/7cmj9xkdMM0EKaJdvdQHFuI9OoalHqG83EQ2iJx
ieNWNCqJx02PSkgh8MaAvhlNNZ3iuxq+jSkfR4h7cOmPOWemI7ePygFuoin1+eKn9Hb9YZS6GJiC
kpxxbn7wViT7qlne/vJWc3dwc6xP76WVF3XWRl7KgD2Tvf8wfLMBgQyb8yE+QiyHTuVUWYin9ATF
hz0256vSKGTJbGJIAFnvpYEct3kIa0yOpgcFq8HbST0JEYFa0aolldjv2qeJvynUVXJDXU+uj5Ow
C2axSazMUiMRJ1wo+3rlpjLhnc9arI+F0duAYbsnrC2KPa1pvdIJc7BbAM/tlsIMkt+Qm8T/K51U
8wP3p/6eVxBEDpAo4kwpx72W+0M1z+7QIsvK7e8czpo9cmzmXBldDAsuPTqqDVsvwfGF1DfPit/R
JATSJIj/gUJ+slW86vNBgwpljNmpPrxcPAONdq+ID5mASw+mFj5tyf6Wdmz3kyA91C3TPnAqPmXJ
L1FLYStmLV07UvRjS5DFkRBo1ZMKN3bfuKXUaKQQBq3uc0wKP5cYxRtjnaOsdNEvMhGxCuyccxGZ
sWVKHMG8w66kmGRuInYyyhFmnj/7+HHQdUz4/1Fg1anWE/rKkWQ/CzwLKzHNVMeHxvPFt1/1KVXN
StjSm9+TNhQoet3cRPxgmkbjLsx94c4MTa97XsGPaa+K5QxUOLX7UG/YCZXj9c6YQH/B002NORjB
pv8/IGT/E/7EBGSHgD92OG6jhl5xItvbK6Z5pNTQJ2Cc3NnaHgE5tYdXCA+XFgdLZsUnN8e/hL4o
bptiIcwG1ArY6sc3aLyYu49VZwTwoNcX3nv18KE1r15Plxe8Pl2JoAK+GQvM0VfR5U8GhA92Ys9T
B4T20nALgsLTvevfp8QVYaKOuJfRTgycOhuz4i03OCCEvzA7kIrcXSpywhndyfRG/ZyV6VQs8cdv
tsfKsFbfkx2Ryp0AzL+7QNfT1mjVYcMfvxgE7h0B4HyhadDHypspwmuqVqFpHxeLcYEeWvLMu+2d
VFq0n3W11zMsiaS59b6Eg75qhI0haRH6weXawY9PvRJVA7Mha5T7RFEEiOpl5rFumJenA3i6hDUn
lKmJtSysH9Opd44wTWGIDF5mAwviAugnOF6xht1IC8/13u0x2KnAR90wCzILAEBLmFrFYmUMwWoX
cM1gc2q8/ov/zBzvQQ0H6M5TZnjk/SIKidqvjrH5hK+1jvkxvPjlYgYGOJaG2AwFbFvH/UV3H8js
YLMRAWRDkiDHHCbwvoGmrkbK9qMZyb0nL3z218TE6kCLNP1RLnl6CmYSwcCv1YsnSKIEiehoO2qp
XyCufi+aohyaK3TXp39aNbzIFbBzvrrrgTVMTlHKE109mTSlZs2E6AmWmj81gzkSYk5QcU/2IWTQ
FS2FvkkRnSSvozki3+X7j/SSZ43jrdwyG4oX5DZsuZvqS36Fq1BWy/Nkbc3TOqn2WfksN02FBRPV
RHOHQtsO42pgGVGNsVty1dzMsyRJfsWcG5HvLhZlZWXqf+buIq/6W0mOHbzflVu3fzq4/Weflu5A
soKdmtutxZgV4qdM5BgjulSlgrKyki/5ze1WD0F6/1o0tYGIbn1VzKk3RyhActb1wAXfhcR52/z6
07q40MgxOpN3edwUTk1qgo8AtOo297Ir2g2Jr2BjzN4dxEHbD/k9lTYCsnxlgU+pvjtqJIJgRI4a
l5cqYDHzS1svk8mad76ymqQp9aAoT3KY2ESet3nyyWZS8H/GTrMiP23O0KrK9D1sJAaVUNAGCt9d
cscl1eudofqnLiCbst3fTLCpVXg+5TsvPk3V/5GPBpeXknenYlXsz45X7PgUbLxQJ4CphfQX0R+K
iuT0RsZ0At89OBTwgjVj3P6ofQUSk1IGX2Fcx4rdAuR8qO3+dDfbVd7RgJrpFd287e18tHYRu69f
m2ccXJmxHF78kPCFJZOIBlOJsN3Hmt9FjUBCcc5B5uDcaIiu/DdfeHykg1DCBbl2UZpe0rf/Yqbr
YWg2dMx51KjPIO1EC/wlm1xLW/hfLDUX4wVEJMPOu485HX8usLKI3NXVObA13JSQ+U+e5wovGLmP
D5m9jPp7egXB7BmH1Ur1sh8bbnRgzBIhHdKOwgGyVNLfjxAOgTNOINDu8sQGGK1QeydwSr8iWcKt
PtZUjkmH/sYqVQNtG7G4igO12zJ3PZFiO6BfADHVjx+WUTBPiSpFfVMvw3ACDse/VlpTpF7HdIw0
QpTHEwqPseUo7hOO1rUWw9uSI09C4hm9ch/whd83I4pv/u0mTNku6eGlsD4PF1B9KTiQKqNOz4wZ
iAf+MUnY2gFmjmFy0f3bP2QBNQPb2eiTLLgNhcPKuiIusu4GJCa8TTBhYBeqBZKcU721KxlMFbJI
QtRIFd4HE/UJCXQBd3T7XtJFeKcVb8bId3EpliWsng25QJscW3vRZ53PVPo4M7QzEaVFgL9Ey6c0
bo8rrLSR2OR2av2jG9i/ZH5sRxZUfse4Sx/DP4Y61q1zW+ID0N+t3qlijP4bCKGh5aXMo3aR6U6b
n8gZ3PthdmhgrbXpXMYJ2+Okt6s0IQSHAR08ZnAxySon/4ReQKl5BZFIHXfu9oi8kqGPvjn2g0TC
475Id51QJsSGVPR5VnHijD1kbp0CfXDT162ULqR0yQ1CDUBKgEUrBoU4W/yDalgHo4GWN4SzxQhI
OfXUV5GvtWCta12F1D45kwdoyFLZKZ+7TXeWoVlhoqeEPVudSTP2/HVGzh/VJ6rJ6MWlZEvD7bpZ
eaLQvhyEOsAhBlZ4YhZeErGGwyyqtFcd/F+J1FXpPUL9981kdqaUVHK2SYOJcay26cuSmsHSK+W5
X+Ts/0xI1xUhmC5oDBMmV9I/HRCkf8xbqkdzDsR31cDtj0tD8Ba1T2lmYjvOCB9tOuSGreeXtrLa
y6k03Aulo17KU5VlebmxgeezPMbkEwAx/iuFzbLWigyjTd4JMC2QP5rHoegeQ3ZUiqv/q1QvNgzC
MHDj7IM/td7B9pEprR1GHAD3IAY6ahT1MHHDiyemiXGBDZ6uMo8iIzF3haw6d1Gkx0tGMpltLF9t
bQNdDHV9LS+l47wSAQ3qxKwhRUApajjOC5mc0hoJnxYVUdTewBvcxaoDLczsc7VlFglsBZS8zBnr
RESiaBfaMv6of9Wtf+cwsP07VwiVgdsOEqtGM/2cSxUt7Gw2G/1pqZYZPN2Sb5/W50auztLzH7z9
iKYosznVbGurvaWt2n3YcYjbEREcjtShZsSVsExzss3aFzhREKyAnZAlZB72B+IAY9qS7VEE5MwE
0nb39CA9Mxf0FbZKanWnEmt4Qs1ArC1YxzhHeL6IMAgko+LK6XGPsf2PsGx4SbSHisfmXA2ctUtR
keQ0yCHq8Ew7ySoQxmoYPJ+NARmdxAFIDQScJQ+F9+i3p0RpBpXZBlGPXzmUg2AOg57I7Jy/TFJE
D+saMS0i2pr2IbxDTdH52rQ5NKJWNYAPKWPlip32esfzb2/TmirNrk+UkIrmiPPL848am7HK8DO2
TBGdH9OOxlKd6loEWvAPOpCb7x6V+8kZJ2EPgRZrRZU0jcTDFBuKjYpVTdy5cvlHkA2QIrCJXdlT
5Kj9sem2oryj7gahThXV8J7WpxgW9mpqWy05ucQOXw6ZMFaJmjcJ5ORDKAAqD3PiJv5OGAvhsDUD
j2skp+SANwU0SMuwGli1EJAJqIocx9OrWKIn7h4/8sDQi8b2lS71ATLBhz1gEJAy08Fxo/L+uJl0
CcDTwtsui1fRU0T/zxitZPD55nacQK5o6NUSuexE2kh60we7N84XKbOChnrd7XbCmNKXmKchvExG
3dmic31DepixTdJ0tBHNdSFkm2MC74PN2xmdbCupIpGFtI4PrwK0fgN8/3WjJfc/6d9gbalPNT2t
tIqQtT8eg/7Gf2nWzIzTk46iKJpF9CBVyLe8SXqenbZJ5/W3JnpZ3aApr8QUJX1G05C6KEHVQVFe
xWXireT5FImKlqKGg66OZcBX1z1E5SkvHphGLPFFIoRU1uHkqeZoo24b7h5DXc+jfsvcO4y4BYdb
Wt+DC9nYQ/YSr69Ru+D4KSvmbC5pRYx5pZPTCFTvmtNmwUu/lK11VAIgcAoO4l+lzkSxGI5I9EyU
XFpUd794gc6K0T54/wX4V8kjm6CM8TtviQc/KnMjcAL+QjeaTs438jrhEJmQdVl5OksEAxWNT9r3
Fb252pHJy/ajB3K//USXrOgjSKs1e1drYWyjInYIeMJmPBbcttQPg3xLbvBmYMwkd4E3wHBqvuJ9
9ROn31w70xlTSwxr/bMdNtRWJC/uq8HD35Ttu4KidOw8V1Mr6tSq4/mECV/IgmSB7m2hWyZNI5It
gUzHybx7Y+EKxWE+VgJGUQTPIcFXBRCG2MYbf6Itp9NwwRAur9GiPHkihhrhjuDLohrt97KIiJOm
abqljU3SdD2jH0snKfdIlc5X06Bde0JFxrDs5IMWNPZl6QhNVhmG4Nrp6ZOqjGwsqLWo3reIBbT+
dyY4R+IeRph0R24TK/md8McoS5XY2LPSpSBHNye8WVrrEXp6VXy1ZCTkffHYa8p8y2rhzrbYJvnI
TuQETl1uvnwMmoWNKb8s/nfArnGXtkYc4cRmaRU0Z+0gp+zss2NZxSh9fSFcE13EJALG1AiEkIJf
roKUL1QzfJ1fM/E9Yn7g3Q2UXJ/DKCAiMkTGhA2MmDmORNWnVqCdsE8eIIDUYnqZ4I7X6nCTMW6/
+h+C92es3zkD+qf0UaeQ1uY9XiV3OHPcP7hJFE55RWCmhnbW/nwtcg6dNDHuvf9Wjsa+JrQw+CSm
fixgy9YXaL6+k8g4JDWmAG1qBTJov1Aihif6v4fhfe6sFADvklCrLw0W16h0AG92Qa876QW5eqKL
r7KAF2FRMzBOy70YMj5iZNKgBO36b3To1OaNYMhY7VxWyKY3kTQi+rcpjd+/ShvXmQwqKcLjGqQi
mDbqFed5CE6a04M/Wta8alA05caTfpW8Ksr3GIjkd2Fxl2g8UiSMBe0Qef6c/FV3rzQQ9h8vT+GO
GmuW7/O4AG4+3+T0IZfiMFoKFZJjq7kUEQFL9ev0a6wZooLV6Ol0g5JemAF0VsCDgRoBmRulg5ox
TEy3znz8BUHWXqX8JQHBwwksovEwJBcxW19mwelVENdEQVWSDV0lrPfScvIe3ASNb6B2gCi6LJcf
VCVSy7H8ztKHh3Z6pRTX4CgqRznHL2izkMKVbHctvflpp6wLaHVDHmpR3Y2My+aZrX9itaRWEAMf
c4y8W+7g1ZdkHMz2ndpCjmFdOVXUvFnvettvE4OT7ElXkyTrOHZyuFa1+XKLbLYXBtk0fzmb3cJq
VG0RbHruiPMpTsp3gPlJVcKT8+bSxOtiWWeXJJvROR+SBUed0k6s/I1+i6jly4H4X9AzwgLiGYRI
igg9j6ftUNio1RYkUR4f/P5gr/iZY/7MXrm7MG4Akv+WpGG3wREHf3DNdNnmdzSCGI1zpQtYlKqe
FgF8inhH4p4vfVh1N/uwaTyIVAxlD52bDJTvtaYXVCH5wTyL3h+v75W5UweGSI6jT+tUV2vHYx0y
z0QQ6htGxbM/ee4dVAyRYHzNchu2yfyof+re7QeCoyZhZItho9hr3YslxCQL7dagm/UjnqN2uYeN
qqiveZd1QiR4Y07m7YhVXx0Aoa/WlHGS3xOm+0hSBjfBtxUz5Is+mjDhj6HPAuiBJhqFjVMdNetW
YrBs3matnCa17pvJhWVT1ej+sQOqDAnGBRo8sgWH75Iheet4iSZdCPU0HV+A8fk2LDKREahsAm4m
QgbaRyiYYgawFyuaGChUDfNHYztWG9ktzRzGjcXsAvBmoi4jxsMlZFBjBSdU/IwvfDFlwJ8RjC9t
IN9p04GRXWF7TM/6/vxy6LJsb7NxtnNgG1DWyzutYdEV05VdTIuVpajY6/UTiT3PD0p7aQK/KsNP
HCn48n8d0wcosDzg5Zm9fnfW0Yk+/jIniBydnFoAR4D/wUwfiJI+YRtvWUGGF6RkemYfz7lH0Tc7
eTTjC74EiKmZiRTdQY4BT22pjKgavy5sen1wPW+8h0G/zQEKULNPL3lohd3UB9tFzuAAgE54L71r
jlm+gkdw+lYkhYO2zE3QeEphad5VZCu+jUSvLSDeFWFS/MacTaM2WtLQpj1C4tIjUDxrQbNSEPrZ
7mfehDB1IRDx7QMtwtuExJ+9M5JcTrjMxUsTHWYKrbwMRoSp1FVvUYHaw4TLUVGlXYk2EBsjZCwp
Z35VrWYSbFmQDCm5kfKPzEXx7PRT3YQvQJ2xDD/7KAt6OK5+hP9vTXDDYAouckRHSHU0spBuSO5A
6batJbI8Ky7Ts5oy5zvUmSGSQPrLXRq2UNZHrgG7npFIdjsYHwRY7vqjL3FHCWLy8KqA0TZiOXGk
tzS4vAh2fUeyHLdjtEZZa2R6UcCxWqGua92Cf8mwRUZqmLoDc70WMxZLVILAO3FAAF5IkXfsFBsX
9pVZI6PVCQV3OLtfaxhC9OgZwCfOVeB3fy4RTFLlduX23luN60AmDZGx7rN6mKE+B2i5Rq1OwshD
fHS5F5dI9PyugON9fwOC2hiN2xQJpLWTWhDz3bs81323jrGQRDrx7u7uG+2gYfWozMJQy/JHOP0M
eGFtRPyUFlLS+4tnvCbcfqm38NkVV02rH4A/4hExZ7+mmlDc+R+8EB4m1tBAHzz+RycS/ezHYQh2
EWderw6HyU5nZsj5gvsJdaOq+iGbJXQnSjLlZhdw+mcMpit45E0ejEftLldRMc3snOK7L9gbg1uL
uvUflzs4RR7hSNTzDCAzR7cFVMuSwDgQY3LtrE5+g68Fi0v3ejw5t2ToPqguYRZDYWsfmcwUmDPM
l0xOprWAQgoYmb6WH9IWHu+pRwkDcntBbIsoajnN+EDEy/34kl1AeLd7uyp+5GN1WKwgL+FwwvYi
y2qHOorlLgftcPK09QzWmEmnNkXVSKQYpcp6oO44nZdI8KgJIGkC0HmO7jWJkWnUjQqbHYHuJmFp
WlnNJHm+3qazt0Z/eAIrHKfA5kRuOFFQv8d+k22SF/dB7alSlT+4s47xKazWdOZO9ffEwhLFXE03
MWF+P8DNMX5qk6GXJZ8n7rDNp54x+SYi0ZmDp6lQAgNe0Jy5+NQ+hyjZt8dk12ZgGs4EIR9gvYgm
xHqrlRnPfDGC8C1aO/uXeK+a+TkGQD8COHIAE8OjA3OgOm0PslN4itADI356/YlhOq21+1RKTtn8
PHBpOmrs7LihtKBazyicJtOqPEIiIgSVX55IXr/2EB5H9aIG5HniNcVRLa0ZV3CJBb1Qg1jMaCsO
k7OwYsAA1B/XOCHA/u7T+hz4OeWQyW7CgvTx8//iu5I7bwH/cF8C60F3T87XU+LP5bc/Mf68j/2B
0ePHclb/d0+DJmhtrwMsX+lIg4WOQkmrUwEnx4Hs9o9aAsqHFNW/U7Wkay4MbamUUCBA+lv4D9Lg
OlJ15OEA8S+Me4NAPs54ysaNlG+Bn5OTGLvN0ITq2pY3l2IdTyWk3bCSNgi9ux1dGYbE385+DcRX
vxGw08Bv108MuEQEMgCU20GdFnIXw/wkmQAZqyV9kH2aCu5QejEpKA3cdIW6iVHGjE987yeNxFK+
8PbQ5jAPV4znzz5XbShOhGMCDxLbKRk8R/c/V2WtbX3KVhxcFW/nf+ZsyVsoc+G8HlE45PkwVxDN
xFdr5+P6ujBGzwHABS6sJp1qcoDRvfFD/ZEqRkBTSZqcbbPTA6CldR8NZX4dcTGtcBLYk+V5neFx
CiTMVTrH72uan9Yqd+Vg3Rr1GgM5a/aPqSv2MkumeiynuMZY6iAcIHOI/zxq1UWjyDsVicu6d7Jc
YXcnMAXCMmFk+YEFbL4B4WnPFMQmDLXmfOmuV9or6r6S3np+Dnzq2Q+Q/GtSxhZEdTElJ2jj/NXO
HpwiGeLFVVIcGC+roSX6JZ0dTZIJNnZbnYdowGhgk3Cmufe6W2u/4jfRF5ZjVpqbEPCYtZDDAoTv
5QGgwz6WbtyB0gPpDD5vSyBtXy2/ngvOl2Ar0Skte68AgXlIKu0Wo8dSeGce1X61T242tFPmQzTy
VDDa/aRwe6py8LQmtt4TzVCB4oYBOv0fue1c2C7cwIgyMyYrUWF/kgXRhC/hc3vBmrrBAMgplyuX
BE4MlGdMbvuB4jhnofA022caTOwUO0Mj+pXJVUzFPp9Ggnm0Ffx3If47sKXzRe5px0RoZpXQVhOI
cb5PeSbH3BoPVVwIyuqnzmnGc5Fkz2hXkN0FlfYpOygTEZn6qdo+dv4o8cjaJ41ciTB6xx5K0TbF
Y2r643EmagzttT0CPp/QBn9oF6zFDC9fr9i50o4LbvrEARixWaNiYQXPtvQBi+Xm3F0kkX/hERu4
Ol6y7UpCw9jefFoZL5hDt1PqaxFv5ZnHw9oZkdO9YyWZuS6x8FFFBFdtyZZVSmKEc6wek4/kISFN
eHi2j1gHvxh0zHkXt2o0xjdK+HmBKJJfabLU+nGJ8BSPJt5SW1mwe2dG8cJ9yQzvJTm355oV5fji
j/HtzxvBSNhNVaaeHT5InhP+FJ6Eo6AGdwyZteT4F39oNUXxPgPjFm1RBDfdyppYGSqIavX65Rwk
Ma0lYUY65gcnmBiQAaeaxHRASHmZf7M4JmiXBzKfXzMnJLOrERihzTdPbt7e4fYupK4iE/jRafE+
EGjDeYpGRilhjPsaT/N0MHNgQaOBEpq4d2l3geQ33Vg+odgIsysubWE04QqDLD7KaVC039G/V1aQ
EwqurIOF5m49dtC9NIyK73BZgbSHHQWr1dB7slPGOotak//JJDrNMnX1CHm886HMXmads0nCzPrp
qQQVdhRKF2G1YCyBLp7AaZ5/lcDLbmfiIvAWSThj3tixJyUAVpSRnpW4nW7p1ZCp0bSlHK3QyBCE
WN1hh+QuU+DicdlGFzwZSaF2em9NoTl7HxXsBApruPIyi8WqQ00dg/Bt0Grpp0O3J1ZIGxZ83bCW
UO7JAY4vYp5zDYBeIKofYXdEkqUV5YTPKjzMlzV7cdEQxfxwu5FxhrTdo2A5HDR6SapMCFL1e/A0
4YEnpxAFIsxNfbxXWBxa3GR5dTU4oxhl0NX7PVNA/smKY56fTVPN1oroVSdjiIACTqcz/7j18CP/
jIVJjcfSkFm0LFGNKvaJ8itCOWRmJJf8Q0TPI8cTCu4MsWlK8tPG9PvmKbf+W05BbkeUKljnfptY
WveltXQ0cIYnnKuLjbphDLJ2pVdYCrG7zqOPaeX6qK7S93tlFICyAXekc9S2/fqyvP6soYReaYRl
8+ORedU67zlzWRk1I+36feqmrsf36WebBr+WJGK5OPCLKJTi/DF6TYdYg/5Gwl8vVPInNeDG/t41
CdlQGA3n998i7giKAArkBgQ5/x3y9UMR4m6lkoZGEnifq4IRklnht4GRLcbiLb3XB6y3HbDarMCA
334FUzyf9T5bcpSnO6do51HrrMijHowGPc/iQ0b3vLq0y7Sfb7eSOCt1W705tV2cy6awZsMxOHL/
7IkoUa7kgIcLg5/7WiSiXX4z4dx2a6mBMxl41LLqQn8Rd0tRKWw2WI+siYLGKwT1/DBoBYctwSSl
MmuZ3h6ZF0ji1rhcfogRCODcqGecsc5aIy90t4NXObnvR/6yZ2inqGdIHBDNy8rBpZFzgFCOZxnd
xeQO9lynsb/b4R9wnUQtHF+tjkezU4pihcxPgCxnPhDz5o61G+mRTDgTBZXbtDQdmRghZrZginjY
in5xwFkqq8/zykDgzwyGn3iuW89wrEdZpRbbZ3ypHLsPNPiFs4stwx+1dyGKLf1NnGVTSi/PB8Ye
cwvVTmN370qvMNNBR2XrCv/xUjp8fJ0YwWK427XMSXKG/ihWCvdtw2Sl+DI9RDgnT1vHzlTLI8cc
JHyG8w5M0xQVY9hZKZsX8tUOjEsM16UXmzor9WPqxKIkiWTEtvMnBS+KK5X2PJGhZyTsgZaBKtF5
XKhJlFG+bPm+RJIixk57G1ozagQGwgRD29TxtyyofBU8SGHYI3OsilgdGyHf1y7tXN3r4LC3lNy3
mYtor9RclXtYQaPIDZxtdi4UhpxUzRQpx482AvwUFTnLrD3YOZLPWidYKSQfZTJ95Tf7Cb4pm/2A
AhG0AqKXnX4DHWose+SwdnviGGIJRwebN4kxkA3XrXaNffkWo0Z5rrtfi+J76gG/WwbcjJhAAXtp
b+tGlxdLNBXXOGReN37/PqD12nsKYFF5CGV99vh29JkrOwQ45qmdA5yI87lUFZ5PbLjbqI3iu7Wh
qzm4JdWd2PAf35hik52oOCMqJXCuS/jlufZEclvXps0s9WqPAy4K5T4wFBTqwpmHLsGCoCNubJ2o
8Zf7Grb1FQqxf/jJOBHySACnn9OSyR8guTP6DA++XWMK2Ikr9Kw6w9XKLqX3LfWLzV8iJY4KQemv
jJfbWgfjg5zXd9SMvD75zfeNJStwmdjobQ0QAhiClLHeXxkA8qAETcnthT8Hg3h0hle3rUdYornx
R9fqk8B6diCtcw7ILosOM20p1tArT/vfJqDDfXXsmingywoIL5FVeLiGYQV7HoBv+ELcQsmRGDjQ
/AqYIsfisb7FILigdsA3zJg3p5bBeZGDYEhvWYWrHwkLSQDc00M/oRUNdr8hl5zfG76VPL252BWS
jAfGIbK7wrIgNbhTuRWcTzBnTih69VCoLzwdYpEoyu01kx1bynLYBwYAOdtmJ5nRmnW83G5gUn9S
X2gOpx3pHWnnjf6VHTGKGmgDIAVc81Ce/XtwAwyeowT8BM+rLKjoDwSym7KHAqjSz5QMMiMtWAyL
C5IFqnGYn4qO2OrX74hlvro3ZQRGkGLIzHQFbOPfRnCxsXTTGxMZV7V/SXeOeXrBcBB0Ns8hsbcN
lI3oS2zXGff3yc9aW6rRORXuw/NInxxj/ctENKUftyW8g/byWaWpMV7SGQmNjhrV7dQ2L0FdOmto
alaBGNnSI24Aw4U4jAcWdxuL+Db/nig2vMcdW+M+aEtAOGQ+his5a0naFBl4xbA8vCRQCsT9/NjV
OKRP7lvLk+Ty/Efhf41E49gAn2R02tGEykv9MGp0APN52uINZ38zKnz28XUyU694aaBcdPfZaYO6
Zk6GXfL/Cudn6XHCKpJXTbWHn3o9ivkK0m5Vs0IS40qwnPdrKGJ+7C3pHYXy0Ly4eOS9nKr1Bm44
suaLbfuEWZxkvKiSBz/HAhApDtkBxv6+p1L166SBO4Y2vwJsjPJvHPPVL+dL+34AnOPSNPrNgt4g
hWNJW7c9cMB1FxQ14WdyYuCFV4oWw32RTLiSkFgEz/X8exWZC0BMybm4G70A6wXQkTldmnbdBPmi
6BT0qzgNeP1ouLZTiKY1WPkptyA1m8e9libHfeFmoLTOL3yHzA693bEonIFShpYs/ChqLlb1D1+E
SmBmUfz+1wIOdBLfuwDk2lAD0XINLEN0SWZ6pR1wJXRfOVn91G4XuUCg89yZlp1KZDkr2JG1u9sZ
IqtM+IjIExRgHyOMPvCmYK0ZPPjoVlomjnnfEtWOQOqRH3pfZzl/MuRhs/toCkYENxxluYxEL16d
76oPGwCrHxae5aDw13EMKyIGt92uB1V/PHBf5UaflUqCwjWmIIVWkzgdaL3kZJp/uS4DLhLL6VP6
A3gr6SqV2j0EFzlGsdoJcL12bF9C9lT435Qk8VOcNh5riFh35tW7/WT1DOghDDa3fZxjU2VZCnh/
nA3Di9X8qlkd5IizlIdmXZ27Qk3o+fYHf1ZjmOfT4JHbCWP26pWEe0/lZCDGxxvsW78306eyj1lf
XyG0hzmk1v8ZIFBUR2VVYLmZyaHfm28432rCCcLntnYOkRGZCHuMrYEf9WRkuh/PSIM5BxDcde4t
3h1/P7mBL8VDNxErA/zj0CSXC/m2nb2ebda3lHtWQsi619CKxLy+ZBzAZPUI7vCLyNOJMbui0uPj
vrwN4wIXrlgnVwQhthZbRsMTg+AdWkkUsQ1EuB4fWpFSUxFk+/gankhNRFDQ7v8XqXZRgv3/ucTS
j0S3UPa9uYgCR1uqGf9XpJFjsXxm/Wp44JTd0W+9lBFwvYgKstomIGj9lhDizKyq1mt9RNyzSw2o
1G7CTqgZiSWM7V0wKsdMXOn59Ld1Csysiz8MKnoYB5usxj4iC4hDN9j4yTpeOiy2cE2wTpSV4Wy2
bP9ABQTs/MWfQLyNKhhwkzJtYGLGnT6N1hNrWA3DHk/w+l8SCtdr86+KN179U2hibLZNrT3kbByU
b0Y3a/yTBDCvLa2FxAgRZ+TqQL6bATAZ9qQKr7QLEChgrdJ1sMGZHanA0jP+CcsmLFfqBSZAy87U
KFYEazYzbQOZ2Q4q8/q4YPB2Llma7jGGIjJze8NS2c29v4z1hhQjFz998LznT4+zDzW23PARvQaJ
86mvs+fh9Io169QmXrq9NugcB9PU5pIkmfTQDlzkPhkVIewMEOjDZIFz+y41qlJiX/IcwT7xf1Pz
YOcxf0Ps9kyy8wbhDR+ksvIp/9zRlTMyYnV1AhOL+fQm+e4zGd3WLRGDMGFPj7wOmAOx1+7Ua+dT
JLKbePLpJiXvy4MWHNro4WMf2ReaMRzcbPeq84Y6wguSOmgpzoEth9e7E9fKyopPz32V+rj5vMd6
JHQlWx7GXZEN5GDI0II+ciPHwRb68JuNt5YYuwN/MkuTbdyd/Y5qiSATnkcUklF/Xs6dJm5GKBOP
sVWjqMx02UvTGlIpYnaE2ML3zYENmxwQkUvqWR7mPv9LsHg0dKQ1mGkYj6NDSU112IHn4sAGzuHW
zRz6gUf+AfIt8BrzCykHHR870qJFglEkN2uGzrh2eUOqMAclcVG1s5L9Pnx9SVClfc+DpWVSkrof
+VY6eTVsWWhXJYvF3gu0u6qPF+vFOeaR2v2exsbNM8yL5WFgPXBD/8Nb/f6uF9qD28q9a7Xtr7eO
THzxIeUtLQlMMCwIJ4sEwsh+vZobDlDO7ilSSsrNHDJx6hR0+/Ozz6d4O0uhO88ANXadafgbMcYt
Yzivk4YJUla3a1nJMka1lmioCX2cIsidscC2h0YTUT/DLsKGb3Os5HYsa7pcB5zxyKsQeY+dy5Zo
7Y9jwN6ZHKKzkxYuU0yj4aVTn69PyiDeVVYXEkPLACoWD6b1sbNLkZ8GBwWv7fMFVZuRr/Dap5r8
Ws4KXYfdQOYB1QIBri2TQkMacfj9p4GUCL3ZIyJvi/dRYecnPWHFhd6B8ReBZysZp3CwOZZbjk6g
axIYh/9W+c/U+/6xNU4l5xgAAjCjNgcNBE8Xn0eb9/S6M2I9RtjNcmW99U2rpK4B646D+2s6Pmil
1ly8qkHmVwyLBhwGkX7g7ra+IsVi7RdZLj5n3m2fOO3t283rL6L0DD92dirvd7XiL0upnODTYQaF
6ALJBIl4xXXfkAOhrIMAoj1Vb1aHy2RugVDbuAe3PAKzHLgOfSSVppRnp2eLZSFHeyvRaOVSBYVk
XCcmgTADmJE0M7iJLXZioNd5pbjRKxR2QOpvjDUGTxyhZdRRJlphocLkU4ZRjeoB1GnFEn0V0kwN
zYFS4M0Q7PdFutr+YxidzgypLD2Bu8vxd45mrMZNlYGT4sxFXXXQy8o6KZjmMCqimwx1xsJpvjqK
JMwTnc0lCXzgVt5/OXIgI4kPFo/rcsuIzy5/APq/GYm8jAPAC4y2PsZZNw0WfIz5MXm7Al3Bv48E
Fc1TPBeAACHzpz/Qz8SALU4z5jqVYTrzdcg+ZSnzTzuy7GQnaLT21XRi3KVsN7i/Yv6CZFSdlJ0v
OYu5DY4AiLwHWrhtK2y+QfPiYRIRSf4LVGeIHDcahqdc/ihJ3Lt5ngGc9vwRb86uXAaz3IYpuwKv
MSHOCDBOYELCotB5BwGbatLRo0/RnUyD4eGYgA3l8X8bssgF+wYxyZOeQYKk5mw/bTh4lo7YLmMT
qr5pW2i5UKG5Zuyd1OACQtaYmnEmncqfn3pficBR1MDstJqHVzvG5lKoDhvduy0Ikk4+MKEBV+Kx
1jhY1YmCaenkvu5EQaJlKAN1/77GbQ4l9pKu+0QrKncM0iVQuFNqAU9/XxoQhFRIJbp3FOgcsL4j
+d+15eMfR8+/jsQ4dOC3HDnsn0styjkwKo382JPDVXKmEKO2aiy6hQD6kfMHtQ4D2x34euKbC/ih
fkFiLsGvRaIo6WA/jX8TR7mwqHAq2zfbBYGdOXHrTjVrcmQJFIEgq1W+cC+XJpSFgvjTUPe8SeH1
SVVklj3Hyn/TpvrqV77J/15tAlQxHdV7pha2OPzPt8jnZwY0oVT1JzULtQNCFcwUlQvAUwvlhO6J
zv0uDcbNsc+sDL7kL7suhHkYEP0XbMuBG/LHv5pfy63PH0OHAyz2opt+k6L1kes1PxoNkLbHsdVa
KO9c6jdYqNTy6cHqIQ++B/AZrg5/Y6tWpsO357SgUZK5zDVYSFAg5YkaQxkUC6JXCZ1G+zmk3Xdt
plwNsEGBeJzyJ67qt+hk8Oj5DMw0zSrUZsnMH17yzqBHJKXNNEYTX+JMgmL9ZDmSMkCClJKQtOjL
5R3/P3MtU7L8F3MPGIf6J/mMBFiggntBgsCiuNjxYFZXg1bYNc+yU/g7EGlQbXIQ0IS0gZ29X5EZ
rjnXsmfRnEWbY/9TjLahDoJTvbZ4jW0Tc9hbU6t9KiUSPjDcoTRGx8ZEoEVUC+a44JLWSgGNyhD0
iqbuUXL4GZE6jdX2x6hCMEGRNUEovsMYD7anM5HjBtQy4j2rzhMt+b3k+vQ40US0o0QN7CVfZ8Fg
qSlJ/VA1WyVQB9ky/GitdW838faXX3wAjY5yFPBbYK7l/DWN4LUzGkD6qBdD9tEoRk3mVf1e7Gmh
f21yvlJI6osLNzkTys+cY+LTosqUlTfGeR73dqKofMJDqOATKgOO12vvaTNDg8KVyTdN4nqmmviR
qKzhoTlJSrBrr5OFzS5XuKsdDYKU/NYy+kZ/wjRZ2uXbkYUs43IBR5I1bDgyz6g6+rHVvYLRESGi
lgAIwB9WBN6Sbxkd1ScsVZ13BVaizko+25lx2yvAOsakFY19wJkA1g0L8TE2eE3fXkOL1RXaqziZ
h5H/i07ZW6/R5vSYG5qAlmVG7MRv9nz54reIO6DKXyJFSDG5EP4Ix1PrU7PHcX9RhIoGfvxo+zgO
RM2NuWw2NE6kvvqnv+j4N2ltjwz9VemDjPjAaPvjHnMiEQ5jqEqVigNPdtAeCnSCSyjtbiZGecZO
Bet39gD8LR+Lx77/5guWYN3Eg0szrQ8Jf2847dguLEQM3qdxVNe1ZpUEDxHviny90lo1QRshIrin
CZx1goKKV/4EAWQzGFqtMc53JoJnG8JPRTzZyYze+mxOS0HVm/o7rKbMeIaclcHc1yz03Bg/M1vn
pK/yFikckUzUBWBmx7FUQP1F7oZqxb+bRwQVVRHwHRCHorF6MTPw3iZ2W4uVXBuFvj8+Fh9zcb/d
yz0XYyemB1GqMdvMC3h1uxbvplNgokMPMkDaNU/imLud8Y9Afs+sJHFXQ7+6rFEM/VYNvVDKXfRs
J72b2rq+EWt3YAnNhlgVvttDnq6V+avI+oyQdssBgEw4NmjzedKEspxlO5TyXgbBmkTisMRRZPyp
2BS/S1fNQhiinjdcUj9n5Y4kbbth31ksiRiHTnR7qnZ3fcB05ETx8x2H6QkaFZdA4TF5yGgalP6o
9hFjp7Vps/e9Uz5iXBaCxb3VmolWObR/kEd7qmPrEaE26zJpc2MnQ50uvMDxzr3Qw7qJnmHOOabw
66HPoBQ0AxTMWYxqf2MSiJCBBuMwkG7j2f3y/X/xB8xyzqV3Mk0XEwwAwuseBfgBp+D6/N/1cnTn
Q4aSGQr4ky/JdbByWgkMiNlYD5VDJ/vMJHu5SAqT8WQchGcj2gnV8u7gJDqYYU6Uyu6yjhtI5aM4
oWRBRnkUlzuRcZLUJMZMA8xzKPkw/hAAUCnFqe7+AD5HjEK+werpFkqByjrNO9AenAOsfGsU86TE
W3Q9nV3eerey6efKWFE0oGQ+ndMA2behbLbguZAPTkhwrMys4JbApcflmaVecM6CJdWbEVHg6fjv
gg+04sFQqb3Zb3QY30RFbtZZ6HuI05QnVInsD4WibFmsqjXKUKq7Pbi2FD6nJ4KFHm5MhsKTxnTk
BcHAqETAX/nz323vUkFy9Lg4j50dzyAWywWJw9LiqX5v/LGr08KFYBzXNLXbdFISq9SYmv11N/wi
ivHeGz+Pr7LhW+el7fUBCH+jj6naO9owRVr4xJYhTioZ2ktJ0EzEMiedS7AjxD8g/PJLWzAidXQl
fwPcAOyXwLZmq9DLLlP8CbqwFPMe/0yjuS755M0AqccYHYiyQdnnU8aoqU864te4yy/deO2hB/vm
XcKunICeWi3U+pIxVIyKAbBS6rtUXvAQRNTsYdgqR/I9M8z3sOlI2Th8q1VRAeR/iCGupVYGXxXT
WxbEgFZMl0x4wd2sCdNXdhRSmuqN5AKg2oF6QGDk8BitkPEpAxUPUGjMGUvuLtQlL2N/4grVafSh
hTkDQKmAM9LSHTOegzJrN3VZbvL5OVZ46HO1SF1mb99rs8M6WerszvEPuwc2y87f8stGwy/o1PKw
EMY8n1KMlb6FDk3FkzjLSULLKvRaYnL8yzPqEZAXrYq4/HP4VJXChy6j/ldg9/MlBG9O5oPIf+Qq
MWerBlXaEW62GDJJxXtG9ff1Gcz9Jr7Jbm7fWfJ5d8m8Nv03NbpGKb/9DqFRt8fx369l6oYgcIUY
IsKN10JSuut8EOPVH3HIMoTTsQS+YUH3Cw4CtmAX+gCcZEjgwl/EygacJzv4tl4+0bHkvz5KuBCq
Vde0rDeQxcd7Hy2u5i2RgySmeLIdd5cHgW0DXV5TgVwBIrynSTutO2ie//Qro2KMTxROatP/YWxy
iozYu9m1+f/7nFqh/jXmCBowmaEdEjbpaTyPp6QIBiSrSvNvKuqS3pV0gvjv4w0P38EFoVTnWtRr
prFEuG0gzszEk/cud1ITJsc7yNKUUOFt4S2nagiXnP7Q+9wBIcNNzaPXHL/qt2EQ4ZTVGBZOdk2E
Cde6p2OHZhj7+fzVOXZIyjRJDiySii/TDfxsloon4We84CBdUmJo7z2n5qgGwDgpDo32zh1J6BAI
uMguEQ6xUn9o1nNQFDE8/ZxZtHt7uDA4kqNIuGKt9WP4U761Um2hAYVXrkUxBU0ylvhH50cyUFQK
nJa8S07xIq18hCbSjRbUs7RkldMKa/uGNd9Iy6j+RNgFpYFar4jGNniJVMVN0tyNSmiNTsKyindQ
dAJvFTq9q5PouOBLEIsbn4CshFA+Ikc+ckeR8c2DMMRRfYO79eyGj7SYJ26YjllK4z+9qfA90fjM
oXcY4yoqfQNasXOJBQgtzjyHh1O4FZ4iD6gC6JaVFvwmOV/VqzGfD6/T8C74A2czcEc4+Kn2YbPp
RqcgQhnDAIVhZOolf8lq0Vl87wBm7MKcX1tFWZdFE1/E4BAPgPnaKJPYI8jOAWS7XmYgW0Y03QGC
6i1b3sHmxWPNimAUFpnJ0oSA7gWzF4BzcQPc0X/MOpUYmux7TRLwuyHcIwjguV1Kw8xWgCfF1jo/
ivbX25wld1zra0rvUBmDor4QpO32TFqIKPq7XqCVwCV75ZdPGw8T3XQOO0N5azIRWQpAjliPTxiT
ILRLVwbSOAa1cvG1Axvn7GnWBNsQSv5GIc2137tqsF1AXwMxH8ju9pXNVng16V7j4cbobJMlZ8Zh
SgFknpgOZpB5DXcK7sBor9ekXYI18rxpNzJ7uPRk1LwX4nUlaNVdmr+6N/UuyRi1VbY8MYLBihLN
SLJOt1QWZTtN+CIMChi5pbd/yaW8ORUKk3HvYHm5Qg/t4mnO7p+y7p29nwRn4I756bX5XlEUWiB/
cyGdQYsUuct+BU5X8NRM9S0MER/yNblcWc8PvLUkTYqQsw0S5n2NmljqJDDbEqffXZHphVlHIktp
3WWMLNbQBNBSUMkvioBlAq1I1T+6ajrSdDMENTQf54u1v/WZkt7nCPB7F2ImfT5kctBKugHzah+s
A7O4QyvY3jlsiXKm3CnoeRJhPS2Y5DppnGbAZYUnjTzWabcZtzyTuJ9qjA154PeeRd7uaezUIrJ/
wF/M49CZsW83QCqiqiau4iL+I0l2T5zVAudyQCyg3fHn6JxW2Ph6bC9z2rwiRG9Zl+Rfn5uHfs+y
f8v5u/dr5mH+Q0d87YtPnIj+lL7njzO2EmekskG6uqdf+DFYBupRTyQ3WgDZB2fkDwOpaOideWbP
UeFg91L2mGQARH0Hy8j8QDIkiLBwt9NE/nCHyJLSmL4UG4QtlUU4KHByPFGSlX4N9ju456Jvp2i9
/HZA1bKd89Clo+uUhsZ/0qbxC3NN+G1GO596RGU+ZUJPfG5fozf++Odyr9oowadaHOVabc1xyX82
72b4DekwOOL2RVwhMDNFplbuVK/e1eFR2T5C3hsKsOWc08mOfMcKMba+gDNUJzyY6vMBSJ+VbRPG
SjMFKCmTcuaMIVqz2HNEa6zhKEm1h3UeUf8FA6WuKakB1LP9IShyPEmcHjFvwKPhXRHLLOFZ8Kmj
3THcuV3k49x/y1RejL5XbJeJ/JLaEh84KcgRcj1rgTaVqbFnypvjmS7nMi0zl64Qcl3nVWtDioGq
9ulzGZPiPkHYsFZ2mSp758rJ2oAc0QKjFQ+kyV/iplHwAQkb0GDqFO3z69g8jmAKc25OecnkebpP
89Shjzw0S3jqbSXjfx8fNRmDimBsEa0mk/K5dC3VaNlCgUuYWiT/NY78yMffK3Ji5gNuEu/jZNnx
DuHXyGGMCbZimpa49+DlH70Ar3rvuEg4IS8ZGxuu7+7NKgNdkc9dbvz7Ozjuv3KrNax9NLv0LLQa
buGl0UXslKEgGaHaMoKBlYFBVFFy//clgpWnI5lDHi9a7y0ePl0rjcrt/CCi3o+ltq1APGZskdr8
5nF50u71XiQHYdfHQr5xrpFpQFyUvVd9BTNsppXcPeGwYvhKbAgMyzbpbF2kyIT0W2d7yJj/nQgA
hoY7WKJyp6NrHjEVreKThB6eyyaUvvdfqA+OGlldDoUk1FGsH3+N8n+WGI79DvWslPY1shGLX3wZ
2q79q3wX6uiXGhtvPF58V4BoQcdjVxz4fgb2W3E/ZVcYEvG9nSQd7wZ7Kb0qFYqMirzbpwrU+1uW
JzKhiSbcPxfxbe2KJcEaAVqfqKynMyr5bYvAKJzXxB5H7+/dm5RkZF8UE3F9hlc+EGzH9dR8CbzM
JUwtH/StK9kcFtkjS34uwT2MKmhSLnhWkol6Mn8bxxrn+c+x1B+bhfwbHGcbaFHyS+Dm4MHwdp5E
qsslwv9R1aOgQTzuKq0Ge17BYT+CflVR3m10St+xVdoECtmRVN/kEpUE/23my5PWEaGTD54bPgwe
IJxytW7Gug/T9YIM3qxzrfuV+BUDKEDjKgOrv91dkPnG3ld/h+aCGKVefLgDLbESrooRWi2fMtzP
2/lhoZzHgmtHxHc+9RA4DiKiQGfbhd5YQWvCxFtzX09c7ZxBBF1fBMpI5WCKl7IZpp1qGHUAd0I+
sFOgyA3/O5IYMYZK7yHco8Wu90IgTlNwaYdTjfgSSHXNMOqARmY63/hMXQB05cacOAXJHfxJ5lcz
be4SIfZSYvarOyx3nr6kGM4cIKRuPPSvxfc8W03jYFdp1FxHgEDC/M6gdlObJQgDINeJxqWsPcDK
A9+zbJ649fgg7WUYSZoOutonkkegr4of9Xo0/8femlWxcCgFKJ9XYDmjtxQx4tHKdBJxc4Iv91mQ
Hb8UmtfF8nx3w++BAXlh90j/ZYlnR93T9TNSNRx+Gv+5Tckq840EaChliz2LpLxhRS6SETblaWZP
NH4SdFmgEJg0nnLCnlgIK5z02Z82hPckNRZNDd0wdiGr5KNuWyho3FpEbRacdbLt87LSvdszF7Qk
hhkwNsSfJToIU+fHjUKskc4NqcYN+vZ1VQ/TFa2GLtJjWwmWYG2qZUhYOVWUoZUlivttfs2a1M5P
8bhKq01rYbJveHJKCJ/qWZ3oAtbAciYBzaDU7B/i1Rj1JzmSLRKdpK7j7ve6RPMCrBfWGiIReFNc
SJQXk4Kib0n0Df/pp06pzt2IX+itxfdnFWQCgwKoB6V7mxXltqdaSFP6wRIWZDV6/IGoPiGOmVZV
ytkKBtlLA/Hy1hU6GxYMhWPuH7Job759yPb0GVb6beYJFaZ3GyYUQcj9YpQMwLdK6JMJRbUmS6IZ
PJmPV5NfsaP8K6+EhPHNLMpJp9ltr3RpT8QB7qEUti+Rb0bFFiICcgLIsc4xw5ln/gkPrcZOMo1f
iFjO+xp7wv21FocO82jMqTSPtzEmprxQNy6DPlQFiC+6+ShwT+GLd/Y/ZtMDQK2YN2DtV3pcSdKf
bDyZn+qphUi76REEJzn8ZgvqEbd0tIIwj964yt1Y2SEUtM4uwC0pPj0FyPJhX8ZeDz23NY8PTpXJ
eDH02ryQaatMH7I1mJV8GT5xZImW+7v1A+GNyf1opM2c8QEXaYmAeFGfvhVAjRSzUe2hm4Rrz3Dr
wF/zEbkdlJW/oArRu1cbDgOlXBUhUoCL4ud1pe8kw8UASFXA3kt1TkpzT8lPNwN3UjydJbzDVz2t
5cD5VnMvlgCIqIBf1XOxtXd9nVnS7Vxz/KQOFzq7UYaHMu7haLkF/7ULzDQQHL5U0UZMi4o7beNM
JPx3lRk2RlXunGoPIqkfeG0o4qCJhp9nYfuiXVGb59p+C3B2GDTw59+mgtI43NweRjLIVEAEycgP
2/6Bx9OXfAAKBjNMu8QRU6OegyS0MFpmNxNWyj7E+Tzd0lEEdaWjrPsy0kB9UrvcAx9sOR7xvFzx
B6xgbAk48Caxy1/A77o453pHLMg/CF5SR7JIt0VDmgTA7CbDnkB4T1QQ/yHKDPPs5Z5WY3QcuaDf
Hqtcd70mddm/uQy4DQptsB4zsiv3RoCyFnWwBWZdskSd2tKnbaOXrOUeDUu6nfaIXmBXZitW30gy
WCTrBAQ9mDM5ltELX8u0sptGJQqDb/duTgk2YMx+HynQcqzPhA/vYpyveXMObW/ZGZJlgZ/Vo95t
DdHcCR86nArYJtemf62aWpN7dEXKI+hB1pG17MAKm2xXzRS55lG2zqOgvem5d5yuMXt2h5lrT04y
jVPQjUWvxbTIFgXxGuSL0ceVTLf/DUpUgYKGvPM1vF9oV+XZIzyti4IiNPGQUnmjmlqISIl6FhpN
nhexPXtjQ8FN9e5Jaq0aQPTWv3XFc4ClopeBjt9rUFeLZFn3nSx2cLPMar/5R6uK3QBnMzJGrotJ
xFD4c0Gr4oUsch+qr9vecdB4TTAzkYSTJbqil78gJm7EEjmvC9AANCke+rarylhble5Qwwy07tsB
H5bbgzg1XcKmGR0lmEiAr3h1/U6GzBOwl6+bTI3pAfk29x3nUd7qPXYSs2M1lqgXusoIGYJWgogi
ByqrfFL8CTkljn+pXPME6BcpITZxIfUwF826lSFxlq0thindTvxIQm4ENfWsKzaQiGK+18wthXkW
xRgzd8iZmE95/OqGP2EcLLFpOY+SISnFS/gdEIRhjX35M6O0n/4RtNK0Ubt4xrodG3IVl2Sxxkj5
q+5XJ8JczZt7uvRC0gy5+PMKMYZfKji1MStl6i4HNTuGQb3LNeEa1GEPWFEov11WvmJ6OXARksk3
/aRNEyCN6czTzLN8HCspIJDbes4j5oAvHi4/q7gcvZc27iw4Ly2o9oYIwirh4OEpU3KxzCNeS4w/
YxDndqoiV3Jv08MfbAcd3UhUGuqAl0NEqymTQbF7Pr1zPnwnfTQkOz8yhJLJg+B7VPIO8XOoe+pK
3CX8wC9YmOJS3Tt1lD36fGr/jt8RLdtymBqirV8fTgAJ3Kb4zakn8wii3DwUqX8nzU/QqJuu0gJF
n/yUYql+gV/1vMajPWyaOg1rP0flQ2WWgJ1ONF2SY0seR6XjgNqyP5FYb4DUUNR9vwx5kiOXRKOs
j10YTCfTJ93+3XKwRdp400pocjrm6GlOmEM4X6sdprFJCF43M2MHUQbwataMiHDRuVn5XKhggEez
uzv8m5/elWudpTaZrIvmjNHfgy6L5QZ1/sZfbUBdqLSHr72saRDPhAU80xu/mNUcY1p2jS/dl4X1
3u2hjD2I6/lE10qm9VOrd3HxjPdQQ41eZEZ5Mt8Cyo/aztzePPBQeZH6nzgKN9e9/FgQ20b6ZYXU
XY9emr7HgctDbiqxFFoevRBH2VtEwHDQMY+kNMd4+qltHaXMX/QY0b1hpbO9+z1NcawX/U4k0oy9
eYfpYcu5sffrbvl+QqNuBxC6coaH8fZ0lQrfWsSpUTrxnkwa1ZhpuNCVAkQZ1oK5zqUC9BSQAu03
Hk3YC86HwDgXzJpVLLaitUeUHgFNBc7FquahRoqNoTtTdqlR3wkgWTlDeYgDc5FUex6CkstynZqz
YhT2/9qsOvq15Rm84/jdcgrOWkwfLxD2LivuK8bYKilSEcqgQ/cJVh8zluk+2luJuaODCIF9cSXD
HNIGT83ikREACijT5mLD9npxBcn3DMO0tIqB80QRFUesZ4oZV5lEQPFhKkK/GW4ZahUOuM+4G0Gy
8euEYjtSJ0nzSvy/Kwk9o9VX6zOeX7fO6W0RbcUj5jZ4w2KFazji+1TNhg9ao8Hf8dw+fEV1ABRb
zgcm2jyjcyz614AgbeALTn0DC791l45eYKwdVJZfIs4yqMSCi5x7vqPXfs6XwMERE1EzWsE3Yekh
YOmEWcHgRi1PMrpXyKOHptLY85S4F5u7aEq3ZgKSVB2YlEGa4qDGtiiXH+3wN+JV+xQMAAG4YMIc
AN+s3badnORKpLzpV9gn+KcZ/C/VBvfhESINbYkGouJramcLQNHnf9eZL+jQ4r/cOJS0tM/AoczJ
Hq9bp5rtkW6i4UFxPtS+qG6Ynn9EqxwUGhZlxJ7pxe4xqqBgEOMOADy56cg/+bccxBUyperH9OiW
SqTg5kiZf8IV/i12o91GdukjSFOgUB5THKOSs+28lEpCU1jUqt5T+v7RiAgv34NazgADQ5uXDvOG
AxSii9f9035ebjbU/mB6oxIfMQoh3EKX96K5B9rq1ngUE9dICxQZR6M2FQ9oZT9i6JLTYDk1ukt4
IzA/hrSiFycFzCLfDDWkyaGPPEYM6K/8bsyIe0R0SvFfcqkiXlT4WyKp1rpDO6bDYbcD+LGfRyJR
szcl8RIUgKkTpm5xNEaaEnpxYimKRzEXJ8VSbbCAkaiUIWK4CZ1WQKGp38qvRNpiD1o6gIvAYsTS
jH5VicMLHTwGAnjKs3745C3fWNByQkiH1J1WROAnc2V5WU1A1zbgBv0rrgtwL4v05QHWJ80zAdAK
YCXcaVlD/9jRbLljCBINHrzpQUjmq/1EZ0e8qcaKhAZvPwwX/l8P1IeD/YPyKT77wsoCezoDrHov
EaG+7NgdnODKwrrCzoXDf9VBn7tiSTNcMcYJc40hVKDsepFyld9YQZnAOzcbuH9X8zNbvLKXGFAX
BN6/fWu1qMHlNPKyLujutnGFdff4aRaigSC4ON68oa9vkTJau53Vjh0lUPYzM1aJD3tdNKBd5fh4
bssjsr63mymMFIFRyfdPxsCB+Tx+ahMphcn2qGOAnx2En/GxItoH6J9CcmiB46WFC2wg7EttNbxq
b1Oegvo+RiYGMtb3heas45KCwQJOyyc2IQEZT9f/671NtPE1HGIfUVvg/xOm2WB7F0XJahpqQbIB
qCGQBjkoU5gSZSJqXpn/eSa/aE7d0HD6LxmlBq7rmk3w9V3SuJYUwv5z9YMCcyZxh5MWUOmLS/et
Vg4+teEQ8co7jK94X/4IY7HY5dYNqtAE3mhuIzNrZVQ7qJapuVCroYemHyDNAYqb6GO79v4gCZjV
VXayIBMjXxv6Wm7vlNh5QIZNK5YkGbjx0Uc1wn02LTXBeiR5ak1WVaMsLwWSnm2Upn1VR5f35Wo8
7bEy7R5eAd0FpL4YeFJFzPEMyVayO/Mh/Fdnjer5VSSXYdYMNJIEY42JtAFRuYJy3uV8S6TUtNMo
XjNKqTuodGFq70TJq6b62BTsetf1kmXJf5vTMD3RIc/FIRAkryaMru4GfQyuMYFq1NfvaZGSg3kf
30wwIMWh1VOHS7qM5ZDDRVgyQQJky9gqhkSQ45BKjApBIIVE6Utj+NPezX7lsm+NgJLpwJSu568I
mxX1uwWqp5NPVfb3e6klek0cMS+pvdFPpn/b2w75OyIHi3KHYgkefAeENKK3AcCSs8mm+F7Qe1Qk
JyeyEfsltZThJ75II+MC/s8q2NGlEcf+zSpo08gzYXI2c0k0JyzkWuPblHVZfFnBbkRJ11NVdsvF
JEv5n5baH0NP9A2pKUVeTVk50NhRkdCgg/YnhEYqAhhEX83np2bttPLK+OHGUl1X2Q+RfEq8/Bld
4VAYiK5gg7xwBU/BYDS6gqZmtEsACiVIoUcnZHpDsr7AeEweIUqVla7YgcwG97H6YcFYNkUmuj1X
tvYh/S6h6gA6KvvEVSnl38+EEPzapKlTD8nBG7UdnYEaZBb517lNb0YSLYWtYZK8OycPZCao9LO2
DkQXLcaaQmAUs6mPkR9fDrqIv9smxUYbvhlF223roWAYMdrCbLKjT1X88vXUsWrpinUr0w/ZDdL4
0lDPL+G9umhHYfRkbRZs6co7xaWetAZ2PVv9lA0hHtARDdTQzbeK27+dnDszA3oitifslRTX2aMu
5fm0MypDrTrJ0oH73+zclseW+v3Fcx7ZHV40FXL09VGaOXnEa7nOV7B1EA0lOtjn1PAfHxR5yY2S
B9TFCOuzJFZq5OnWqJrSdzQ6PBYFkSJQlT0yZqEn1NWTbrEJZktqXV4EAAPlgdHxPqGqtLAA2Yo7
YAZE6y2zstsuU/QcD5YFklKOrud7f/6RHJ0Bd7AeK90hzyv/At25zj06wtbBVNFJddBzD+/sIxWe
uolGeLWHIub6nC371EiMXNt/6S4S0Dz+gOh8HKABVDB2fGPetSNO/pSvw2BgLLELXAiBWMpvjz/C
GnALfrZq/ICoa/6n9kjKFZp8HZONLuICxLd8gUt4kTJIKCgL6+f30tRSLO+N01NYZQBSDaHVJCBX
eMmP/qKf9aI1Is6PsKJW3NyBgYELUm4viJxy4JdBREyDKoDu4ooyJguw9d8ulL8BFdH7HNUp2cMJ
PIcv6Fs/kqq7WEBhfAxZrvg+StnMAUMrETaUuQYKCDJresTIwb4FHX81YekamoPmAwM0HdqhXR6Q
HzyURxYbyHRZaS4+esDimhF50a8MzuSHZkjoFUb+USVZEGzjoX8/J8oya6vbRHBpMBbe7haB7DD9
xzbq7nT1PS+Cnh+x5HQSCyZ5VuOPj+dmn7cIWKIuW0EbR18bVPsN6rRaeJbYOsWLWL6XDJrWAhXo
tHEQ++mIJOUcTLpi2V9dZ/vSGs9Pm5WSQF+4mU93addx+hJyQKwXOIMdE50hTWCDcnneS5b9alV3
vtL/AOv4JF/9LeCqbjlOA8OoXts96IMDWmaWmT2gwbNpXOXh0LvBH9WrK7FxrwNMEvpXC8HksJhR
SPvBl9QdoxwgV9jLYgewyAgTG8/z1USSIwygWBqZHL7W/OTThxStgtO+hsyySYw6xf1FMQUqBi3E
5fGkmKyZVXoBZkkx1OXGuK/UZvK4w8b3pA/FUkPqJVB3SJaPdRxpHDJ0KRxUddLAH0Jn27Ub2uPT
QnvzIpYaarkbpJ4rqVbM0WEqBCEI0blr6TVxGd2obkZKFcIWE7rG7HWPZng9SxGUJ10yBwRbhDSW
G+78N0bqdJedbs8K90/u+jL7nry9RP38k3zAlOy2xVu2Sm9+TW3oYcujym0pmDLubBQ03GTAwmJy
aIDLvnM78riauEwJmmuQaI1yAmajqpU+XaLohOr2QJAglGVsCW2VF2V5NxnreNheDovO16rg9z/l
/GU+QMbj3AyhmoWMUq2f7mbH8hwppAp7nKgnYBzlOLgpL8DQncvipZxXSslT8PtJYPeNYqm8m9rs
HaOhcnOvcrDjNDKssFYtQcJHr/bYNIMlDojKNZ/+pAI36GX3QBQDSs6o8w0sA+Ekjm0OwFsCOQJq
ZqeVmA4HXSJO0wEBxD0c5QGSNQ/FjDRKnB+Dy3U3xLOyWEvsbdBaM20/jzz/WpErIVWbor2GX2ks
weYeV0sRZnXENrRKYvSPfBPSEKQBD/Z/BPvY0rxp6kPM1NvXi4fa5yWHZkCYEKTy+sdD5PHUXTBr
5vsiqNvbFbHWrIv7jTXVJLRxyVy3n9Pvd/mwrDfobpU0f/1f5CxY/ae+D6eLWvFiZFC8Qxji1bcz
Etb77FIX5SIhb9uJofGtwKYRn8GHv2xg1EFtkKj4BdMLGuW8zsg8yToWsg7NxMH3TDcsTSyKlOi2
s+LnznqZXiDIVjvCGBb6k53zBIf5qUHUT2ai9Gk5djpx5OIhUn5DjdbvFekaCMxcCI8EV710U6sV
YOzvuaFhb/dFAIIORuJugG+OmQoBwdJcWWtB6yYQv6d9kjK8E6ScybpTmv3mGzbCF2za7RQ+oVJc
J/9qcNf63Y8fEGjEvYAdQc7vMX5fIP3JBp/jJfz2aWOP0byf4kW/f0KbMyeyn5qAiWykYdfsDLWX
Gi1DxPaNIDSSZBvFTmY8zm65iM87MJbf6RrvND0IeSy19BxzEsEW6dmgetXkbpkj+1c1MGej7md3
id7MwDQT52w7fhiyGPM2lQUuuRWR0ZfplNGouubkrg/wdwIMms2ZNVp1lQS2fBIqaKClddy47ihO
nyAeMrjtr3/Ck63grAlzaiuMx9x/eMucD5EuR1HS+5bGahV0u4PZsBSo79jWoOUWxeRsG0ERRwK5
lq0Z6JKA0peT9yQN3hPMHU7b1uHYLp90kSVd6FWDchlzN0eeYSgcfr+9zJp2ff30lM9Hap8lsrfS
KRWBKsqS5BSQRgRg0tFN+2NTSRFVnapjr/XLWCRbQyC/B6H3spOEMHqh/TJngQ1bd+pbTfMFeplj
sHT0c9HjjRGYb5hvKmOHorjmmWqk9Y1n2TxBEDji1wzXGD2a3oelraQI5qJfUc64RRacgMxbEZZn
UbkTEK8I+JgvGzlu9v3JznhI3K2I0jhcrY6np0A5jxAWEzipGf7BD6Wc0vGfJo6uJW5AFPc9U5pF
ziZHrvBtK5tUqxPjUNILsulx8kAFBxxX1obsQArMVBtaYzQ/2nsivo/ZMpCzIDM+r1/qR2TGpeSw
+KMr21zQYXsktLjsMWHYtNMukFgqnIefS1TQt6vUePQ/fOVgZraZb5QThh/k41gtNlYGKcUT0rJi
DRxdcdDvVFUQGNoziQD14W0wbeW2838OPog26TzPnLkT45irSNUTtKus3b9YNmS8MBoGpVMRUymh
OyKcYZnsy+DqOr0kZjhyVb4wOpnYk+K7MxCt+CtvSk9Rgt3CQY1XzNKoQVtJNcYu64uYWyvyZGLp
8d2rGF189NmTYhYk+BRKfxD22BkkBd761HXk81dVho6UVWQJyC9DT2f28kp3g0j0kM7JVugB6oxa
Gz/bydN5KcAII0/984+yioZI5vLBNc7JcyFCoWhUQDIrRqEu/ZDcZeIqqYS3C0JTD9YX8GO2/RQH
7NvZEvW/zyFuuohz0i3MRpUfA8DL8SRwImZ5Lu8S1B1Fob2mVHD93Ouwe3r2h8E3FD51yW20g9er
TVlS0GY+R0cl59oCOlegITEE+XBWjPfhYK36OoorS1W82nqLfaDlQMPDewA6JxjI0fGSvy+6YRge
k2afGbS0fHj0BSYzyHneIB0mBqePHSy82ykKkZELDv+QQ2vBdUa6+Oa5CVwzkLDN6vDAQn+tvWan
OVDw756iZJCOfZoKZ8QHghGWteOhb4wvD9kSER956qcfVJ+DQjz0rfiJr4pMNu8lgRBo27gQwbqk
Nb4b1Brc5ylSb580SI3CV4Pq2fbuSK5Mqq5q3PO4WR7UJwdwgqisatcnpe/bDSCLw5dgEelMmHIS
0Z6bvGIGe/HBaMt6alq9o1AsfVzTYWWzXUXxdKhB/TSJGxh8bUS0pX4QrjLXpr+VKqaSOemMWn0p
vUDsRJU5CGSM3PfnnD+Uhdekgb8+wz+Tl5Pw00bVGdEl4xq8uMl2X75cDO1vC0x6e2xaHZQILCR4
3YHaNiNxvYCxXyRQOwg4DA0/tVWGWTxgOxdTt0UTrYf/uA4iimUY/sxcjxJ3RJPWCiQWD2tt2PyJ
VNFlxfHoQLnAUmsy3i8By0wsuAlVl2vRN5hH2Kzi0D06u2w/ihth02nDx4tHCKTSPvcL4+Py5J5m
63/qwPpzpPOpfUG/2pndTR+8A4PfIlEERTfh3cGGCHSjpzrAVlkmhOyKjSVXOWT4esGO+I+kjQdt
ehEHIQ+xeDY21WqLgQ5b3+Bzsp4bUk/D1i0JG5j7TC1c8IpIfJbDrIFcTFBou3kbRL6ZgkdWfu12
LGDLGpWKki4U+/y52v4EiPbNq75rjpYXOLk2UuvqJveK99Ak7XQHxB0ylKrdNa8dhvxH8ZbKDI3O
6ZpRGFzVP0/ogLKkIcS6aYRGGEX+/fP3Jru0txmtMJWt82UExWdS2kpzLZQThpCfNes8lUf4ueE4
zrznFz5t/QIW+oMGjFnA3WKiAXtCw/LseGHSKle4RpbU1FtFIj7gAjabFNzBj3jFiiroL1gNadm7
ZNRx9nr4XR+tj5+8kuIgThQizz2o4roRu/wZFuQwWTKYznwq0r+g7sdppQkkXzXrdBLc8c+14EeB
idYuZqGVEPhGY5zK70L3qBqsGX/LDCS6MnxpR2JyYMCGC6dgjmTsoK6vc9+0DQPc8AuigC1cFqMK
FKGPosfxp7zCKzdlAmWCY7aomgGhxfnYqdgAIQYJXt067dYx7h54ey0oWc3CuiuRBD2fSCIMNfs2
6KQM1TrXN6WDB0CMNWNmLZfOdttIq0n4x+OyzefiV6WSWJLpQVf7NqdxsZ9LjqvgRaarE9VMebS4
mQmh58HHOv4nTVVdF5tXjX8Tcmw+AFm7bfTw4JB5bLhP3oL1lnXrnJDkMlTDm7tr1pTx5jhXGXqK
cTD9qr+B/VgAPdjq0PIJDZkVWbTSWjSZoFQWl8zwxuS/QIUxjvfJNJy9sGA475dlnffgPzNLgmC2
bdmbqi5A01fKF1fnTtOJEd0MNil7vcZ2LwGamRkz+aS3DBRn3qU60Rzzrrxycg4cYkTnMEYviKvs
V0Gz1PIwLtBy3ANDhRTpHGKq3CR0EftcETp4NGH1Df6KofNWDEYJMqa5g7kBS2yqNy8u0Wpv5oDo
ylXXfDnbTNdDbNipWyuG/Ks/nyZymBSAbuTi+UukKyErOWHHB+v2YReB3NbVRO5P5JUXlHtwMVcr
Jzw6jYqLNXirJSqysbXU5gQDmJOsZ3EnoYXWjVuUQJVV9v1ZOrKRquVECRm8+IEViRRv5hpJtOvp
6i2yo5xgrPEGjfWQSx52doM4n5UwIYIYpPJplzd6wn6D+TKZ8TtzKhp2uPjJqCvj4UE8jfKw1ep8
hc7KBC3VEIYCOEJtW6081LSI2zvx8LG9XcbzkGn1lgSlsREkLhTp5vAMmMnOvuvJPvhn6NnvL9kB
t/x88YPLPVsZSxVpnL8vzNIinZ/U3/9HX8jgp3jGCbmM4lCb0hDEJ9+IMzsAd0erxi0tXF0dNJ5R
sYr+NaV5t0VBPhWvcGTKSNeYexNT0N/Q49kFglxBvvslHNiYiXR2rAWrtsYWqWJUhJxGGqHqKt3W
6P5jOp25IMVCazS99fO2n3DnJRwUnyRNJNAQmuWtpUmlEUBAdA96Bw+t45z6iNnEowpWycdjGnKf
954DiLNJ8mpuHE6Qlhb3kawGmOi/8BtCV09p5KcTmD2dht5gxhEvX1slImY2V7RnXoVn0hJymgux
9i90Br5Kjxp8WlLrMSY+4aHUthLpbMs7tlpqEwfQsukXYT2Ra6/l0JEid7ro9nPgApY3ozoWQl4i
Wi4G34men9zU1gqrp1AmJQNxc03/WPRKs+wutZSgaa4T33w0vsuCIbJ3o5D9kjXK9xI143B4pRCa
MDrZ7hQx8KxxDQi7DiaRvHXHlj0aqNI/kFFOOg+SVirbc1IuU281t+OSyrWS5piK0K37dh7DadDm
KI6NPT4sERiPOsHWCe4NWYJJJEfPnacc0yfVjmNNP+B0tMpCexvAQs+D8ImJFYYZEHJYAiES4KjY
6tmre6/TboNKi410w2g4+A3VeGObaJ8M+a4H1moaAmXKUiXX9ErVBv52ihMt0IXQRatWLYOgwbX4
xrfrIbKzCAKq+yHRedYik0d1JcqexbLHnrqzOGMke64e4DM2ucwNXd+cKeDQXZovcd2RNXg4fyYB
rC1trZmbCYTz8qyjgoGFUhaK9smKJs4xp9MDC8pCfKy9nsWNLiQTT8lClukW1dHx3Cgam4aQj1WB
y37RbU7Uu4UO+yjSifL/0eDWTECCypw/6Y7xhq3yvDv0Er0Lc3FAKAKzrRgcqDte82QRXxTNgF3a
7No7H+eogsI34TfR/MzTG9ajCWntQTqOMSo9JwkY8pf7re3sXnyr2YyjfjpZTGnT1PBv3toouzSw
ZZciyU9hUvY7mlsZ8GgY3UikvxMvRDAoD3Zo2GC/41ubuw+HiNXUd0So3XlQ1n0nJ6YnD1aMWPpK
/kZV5kPuQqOEJgMGz4yw1c9PGX7onPMPGCRSKQVJm8+ZTwh1jClH/UeffO4JrzN5sGlJENkoqFGA
pvtAj0SLtivjq+VJEE7iXy4EQIGNPV4pE40/C9cM2E1sWTO2es6wd2HwnlJUKZp2T6Nis4x7aZSW
LgxLXbbPU6UgW6QogDTKVZJvkD883M2K0mIL7T7DPC1F7H7FAYx1kUZEU67GG40GWpwZ6zfjZLST
VEqJ9KI9u3c2VvRuXYc7ZEXwfwbVvQS1EpabfxKSaRbp5++cWB3L4TolbCKcfSYdazEWnGRYgAj7
I2yZZAgmMySxj9MZHLr1QmZ2IUif6JiaqKzrFCkJQh5AG6FVcdilbCBTzGYzQ/MDWB9d4s0FqEtx
9zYrIrqceGYsDe96+fLBg5w2ofYMASYAREtEkFGSPzJWpW18kuqwuexTh/dy5RAD09E+3s3jSgWT
pu8F7MlWPJDBA1j70IRcI3K60CR/qsEc4Alo+3XtSr4fZTQX4rfSOrRSvdtu/LkZr6LS7ySXQfRl
kpt5v5hkakloclNi2rt+UdksiI1KGlO5ZCGZIoyl1gZ88fwPvCXAV8BRnhCc4tNLlgYz/jeRvhcM
SkBkpiO8MUldthCi5DOnnklNhZMEA3MdOIzZI8salleu6/GRTK6sX4WLrOBTxIY8LalutJh5kOmo
QiZ8x1qupUFIHfCQxwdNwCiQ4q+NA0dbngREh7IPqcByaBSSj8fdvMXWaA51KPARUVuJK3Vcqvnc
JoOHhRbT5NRrT8XtEmfNQ3/ZuiLb78ef225SGi0ICk0TZ4qF48I4W22CUmngL5lebiRBnTmKVjBQ
QQhrTPuvs0BAZKrE4o6yQm3xVo57Wwku4EWtBpY1NapDSv5KvO/44JC3ur4jriYXJyzTzoN9hrF7
MBxI1xiciOCYMrw8pA7o1GxFV8amvmUvLyDygpWKKlh0xOJ5+XKkHaF/2qtrf3QgPJRffHfQ/GFU
gCPJQCOrvxzoRCadyjguQAipWzEaVadtINVl84r4kaKnoDtujPCRCFUKvBDCYsCnAQWIHpDwKosN
BdlNhVs1isgBfy91qLQ/aO/q+NaeogPhXkt4gAcUkonehmslHcpJp9IJfQP4J8tGOGuVcHLe8CAZ
MGk2NCxrTtHPBQ5HUWN8dnfWhvvaIvgfDbyquvv2ktW5TiG8nLSmiyKqQOTLi1iAs7lzFi+B/cQE
PFFb1WKIVrNq5XJ6h0xMatQo/Qldull0ikpNWMa53R2CrpwDXaXvrH6qOzubtFGr4Vc9Ret9+KMw
01rbiLYHpjual4c+QjTGjqSwkg22Jydx+7E8qwRXZMlMDQebKs2hzR252vy7iCOEI4xZ5FJxBt9K
ZIq9kt3Lz3PkbbAFO2u+pSFQ7jYcDUv2+YwpKiWJhSA7In10e6yIbascKBtw51uKbGvyiTtnEw+y
a3VX9ki74MfuxRIM+BczJT50HxwgvBpC8BBr8QQwJkVqticWf62IeBi1Bn6YvUIqt9TwfprqmLM4
T7/ONyx0DYsvXJxtBeVdax0KYfSrzLXNUvvJthl5EqB3KtZOkHnivUDwyvlGdB37osTneu+iQfO3
SKg7ExRqc+Mk/UUQETnGzidIINUiDFZMDTi9wZ7nyjxIZG2aINA3kiFRaTrznkXbv50+xMX1pDiM
UrngqbDK8Og3Ou3B4VSEBcmC6rRpUP+fPMNVBCL3bNZieKKPam+Yq6HceVbx4nhVEpO7KLWuBPIV
ZoQ+yVfpH2gIP+7EK0MYslQcsits07hv2egTR/gHJhA0XiPBLHqJb7EBsdSC3ODzyksfBdf2lr8D
8aW72jjyUuqJ4Yn8XFtp3S3Oo0cgcj5gxMsxVqgxWMxd4duqFwfBxCZ8q2qYuvx99PlfapVl+pqn
vmgmx6twHz1r41aj7lPcUdy/x4RFihGWmzxPsASy28pAb25tAoeWIn6wjCLeMOhc7SwzC+GObMCI
Fk8gf2Vhisx6Y8pv3KboedCpLRYCMoFDl+YhLixdX5ZGPYDoTI5GMcS92z47r9LtGKyRJZLRstuk
VDPIgyh7BF9bDjDq0jzzuZhJTZgjWk3vT73fBIQNPxg8MRkeb2g1+7sDlZHGVcIo3FrdzdLBGJ6m
4aTDWhHWFddkyZROhRat39dCZrndVWW4ngoij3M6G9UU/uCl4XBPwQU/4Z7hMOh5VlJln6llZYKi
xEa1XwAT5I6bY/wZV3nxHpS5l63ui70i0aFaCltdOWQZfkUU8X67rh4K+uLpbQ9DG/5kQhtsxrkX
Z49aP3qLAz7IKklhcTwH6/2TI57OIar7mXkCo8XbJiTzYG1njLYSo5sryaxDHp88YO2JhTDz5Pf/
Hbbvt4oarcecL3bXOB4KeRBf6Fz0edgMz9cqoPa5YSoIVndWEfAfSZkR1ivbtKgNPmrd3EI1/Pcg
QowlcXD20MZUAtz0QXZE2e3dxdpF67lHflEyJUebAtbkyViWm2w377iEiiFPniRfqhWmqu2WHQga
XWTzA0/yUUaF1yjAlHSoJmYe78OOV3vjwzkiGf2mPI6XmorSE4fwI1EJCA9iWU32N6amn9LuNTo1
7uzfVqPU4ns6xPQU0vkj/leRawBuMqbTZElC4dZdAe08VSch6432mnxsLa3D+ix8XwO3IBh5XFZe
+IJJ+hAWIIeiciQVkH/hUQaEFfa0k9oBZuhYE2GlymwxByfJFz0LR/B/hVEvGSYDpotSPcBHCPYa
IfWZlSTzNJvYmC56+I0BZiCnt6c2DKGhbRGnWzEZ60IKw0RLMIvAmgK513lH9FiIvxfNbIMQHJso
WrH/Bs6sTejvNDbJ9IoUX4UFr1Xul2V6E/M7QeWORyyrvFJ26s+Pd5e6Aef+RWGYqYOfqzGhVHNV
p+z78SvGmy49tlAkRdThThgJggI/RXjDpjztNPFwJNJpvs1BnRveCTWff38/UwrvXj79uAXXKduo
2CggIEwXF4YvPKdUnJBcpaUTvuN+iDazrUrbxdTRCCi6+7UuhuGsZ7RNnlby947CYe3C5zlLhZvI
rtAB+FueSaCDsSEEcc9IRRRd95vwMlCj+k0n0QU5Pb2Y9OBAk6jAP9OhYx+9t2Sr7LApBb/yEyg1
8P/go/3PWYtccnpPRiTUHs7ZjzQuchy/4k+GdD3DMGIpWcNU1koa6wsZC+9CGVlFjn0ACSOHFCpK
1JkflWMewr2UsLZiTFGKe24p4LErOgi7E5YP6mdEnXCAQ31zrGKtZJwOR3+a0FiDRwSIr6VoJmbE
RtJadbl+klNzRBeA+v6CJJCX6fNsLbRB9gyEjqT0ew9jEEf654YYtLQLR2o7sc3wf9htblIVH1Lr
9QfM1jeZV32gABVqS6yZh/HMB9TwVyrRduZM9qldiuNkAhE4bSAetKUrzrRcHLmB3yADnTjbZ853
8eT5komze43ezSJDp+dmpdUcshvyIaU7BgAIIBRdh7v0ZM5oxKk+2f31WRUO4Dpd1LyLZ7sdkx/u
y2gBS5qxCVIJKxu7/5jPQaddjj2Cqz1s/lix1lTRJVM01OtSa1CKlX6+Q+yjYUyKbnGvoeVnoNyF
dhxiKzsZIxYwESzzYO+/y8yrKD/xl8Iotumi8JuUAxO2U/+nIi1dBMKmK5PcEo83+fNbZKNELTAg
HxACJozfmVsXQUsXJnVHUb5h7QlNBV7cY4KbXXYiLaRMX5ng0cC+cbQ0cHlBlZ9+tkhhyIfwM0TQ
VrfcsKd/q1Y7LWDk5bB/KTp6RZuSuvhqZUadJNQYUpk4boS/+jiZ8t+wYrOnFuf+ZdxQZLOuUkF4
rflx82taF+4/Xuf+BFYuk1qDIce3a8hp/u/AcmT5HwtFVmWFb7ia926QNBWIYe8RXJTQLX0iSyD5
qPRSzbEaVXnK9FlfEHqky25mNqhniuygp6lP2JRgLNeCNRgZJerJpJSOtU48XINvTtUpidP4EezH
kfa8W9BTTIYm+1uCtA6/Sj7gUD6tMiOl8u8gH4i0Zi33FOQ2AwW92k5dDNIS3oJGI5xUks/eQrSb
qgyVQZeXDPsbUgWNMHqZiLT+Q3PIjeKz8a0sgKXiP//Hs8kv9gHzq1Yy1X1dnRQuTPF/JgXvjfDL
Aj1Wk0RmmdPO+T2F5XJ/GaPvu5Ns+g2hR6iW+pHFeD3Nn7iCp+KXN1o7WVqynpKo+w0OFgWIHtXy
ToVPbLzAje+JLs34dAs49HtOWLd5h/8H5IakSQp9QjZQEtBHl/g88Gbe951HXhbKbNXWN37DwfgS
+pbJfUYTdJCNJfe5mmzT1JcQKoHjwKk7EapU17yHEH1vImcP4KZUPm1Dhcx1ZlyAkwF7DDJvxgAz
Y9QzJw4Orl+uf+j83mqnWbPKqE7dVFFI152u4CXEFK2rtTLyWQHrZfCF27SCUFXpnwlnjBiZLOAc
BGhv97E3lp0bThJRJvNhiGqz6BkD9Dyf/XhWp5LuOmVEnrhm/uSHuA6PQZvsbb1VhWjV85fK2atG
SJsrdyAhoGttSGFfzasiQUZBU9/DAPxY0dH1B0R4/+Goir3xFRcLFMM1ZYXEY2yMLvtE+QuFKu1o
vt5xKxDsi87jvE59iHSR8Hc65eU2++/fAkj1N2Lv45jTZ+JLpsJ2M5HR2FCVrtE2rAMXAMpwZMle
QDynzkgVhasplhLowYaLoUo/cQxxJmTFgGDf6UZ5ZaQqFRTPih7gbGe/DqZfFFAMozrJ4QRckuyz
DKgJctGfX3mHwxl+cPgTweXbkyioLhBZ+biBt+TjUmk6+yTepgWRxDvUAB2WPgCGCPorzhg5xrru
qoqTYYGaW7+DHee42rt/odJfeqoyXPKo7GkBo0dKphccCS+KPkxeGb7eveqbfgu/VNO+5jEZjkVZ
M/4pg0t/cLKpQT52EzB+rlEG5W1a2qf1Q63Rcoohbic2iWsBNmRfEyrTCkMFK9elwZ25Ydxs/vmi
WS/KTqc94gw+yMTt9TNb4YyKEDtUVg15X1lTbLmV3ril4H8C1uIgiIsw8lz5ozR+K5LetrlKFXTT
JH14n4NmpHN+FrGjmniRYAAFEWsYiIh3kQvd6PmotwmiDkfx0Qheq6Dkr/W8KmeC/uOU3KM+xbnb
P++a4QfwqcAkSBrbbaMb0UH/g/V+0Mlh0IHMZ1QXAKl2C9MoKYlnaXMBqQAvXrKxLWle82Hjh7pn
ldHKVkvQBQ7BMvafkYj23frmJwKupSHPEAARTTVyAcZ2GBEakN6pfbLlDEiS9idYYnSU1ah42crL
VGQL+MIV/fBr1otgEVBMqinNIJTNnDiGQQqf88X6wMvyFT2aDwpnYiIWuIDhe8zH0HqQ3VyMQrgK
1L4l7uh3QVPQ+lVPToZ+dY65c9xb4PG1objzKcJPeLvUKumcq8Z6AlV2XwBU8n4Q/Vh3KWY0Bc+1
JJnHXJ9CdhIpXQqWf1BFt8fFFJY5G2SZOkoLJ4q6manLh8NqA25htHPXa8/1s0ZZ8kXpKy1qurXa
whxnmPNxpsSg5N44CXJ9b298smfBXkhQ2iciQ0GipSfyTXUY//cMiRPgKL9iM/mH3SzmQ8wKn4Oz
lSAJyQ4zr6XiTj7BFFUY6/bZOEcJ1XFh/CQyn0PwPWtRf6yvPakOk/iSBiXOOm8T0hhHokH3L7r3
zM0iLNtWLsHlpiX8EqCt8bLuCJprAP/tHmcRhAAUEp6/x5hP/5G0zbi7s5Ydap8Uzz1i3fVzSPOl
u7V+T9uHaW3UynkxAvh9O3C6GQS77bPx1xB5BYNPIeiX8mGcionwTY/jYft+TAUbLK0auxFEqRvg
VC1y27aAcusgJ5DLThIfKzvxEMiOWtD57hQw393CetLOYUyxlxfNXD4ZytZSanfJAFLfhtVuCbxY
rBpR4gpzTzXT3pBeJx+261LlXIjDQGcWFRgcAXIWaaa7az+FEVw5lZqpsGe+kPVj0NgwgGiEnOx0
CgjnOfsGZ3eqpEnlSR6G9EEp454x8KllwlXgtgv+h4YBtM/LXI8TISHLVRC80p7UfbFmmL0MbIyY
ILDiHsHyoam7EgLLYvQQ3p+hs3/LrSVcMae+TPBXBuhma+G5i5tNaHRxMGRjx+9xstH+NK80lrXD
/ntzDRleHQU5UEtb+4o1WqsteHVElebTUnaVxJVyIO5PwZN5K4XybGFRSUKHxs59IxXfvo9cXhJc
9rT4WiUgMUAW4CnfTypBA+8aOI41ID4vgjKIGw/bfY4oHZA1tvD8QpOZTNByIJEPSv643E+peP9Q
iQI+ShhMYUJhs592DZ8iHG6WWwK82eQPR+jLQf4ECswFn16aPLGT4a03Ms20YireQEb1eCDVXVQQ
1HYqR39K8ulLMtIKBrftLlLgEQbDeaplrvxSQaZRyi+YJK3OegTtTGSUgQpaKH3FXONWiM4AjIvE
nxa/Gfg63pwHAAhloPNMAWgrJo79UESTx/VfmSKBmZC49OID1YnqdJHl2FPl39pZAA/8ujkScYnh
yyEphrleOWU6e3KgpByHc/s9rLyIvYncKlKji28sQz8AEAqRSFVUk+QUFVB/XbvxxIv2i09ZRcqf
Byef98pKI9fbHqCjdBgXkK4NYHZ+hMg60LNEAJ6JnG1Mc294w9hrSRgaPCQpnHnYm7i7HRkZqEPc
Au/giHDg8ZQhY2Oi4+5wtkXnxUzFGWY+wUYJYoUEkBVflA7G4l9OK2mmxp24zhCUZLVp14LDuY00
NlQfnB1mih4AUwS1zbOc6lHSmDKdR4AxDnDeYRyU6J25Zwg6jNkPf2ivzFQ0BCS7j78bCGcvbsTw
aZUQ7XOmit/Ukp9FBYoTqemCZRmP9l7ACH7ExS0hFB/dbGLYWvdNeNsd53XcEYDbRyL25pO5/SYL
WBLnqH5KpK1PatHSlKALyhpfRjr2PfXbAVA/4IzEMNzt7Jsrt8p8YlSQjvhATuFoZkUl3yS/O8le
GfTzTP8TkxTnjcrKcwqEcPVzOYpzYDvifdlAhIYTdzn6Map/qHHnjGgN3iPqhJwIgC4WobWO5FiP
nmVJA2FLirtV4gGpUpAoVQ4GxHMR5KgCs0/hptNBQFBm3F2UV6AnqNoq4orx7SKv3lubO0w1aF3d
jBbriYJ5WFwkGjA7g/lklf3GHXEtI5p2sKucVqjOG5iP2nDgYmI4U2Z8KOmTuyYZE8cJEiU09v3R
kDokcmbkkr3x89+/lSnR3nsyqjWIW8lolItmlzNX2nOitUVXit1tNWK7MLe7uetCF7Aiuo5DbT8s
9KYd+RE64+LJttJ0pHBL2Uf8bWdws9/iWpZro84H5KWMoYd+yaivlkVXjZ54nEkORc3FPM0UmaEN
Gjr/MeA7hIeiD0//KjvjX5Eq9fMpa/WkbZg+/ze2VGf9Bp0DWK0tymqtSUCw10YTGYPCWg6otjEi
Y0PK4gRZOwzQ8vEnQ3JqGgpeJ7Ze2W0utK8pokX04GlBAnvDjUJT1cNda55040bDHGVtRTlAPlmD
TSY7zC0AI3EBcPO9KomH8FqkCb1kElBTRLB6SjPNfFNP15eHTCnoGQCHLMur5bpUFNlB99jNuoO8
j88UR/kxQmKpyJLhoP3c5WgtqNL8M7+B8eAW995rOxAgn4lto3MsFYdE7OgfHyMrfIKisvxTJgX2
dYJB3+JdWua7jBhXkbJ1GXBd0G2PG8m8mVGBizOTBfPiVrTdHMpTyAkybqNdT4noUr2gVO42R2hL
FxUx7qz4HX9hPEwg61xAONqMHXYzA9r6kPFl4EJrEx1TJao1n2yts1v/gm26lI5zzAAX5wKewHm0
dSV6MEDT9RctAK8GoINk17YzUn6gJ/ezSbQHqNTeXHN0gIKpSpnQ6LzKg+33IQ7vlG2uaJECnkZU
zs/pU8Fa2RvXehw8UgqeOcoRj49w3zln+irtU79oQsqrq8fysZEUlCqT8zGROQeOh7sW8FBCFMwX
A8xdqTSH0BIgwXDNvqD9RFP6H1zXeY8G/h++1rZRcPJ+4H+8+6gTj520kmw2EC+KVTvIu9/fwY1z
yOCqhtpKbS068lBdrh2SYl8Ihhu2mjKKJNv/rmwI2tkEIiQfZ/KYRX/s6+MbmvfNY+aCSa9qHByD
p42o3mGoT3YYeI7Ic97keioUMY5GelNSlrWSdbISbosbnX/VfnoAKunVuABgKu9uSE9iea1i9CU3
jxFCu3U5N6rEXcrcO4clNmvCPANmqv1qx4gfpEm8Jz3zSRY14R41FiY93LeP0a8WJ6xGX+fziOmY
pMKmN+TblY/v5h3nEmZOqcLBvufvNESF60pKXFrwRAG48XFNsbSLEBArbkJXlih9w898WGjp0k1r
/mdvvILi/N5u1Rd38NzOCHNOl3xefRsnn/WZlvU6gJqBb0Lw0KHUGBHI8iHVvWLnTxaG1q3zSTJB
WzdgTMZ7khj5yb0PxcZF+cb1ArHiFA38cSLp1+HHQP4GuIVjlaCuaVb6u85ntG8RYPLjgmrwh1wX
0LEHcbdgBt9qul5uJBL0P2bsyCh1hyJ578tRPJfd1Kpo4GGmrw27ylGeOWODFfe7cJrFR2UVP2UT
AMcwxSjDPC/cwfRqDQuTFky3XBNEzC7wlE8eJIkf/MT4SulkrkQHyDBB7wtjhTRT0aXK/Xw4VNYr
ztBdWty/CUE0nCPHyBE4Hlwvtugtydp/JH2a9D5mKU7dTqgNtVya7MKEYzVWPZIgSrv4sZwEz/8O
ykY1oVesjb0f23zTSr0Ubh1HM5/VCLxIeSye98pZ1HyjkOffr+fB8zLwL0TW3hI6S3xfn0zmu8VO
7oqRdbASrmCtGN8VY2TwI8hlCZ8qb8k8makRXJpicXa6P20fHauSSIOMg4InxnNc1gZ80QJ5juO5
XfELtxYQkFAYSPXhW2GlPA2wNfpzcCFZNRq61yphABp8CJ3Jc6xDv8cYRozEEFjpqVYgLf45FZI1
DnhHsewL862AhxUWA723cSDt6SmGJTAUIHzkTJQLVXvxoOUI7BLEpETEdheiwJTn+J36EF9/qHyI
1ZbGVN9O3mNo6OiZOuU9PbLNELbzdmscv2TWyYLwt+FSU5vDTQu0E1sD0lqguCtfpmY4GvY6zMlu
2tqMFlEndlk6bPc96luINbL+uG9BSpxpuct95adu/SNYMsKQr0Alco1tyE+8iSVueo1zcm1+BzVP
dGWLxFmYKNsF+yyaxId/xhCnuR7gqqMT7OMfjnXDE9s11+IykAJASU0MohwgZf/mJk5RzGZqfirV
YQc08PD2L+Pk2cS9y7jhObxEAngB6PWy5pcBJXYTC6g7DTjKfDuPWJYyvllqpFWswTWJ386MEByd
T20Sfef0hdo6hKONTWHWakPtJ69+iUMuQP28wzqg1LcWTfxAIUY8txJiEYNLwdSb8TcuGtt3F6Bk
XW5hnpSE2Qj7P2yGfspL+nn0dZK/xlZBOiXz60DEF5mR32ezq/ev5On+IBqIRbTpzVz9xe2ohKrE
9UGydQPzyyIvmFP82zsWpqi/oFVSxDFT2/Ky+RCSY+eNzsOz1XMwjQs5nK+86YA9ta0msPCHOnIQ
mwkL1P3PQlY6ieNzVTX1ZBiCXARfyP0Ft5Ven59yxi1PJFn08G6ZLqkkrVBOlvGIvpuLkjG8BYm+
ntokdql7CioYWmVoc4a0PE4W8PO7FFJ73zgK5pqGFkPx97POfcC5nAunOoH9Uooe1l+0Y4EI9BCt
qLlu58TR8KSVK8Inm2UqRrdzHMJvipfoIGxr5bh0LWotPZ/cDVU+/3abua3N/CoIDj1z8wr5xQWa
I0W7G8Z7/cmZpvbO0HPqnaaYyPSKQ8P4zA2IxiFG/KBLqwR3JWIkNwGqgkUDzL4yxwyPSqFMsW14
YH95S0eklbVXIgn4wZ711zhklqZ+6ZlHqWfX0YTLy8vhkHR5tmKD5cjT4773aVL+cgN1iMB2AB9Q
mhCZAtMzYHkElP24jt2NPtKDcGiuuvEwoYQpePjmWO/hrFcjhpC8v+SDyF3ANaCiaLZOZRHEkiCg
NbKi8gLUXdeukBsAGZLVJZBod7855CPfL+NQLgdsl0MbG7t/hvPd/VvA15s1Fqr1HjSTCKv7bbqB
JcmVe2s+NHiGgCHDNRi0BZCDGph0QlE3zgHhC7dhE/fWeqoeN9xVdesfAS0+7aqbU5h5UtfFyGE1
yt+2DmHiZ3FAZtk99+EmVCKzphQtqeZkCaNqxQNCGMEbrngvEuRspwCKktvd8KiX5Zik06//5Xsh
0iPMcYuSUbRKHiGJionYuwcqn8ugREcV53Q2sS1eaiw3rVxGHuiPTwRitqY7QyvRNyRB4pQl7tNQ
h1VtxqMv0hy6yFu3NGgtaHdN98c4/l6eLR3Gd97yZL7YJs98tw1ruk5riAXKbr7lSB+E8879tyr+
u2T/YRjakYenjPPTsx+md4WyKn2PdKvU2wwpyo7uQz2dl5zhPkhww/wNDxYBeqZcP3LHwiRzSez4
dm1Z07mWq4BbwHEnTsgtytvYXlIistgUlPACMo9wlxOaY/bMsEuVVpPmlo3jTAwzXJzKzPnxHEh4
zI1yhDpfnOWNkun9VKTPcMmT3negJGLUVX+ZXz7+ZBWZrDmsiZo9gpofd507jgO0QV/Frl5eivVb
2Ik5RaYp2ZgxQEgl4dkBw5egpASDWLOpz1R5sxJVwi3il+tM9Wt3s0fz4NtBqTKcsqPd7e4S2Ae9
jKHz69krcYVlg1aK29SZ+kqeI6lGxTtDjeIIE77yVNiqaf+2a/rh02LfySIL6HE5dO8OHKx18wtE
tEDJ0GEAk65GBRf4VsczcJr3oYWTWIyhpjENKwjJoqj/78YOB123yHifYhxfOhY/v/X7/ppdORW1
0W1RRGPpwRCVNM7+gkk6dpk5I1PjiiNyMQBiN2N9WSapSL7RyhngUpCzQI2kkVLaVptxGNZkKq6L
wuvoRc2+JO+71sgLAZ8j640LsG8DIutpDW+H1xk8sPxoCG9DD2KzBcVn2Lt5YhdQAPVhwPeseuwW
GBBu2xgeuVYK+p1DoTG5FsGh5hSOKhLENxlyXmjbYwG6LfRxGs6pL1Y7CqrfDEHUTXGeuzJH/AS7
MajeUz2FI49BhkPj0/ts+wmZCpvcmuY1gdZndeq+jlXweD0frNrn3y6K/muYdbIvac3cnsvSJh/k
mS/irtyBkMeoVggkH1FPjXcTY9F1reE951abjnBFcSXnvLSKX9EHa3lfBVLklnZVqoyj0YRGwz3r
+0xKQPfuLKUBp8PonWG72RJ1Tags6YsqohMc5jNMriyHYPuce2sKi/2wu11jwkzdQJIR1CvsLUXH
FFUK97qHER09CSF4viXL0F2iUWVyK+xS7ez0jLabdOfsV3JHm/EUGtj3zyMnhnGDmSy7MOMcpirS
3P8Mq54z41SWXOUvm57yLci3sv2meCWKLATQGe1Wz8YPi5xb49tTL1wPExAShYN3rMucikvTk+x6
vk41Uwn5ELIKWLwXPbbAlx5JCfS1pps3mCcHhI94ViS6Pqhp3VOtQomm1jB9dn2OyniOuwK/DDOa
cgbg6Xu84c/fP4hCtvE0p5VkXzEAeF6NS82m5nVlGbxbBfrGZeI1J27fgLlCiz6GijZFd59j1Lb7
D3xcV/ONRObT8qejKTIj/JEjDsDWOAuCmeKpn5hgGb/JcrDUdsDv59vN4Jet8zw7vRhf6mm48YXO
WZ6pYMD8rjyEwH65Ry9x27T2ji7kEUMxkmZO5ZvfwznV37AiSS44cpCHm7qMMjf29WNLH8KNh/wr
j9Hbt6J6GuePm+GncA+9MB/IvHGrQQJc8aoZ02CqoRT12o15R7sMuqzOAgNcfarrDt5z0rWE5DYd
6VMj4tVu4zhTAC6sG/w2CQ13A066RuHDwvbP5RU5EGtyw7ZEYjkuGv1BZkI8oLExrIUfklYRjG9r
U7kXRUjr+u0EwOxtXJeg5+3YUEa50KrsI52VK7EIcqOPlPD5wjfAr88uQkhrn7+csmwo4Z96qMzP
4Kor9cn0Kt2UR8C8tnbAiWvaUvLSipbrIJLnDLcanyfgDZEbP9NKsNrk4wOOUNIprE+ObHYfzHUP
tXVZ1cRpfGrRzXJrrYWj3jkH7mUBWP3tWdPla47CBcLkWPkZoRnFYZsng8ZVqk8zZc6tm1a9fitT
u91Fnot4IGFPZMhviHbyvedpxH3EeLk+jEgAFj2f+rKYMSeQyIJOYTMprXkyejnMe8W5R/Itt3/1
ErLm3Eh+vOiP4VO2qRrYsMsgeLU7EsRNU9rznlV3MIw6OBpDK4zBLCAp5CzDp5ARWCTHj9woYr8r
lMVXlBgR41aMWr5hGwK37TaGyoY+BpGL3JXcvj5kTiZC64txKPuf7cNze0NOMjaGKW+yAUe1tXj/
GRriY0N3qrlVYhYjLvebDB6em6g0CPZWuOhi1DjhTrUdmRmPXj7R8+6UXW8L1h0w2m2y61cYb4t2
YJIGo3hMLwDI0gha0/rW5rM2mMomXiLeIHVLLK7Gl9U7jeJeq+jfCKnNELdN7WU123mTYnFr08td
3g3Nsnyu1u/IOjU303hQa1fQJbVx2eihhJ5L7KgaUWGuDdBQ2yUXAheXMlkPNcgNqrbJavR7bVQ0
oMwmgeDOctNvA+Tx07TQSXVm38f57gNnzZeBXbNQ4EbsYLyw+Ykg1BJOAZdQCnWcRVIVmN4MVPfV
D03XXz+Csi70Ud+nxFMZj/D2QeREknoOlY1Na0DMKQN8opsX6VtOYsMH7CzOzZUYlCdMAFrW3j6T
ZnVtGi0aFm8G6cmQ6UXKoVsbOWjrbaZYH5ogcT0GI5SCyExP8MVdQCEBYpgaZlFoDCitRtIYBPmF
NSKAy4C4a84GMykbn7Yjifb/0C70BVLg7iLHM7QB/8c2mYUayAa8KQN0k15vHYxVqgHmDeYq4x6T
TUYS3d0vifnAOejDzWl6VT8Vgftl6cCEVrX7XaH6UrRJush+1k76HwavjLn26ODLTlMVD1LFNM6C
L+Enc9rCVbW/1COZ7prPUbeF2LsnkI/oj2RJOS2OYtuXVREG8dMzuAsreqNGxuUi3VsejmNx8qnP
oCilL+NCQk3i2E5MkWdtj1tiho2H9+yZmIL+Yt8CinPL5pZoBEA1y9orHM5wB9OyMHtgWVfu9QKL
PVsOJil6IBVpMJ/9raR6mLKWCK+UAK7lQCeOKVAyRrJiOkkw2B5kgWmbLovO6/1JyLje/5r5xkNz
vlfRJDWJMgrZObBh+aXncLmjrvmsAGMKLEnZ+2WjKGlPnO38qze7Yq1e5Xd9xOh99P0Bd02etbZY
45VG/KRcvCRnr3wY4HvBw8KDbZNxPLdvA5IIZHaG0xl2MAKtM5KO5PulrmhMpPcr0Qwlgrru/ljY
Z5lkbrom5HUpq/+v0eYsXOcvfKdw9UCf98impsU5762iRdEf4amv3TkjfsZpjnmbimzpDqGhC5+2
WwOlZBz8ZmFFOxbc/Wc/bbnDxilpWURjjNPUGFscOnS+EfT6Iel18pyC+sLEfGa00tDtc+kMTkaS
kiUbMuGRQgiHpSmk6Yxlpi6poF42Cg3DrUQcdixWY31P517Jb/tKDkwAaBq2qi9Cw68evhoa4XJb
VKot08LnSDl7AyB8rYqXtMddScSEJjwfoGGgtZ5XIpkYrYyq5a6l67ORJy9fdg8/328EGoOfjDvf
04xrI8Y7IBBaUO60GivLKRgHUEpFxEP2jCTJo1t/SxUONaL9ZFyc84pGO/5AU1u6ziW8uDmZIEAX
Sg7btc1fbLcUz0OPSObcAHn4xrKSQs+111MzXUT1zONwVq7Ysdpl1dmFJTZsWl2ciHoBDO1MEnO/
+7Yy4t6pMdKllvJ5bU7OT+sKr2qYQW+auaTVGwkkGi9jx7tdGcXzCz46z77TQ5cyY/A7YFNQIm6l
o+cEv5bXA+5n1d+zloZFDr2zmP8mhSW7Q4FJd/wyVvZsS8BpxkPGK7eg/FVGVxZTEzaB7CFkqnip
aHP/wIxehp3N9MmJjpVb8IoEwwXB+Y6KphnvhzL+6+o2QFyP8o7aTNyfnPMPKL8XoyI+tW95JXOn
V5Jd/iNacFvKd39vHCU9R9mykqO9kaiV8S+esPYQFXR5uX2ZyLPI7ZDBFJWseS1xz56IhDC/Ahpv
WLzZAR06WL9qiDKUR4wbxHl0QvcSYc6XFElGw01LYw2xrPTB1Z5BSarQyJPiCeMH7dgeeHCZ9Uxe
gAoo6IwC+MVkikzhzcHgGaqp4U5XNvQSc97n7kFMCGc4J8ZVvIk0Q0Z+jIU3gyrJsh4uGLzGS68G
CyyoPyIXcxQl1X4+bj8EdiGf3Y6SbTP1ktBWBZPLLJ8kZROo0lqhOrEz8aCUDSoySHMGtlzIb7Lc
3vWTFMDeln6U40nDn6FiKLtP9U71RxruihGm3wB9U+ayFZ1+HA3VhIHghGWiV7QkUTcckXE2J+gW
pfGXa3uY5Eamha8cNpXelb6E23cnMD0iVtL2mG6gkL/Lo4J/EEmIPUK2OvMh0xwnrVELQHSqVDn1
BTfeoL4sRDu19JSq6IYu6+QpTxrw7PCTcBoQWrszd89JFPk+GHZYNhFwY0HFvKH0CW6MusKaN1Yr
b8TOZb0gHjRWODclxSnYpRX2fQqbAR5fZH+u9AVLttHHUu1K/EBWhYp/uZbS3mUXqpffLYDVnqg7
GUxO7UQ52mxPa4VntvvZkAd4jupGz/vZ1leikjgHyE1i9mtMlXBa7ckRaFcAN3Uxd9nWvaBPPwol
asbLIU7pVpSkdg4OucAORWMBC/ilxqkg2spWq/uzKS/4vKiqfTBbDXLfTmdH2uEgSaiT78JLe5oa
1M/X7i3I19wmaiPp98rvqrGXJ45Kl+O9NTvO7VK6vrghhWzEAoFtVIy1G+mRdeUfR9gzhsFg0hp4
i+/EBzaIC+F/D0KTwnLZ1Y2LuLYa9IVx2iEmPQRX7oeHEwo2kBBGUJXPltKsbQsermAdaurDWsH6
v0hGIZnU50/vwZ4VRKmpN2xpQnyhw/qXLIIXneQL72pcQM0imuV4gv6HN4dC79N97dHzLFO7xGRl
eIFAm8oEsj0EJSfNAGvfXvtJ8vzXDL5EjI0y6U9GZVU5YNIGDP0L70RwicyIcCr6FUMmp8CZMx7p
RQAR6EaLUOX1mAwVkRUgH3/k75a3su7JMu4qc8/VC2OAbs2npZAG/A8J+7MJzoYAkmAg+7bMB69t
WDRHdXDsaRsI1MzH4sE+ZFXbmiRYO+hNQ2CEQcktAv2g4HJ3eVlsybDiB1wq+HNckA2YbJgHhHOk
d6Gvup3DqbUOnUIQL2EZHKF2ZWuKZNxam+Xoi30CyhJ66IebqyVHcYRRU3JueapE5GfuMBwKglUU
RSLWwobaOXi045LZrrAIunnG5nA3MrJHcR6YyEUv4fe89UA0JcgueKpZpNfrlnlb/ChO7H/Okewy
np7v/ZSMGMf66KgiKFJwPrG48muZs9eHLlUhJYvHdygC2K8jiIn2GP3L1hpFrPE6FQwWYCUMr3uh
0PPcCOMGfuSA/376tOx0hW/jif2bQdPR4JeQAzlsdB2szDiGN8fnsUUuUexxcyv4ZUg+iQkPZpGV
BYeoKDclkLxnOSYA6cqONE4VlHT4gKn01wzw7XZotDhqEbw3NGcJkuiyM8aauu+tS106atHVNBit
C671ASba5LwOVS9EzVn4rU1FS+1FHXzfrLoIkCE1q3TNC/imYVs5gSt9a299U9m6FzWM/7u9kCwh
KeG1OrkykKPSxxx5bzKcsOlpH6BFaajNsq2Hbt0l61iDlI8iYNaI0sjuJUAkyr5RaDc0qv2mbmIW
ZswOQFkoT/cOt+vd9FEFWJSkNBMtwekpOO8KVr94ZPsDPMkNDPhjY28c8joHaTEBiN2d+X1IAfhL
AcmRweVUjWVSlLeFTr6I4mvh23jwVBWwrZ3r+BEFwm8EaEBii7XjJC+upS/VQr86VyenD+9SzS6y
03d5DtVdN313tKBNws2tZiWmVM4bjZ3ARVK0tfXpfD1j9/CCw/Jy7P6dDwGxl98+mO5ihMcVvlfN
p1lPjzZGF0LGdsTZxU/1NOSSefQovN5xmD0ikmiuh49bgpyuYj0U7DLRpjc08ioC5z4K3wdzEmXu
p2WP2D2zXv9IA/H/h8LxlzZvvxXpbedNlIXoL8K4+e/ZCt8b9tgqU0Xc3S4q+5JmbzyxOIyV1GDS
cnRyRH2Nh54Kcdi/StwKEW0LSu22OEy6p6hT71mX81gd86wqMHBtRyaWwtz6W+qwt3HbTjkBIc/u
v+0Z34U5cwgLyDJlrSGha+ZCuhbbID9LBlSuh8jjcsT3iP0g2iKTqStgTQtuYzs82KfACGnCW1ET
pu9pszGHdtgPHNwSO8cTqxqPLAPqrI7nFCiLuj4o07/tZWC1vRw9jR8SlKsdzkhXM3671h8rTzH2
X9Mmz0quSjdCcAmFtAEmY5goQ2N/iXFAvrC6SrXrnZDic7EKXh6amVmBLf4Wn6E4iTOASuKiFtql
tB4BeK9pqGg91W5gsT04tosDYd9HbgwKCEdVlW4k6gEg1LiPY+1PDRVdS5HU1TxWRstoi1wlwVUW
IcKV2SZGgnP3n7w4VTj3zDPJhQn6VwDDcF/4oLbBh1K7ODf5MhoMwmX/ZXQdBzcP88v3v+howPj0
ZR4l6miUeQzDrrWEwBFciaaOtUEUqBZnZfMEH/ZR2+4j5rkMpgxUULn371vv/8T2biBG1hLJvFMP
ABpuCYBs/rI+iSIkk23iA2QiC/Uu1UCx9IEBcW8jRK4/m2uu/Q1PgdtTftfrS6cPa4zTZKKDhJza
EM7d09hZOJE56QpzBsipKjI4jGjWPkjVZQhOeCHDHbeBAc5aJ4ISaTGbS0UTNtyoaC3zLdfazHee
0k+15y+kuR47vK4r9VDCbBlmv7wB3Kp31MnhDcVTxkVa1BHxmu/+/i9tIqHT+M2jakgItwWIuh5u
LsFFPAmJmTBfOTueMOknjYpJp1dhulMkiq4ri9EpLsluzG2NYc7gvcwhabbjGKMS1rE7LWUfQ68O
5t3T5wIMLeha+mMurzlJVt4eyRFAgGGpD/8YRcQ7AAwAofGi55RmEHtQpSvK2lulILR6xacAxl7C
WoIpIalAmV4+lrkpm1Ix8DztGaDaR4mFL2FaNnSsLSKF4JVcLt7SZa8paIIwRynMRzXsfzeismla
eDFW65nDZllXyRU+n2LHEpmaQfJB2Q9QwM0W+0rom/ToQRxVie1P9/rRll2tayE+vSOzuoBhP5b3
bMbOcwO6C0foWMd8y9LQez06uAow8FxZFEU3BnHDDeZQolLqRj2Vr0MPuBXwh/EzXiJ6/kNDbw5D
GJratuqbewvtO/T0fXGWJRXAxYIZaEC6CckTD3tNoRthprYqp5QS3nDFFrzX/YsytZM/fFMiNlQ1
i89If/LfXaOtiE9BxE35Dzl3Wpwmqwva4Uf0f3mpO/1WK5fjbgu6WFGSwxE8wNKHU556C54Lx5It
iHIyXO4N4rPKgM0Jo9/X2SHu26ULJC+DKkCrG1u9gKCJzNWG+K8oeOA8ZJzkVluCYWITWYXMiXbV
+iqtq8oSMfmbZwtoH8i6Bo4SwpEryuseV4Hpk4XjVotmykTUMQsaklk8yXbNcHBbHQKaH6jJGABy
DS/T94lACaIkDVdCkgA5RGHMrNvx0CS/DJhQKnbqtWHyqDjADj9lXeM44FR7RFCowL6IlyR6fk1a
koXidcnEPNJkTdR5YeSRISrQ8qgxIW6xEpdVItVYxupea87lQUPL3rhdYhOMztjQL8zj9aB9XW41
LfoLeLltECxpZM0jfkvnOXRZii/sqZ4KJX2aLIWdndLPSUsCq6qQ2VPwix0XXsPx59mU8y30jp3l
Je6aTlW48HvUQ6ugS+3X7VXPWLYKnX7eOCytwJT3Qaw5OcwO3iu6++606HuaKRU4XWLtthTamKTQ
Rtq4hdrLl6Fnm/utZp8pNyfQvVWNWKDrPjd2nVdSuX48861KGbMX49wDe+U9as85ijmW68aCzYK1
eavR3YANWkfnegdjieXf/ndakDPCaObHPN04xJ3dZAdeQ8vQUzrcUAHhhQ9SMN+DD63jEevcc7dz
hsx1oiHJYF2MRxgJ3b4n532o06aC1y4CN1ycoKIzMTGqWBy50GVOhikUhSpaaBTUM3p7X0Om6wD+
41fbGFt6g/5QeJyKqCi9xXwlQM5/r2j1TqsLvvHaT3xgYQlGclCjmNzxcl0949LDEz85eCYYBG3g
OM3zisaFEJLUwgMa1fE2chfdiVwn/lIPAvrYvBjK+eUlOLw9FgJ1cMEwvFuVJrDBwUFCus1kzHmh
ecsfC1tsy2OfGtw/s9NyqmkGrdZCPILtRVPRUSAdCJaS5MLwclWPovfJ+/ceMFjk+MC/14jbhAz+
LSeu8UBMdGRn7xRqcaWAp4Y5GC/u38T7KCHU2U841tsLbfHZruTx5eJBV8wlQExaSFCFgV54/yZc
foygikqPnbfai4OJ3QkyKbvGC4f4q5sh5GDZuzD57xNcHFKb18nJyKGTh/zecQhOGLqnC2brwNsG
XvvIQDb20IVFhRJTV1iFlxcqLA50wFgvB+Sb0LdB90WfWQczlPsh/Dth9Zf9zjn6MJiwVBLIYNac
JUX5hlN2MKwSI+Zds8RkVG2fDh2Lp1ReoLWMpiucN+5/xvJebJ84O3tygAEE5tUp8uLnaYAI5h5x
Bgn67eg7wf7zZS/EHAcSnYeC0c9Pkpe3EWTMS2bkvCrVCxznPz/uMh8UcB+cVhZmjjPlsCGaubPr
iG/pGYnWqEpmr+W7rI+LkD4ZYGKHh2GdWEHeKhbWsY2DP/C7APN09Pnkb2Msho2/4M+n2XgnFqEh
XQyqaZbqx+lQBMO7I37zGLMb+9KoXMaB6e1jglFL5s5UI1ns7Lrh4gxyydc6VUYEHv5BDMzH8XSf
Me/XyMkGbi2p/LzFvmd428WMG3LPqHG3T+I2awk10pB72OCsU1IwPcH4kWc61bNOUYVrd0oAKJ+0
pC3qdaSdT9BivE2siXnSaN8Qypk9xO24s3q8NXPUEL/oRnMuaHwT2AtD5O9iwNd2pOallsof/a9E
nHdQZKT9MRba6KQVTFvbdM0Of3tp5+qzFGssi1SAB4HOsle9RGB1c6Yokty+0IqoCUFuFnm7PQqw
e7SMOmXgZIP18QULjxolMLHgx6+8v8XKW2qMqDxsted1wohyjhSxVBWNBwdl0CgLjCiExaUkpjOm
pY1Yjqtni+fQIULHA6VKjRnIch0iwoZuVwX/q1BA0HhcPM06Ml6aVwhJsCdH8vfxEJu2G3dR1yrV
f3KN1X+e7SzKINSK+WzBbIzhzJNq+HbnESF5G2PgJKdxO0M+OPHiLjQ4EHvkpuzkkPEmttW6TCIq
h4M/SjksfecK8Zee+jGMl1CbYXEstZ856mW1aLPqWaetGGx3uHdH+zx6jjqcprbGZq6P2QFJIPqY
vgsmZdaiV4UdvWP5n/0bFFYDe0ZVdeBZCUiy19yLlRFFXzxKzliKP5B9EzmJd3VHnl17GkzUgFu1
dHTdTwE5sfhOesbSlS+jq6P2O+OKO7F8+ibQyzbBgHPme13Dt/ydVZyFp6B6ktgUFWcn0RImL1dQ
pbS6yEmWCVZN6tgjbk8JD14kp9U4APYoMFao3+WcYRHG9PrPlsSxJ8gdYMdSSCw/rKLq+HsfSUw9
zNt4MVqyoN5BJ8/G3e8FNgeHZ/QVE9vCyGdWfo86duLq0uzEWqhnXFX4mDFnL/1BElGmW4aLdStU
1FwcJT4YQFNcKfMBcu+qX0hlf9682Pru7Rvui2Lv5AS6VCHl6faupF1MaxEkfPSeskFmJiomkEMl
thv2ETiyhsCCpFlst9GPAlH3bibUZcomHC+Lp5OzQrBHthrWipmKRzFznDH2dnKdMRNvlyYBAV/q
YtytNCyHwDgHUsfQMRA0aT6zqiNydoOukTeGusqdLAUCbW0qQyd4X8oIp5knDu0nytha/5HF2NR8
o7Y4O3vFwGiigS2UNHvAsW+3m9QiBdeaHs42qBAU5zJrIrAyLrMwewlPHSHGVV3d/b2ju8vjMdWE
42JrOQycZYf98MW2A9VWV2n9f804uuXhLnaHzaw/4hI+99L8Lr6t8Nn6Z9VhlDHwV4qUIC99gKZl
Ib0XOda3yDL02jcSdyCxdbEKuzCLiUayZKFg1i6bZC9BbecjIzYDsYbPLmGPBz67vl7JLBTUgJxw
E9u7+Ud4qPKeg64QSCga9Nw5ZUTfTDoFNN+OEgXioq4VEXT8vMKD19/jJ3SxEXlStFm5aM6Oh6O0
6FxB4cMQZi8ymuJZHz227nrsi/EW9zHetOlNnFcEygmiaveTcj7TWwPFsTIv02Ks9vCofFxDABcX
JqL9aPXHXgKUl8mIySGJFEKlzVzjlgNQkC5AZcY5vbRs5IETUUNw8hr9+N1ISqZr3RbFlQEY0sv9
XbIS+V2IiStdtRV+08NsJjNL6mXNyXS9p0vgCSh6XOkOrHIIGYzjIUhA6NklyjRGSyn+Y7B1FJb3
xafyZ8rDRTs7GPkF743AA6UVW/xHQcKKlA4Uwdq4fOredkMRdMMb1n9fXG2N+O5a0kNUtjLHq+FD
xfW/Ep94zyhkT1t2U34nVf3tjj+2CU2maHBocRpYdjuaeG5gGkSqMvziZqtp9YH2pcHrXSHXqlZr
6W8o9c849oE08Od6t+CHrO+5m83XJBEiGgYk+qA7GHHyRmrn3BhuAHHtMBfJcQolyKUE/U38I1s0
HkXEVTsQP1AtYRr9Cw/nSz+pMoW3GAlTWroli9gJWGiJ6x9R/19zRhhn3cq6nw9FpQ7fQJZwKb5J
GgnXJtk0lyc+md2+1LBtEtLffBkqBX0kF7sLhlXwEsp0xEIGShr1dNcEcxKesCDs6wX1jG1WzJTe
kXZKNqo/JecT9/u7gkoF1q/GvgNoU0BqHiCBDqZMWKr6JXs7FO0xymAVL/wQ7MGV1WuY6ARGl4Pz
FMKprLJio7AspxsXdEUaeXDlOoVZNT3NV1RytCD/s9HqjEg43Wmev9CRV0gg7QKZJ4ntfN7VeZBf
SNZc30e+eBdWOgENb2stKwvm7JHrYaXO3WXiVI3XeFCqg+WP6+oC9Cih1yPmtkPz8JEBuf2hqfvE
dnWtzFbJoUG/POgwnjhKx2qDlAXOm+CQqEMs8V9mAglTSKJCWb6m0gG100AonAdQV+DjdRJItRL1
8JnUaBAqUgQO0HYTlUqEwFEy5i93goKCTqDFSAyjd6xhKbNLvcrwBBV74IPtEVG2jwkX+prjM4FM
YpwiUILOtZ9ipT1MrLt+xQLk/MFhoRqLgieGbShEhS38ke+aRN/a8H24D+B/0AjEsbArl1ibPWHr
iOJEIx0s7AMIYXJXFPsvnefODbE+8A/dTsKWQkKGx6E4KIzvS1OCF4gxPl3alhdOOGaJV6U5FHPs
lvdgvDYvXLrLIQTAPk53+tR7qKDxbJc9/EilHjtBmMOu1dRx4LWsT8MK5xT+6vIk7YA/t4c/fEjw
d6U9b3kZ7TeXhuOe3V1tbJPce5dTWjeJnVdnGQFiDBAVGOP/WOyopf3i3qDfKz9VAoxzQ4b9GOsB
SRhICaYQfMbB3NxykCqBUjv8XEfKGqxrhDmCnkB4zsbOS+735Lb7A6830IBot6kwQ8CBNuK0EXIj
EDdPoQ4T3Iy7RoNI8jS5S57/G5DiJ2rahg8sZkCso/9bCp35Cwq3UYC826fCcpu9LxY6pKwkmaMo
XWamyuKasXAAzPLauixZu1gBrBBtq5ZQ9q9lMqtLXq24AD544bEeMxMcTMXdaizY60zSd/bK2CJR
ac3gCCmprvUBksNLMCB1M4G67icW/G2N65N5DUQACWgs1mAwl5NRnkU5b/R0qRB9M0B7bmcgWD4H
+1n2hr/anr0q0X3r45K1g3ixxfpe/h/MdHl79IgVRRUlXFCH4cMsCfjIkSs33s/Ny1vDbCgW1pY9
JOl+BxP2gCwVbuRz8LhVE3m8TFTNkYKm/dnltJHpgncZxU9ycylnOnE7IrXQ5hq0fPifQm1y7TrK
TlWWGmTBL9ydP0dngfLWAafAqF3jfxUPK6q7+OzbFNkXgdd/AnDE38nGlEzegSLq22HyIhs9ACdG
okqM7vi5pZ82A1ICPTtCucy8tZGJxtIj+epD4hSpv4OZRRufjObdc2pNu44fPgbwXi1oAqiPkEwL
EfLNs2+qdaeJxmpSK8vzdDty2NHlb3uVHPmCpsRZyXQw4TWW1P3s5IU+0dqWgVqrz6LpEzxhs11r
2cXjD1HceQJo67U1j9YL3UxXss81RRNKx5qxO3mmMKu8wJsXgYNAs5mnTsFOLsEKjn+0MAQtswbn
lSO6p+SF88ovr6U/GoDFDVaMFYFiOSdSB43kXeIIQz9yx1CBAdCYLvjWdVDxob7+hyuAEUQTA1ik
OD/iHgJxv3TozlePAbtWT6Vm0X3YIfn0MjBFB/jQcLVBL4naEPwumiHEzCaXvmHwFAHfbjP+9wQb
4mwsg1M5jueqXzcqYz6FOXUc732gLCbUEMrxjbQnyH0W2epRERXSfDDb7BtABJGi36ctjH/8VlCU
72HTBzD7MLR7vh+B7dJHMbqPxcKi6pcJuAFOedfRoI9DCAVCclcwjOYxKXL/fX6OA7hPYy2k5hf6
oqh1Iwno/lj+SyW+MCjqnnrcl4Zh/4A7V8JB1BD2C6OQIqmqblpgWBtb6eS+/7RZ4CwDinxOmQvk
zuyFbnwK+k3PtowsseJ6Y29fkcNxnQkOYwyCBMpoABKKrrt5phv2naO6gBYW1942hU0a1yTJ2EK/
7ZOwth0g+Pl4p57lJ+woyxWumI7JcGeb0dnnJxQFXmus2Q0emkDUmXOzL98uqdS+InB8VbYynq7T
4BjPoPB8GdwnSVfrcRZV68YyY8NHVthKB8k8p7b7PWbnW3LzZ7YX6cLpm9ChS/VIBxjkxQmG7bfW
oGcNa4TOgAUkhFUpa67dZTjVXekHiSH17qd56uy+8qY2ZaQKoLjj7hcn3MA5mnqT/7Uu/IrNs6qE
jefeK03DC4VJEYebstUkIrkDLhkmRsE2qNveG/L4lCX+JPkTIEd5k9d5CBeeOSUcRvjINVjwz3vN
r4cpZG7iFQZTk5bMVH7cP41BLmBC9ErorApLBVsDai1AeJspvhiTNM6vrZfSbO141ju93JEhnuwY
hLEF/fU6bKI3a4n/IB6P86EUA3hl4OQ+Qq8Ljz5b2CBlnfurPP0UAnnDabdqyGx3/1Dz7qg/HU5g
sXN7d7f+fryUaHAgtNBDDJ9T9eSl8Mcs0pqUAETGPsSIwQ0b1EiQwTUsADHfz/mqQPoxqbt4inad
LgT7cizok5ysLg5I8iTpdg+T7dTj2nfd/fa843AVdyOgE4fnBziAl9aqng3+8soURTgrMJxXNTQn
i1b6d/U3DEhrtv16oZstGfr6OE1PnvykszqLLWfu0UZYLY3SMoSO3BzSDeNj7+YeECOkxUYD3KmF
GWwT6WVsifNmBDVJ4O39Hg/zqISXt0XawqQweitGTcpA0Ng2YTMnDhQYhjzTP09oVHWWVnNEgg3F
pWyA8hUOvNtX2HzN6sqIkxb7dED3Y2v79jOuY+WQgfRI0nSxIv/ASOXkr9XiVy4W6ahWz/y9/PE5
5QqxdUPbhcXuCmrsnofZX97K6nzqTMj68mb7q/+JIjAHfOxNYSCje+9Xo/Q/9SxAtJ4fRjvBOJSH
h35yPHD45Bn6+b3ws13WJTNJEJB1PdQk2GnUs4HXIQFrwXlc4cRlYaU41X5hknudOOuWF9gvu0bP
yFLgS6VfhkoT7czAJVLzUpqiPWzW4v86GUt5/l496qNGWsoLhmS7EmQc6/1mlksv4mS57N75wrb3
Z9l8FbFV0MVkdWfw+T35IW6UDWCjxsXN4p6I2C3CFPF/a7rTwco9ayt6wDcpSlyiltdsoKFk8OpX
oxDsNiGR93/7j815l4hdFl+yL7Nk8deM4U6FnoMVqIWHsCjvHZ3shJpaN/gNaCPHbkJQm2papQx4
qHSDTWAyVjCVroaeh3nuGu3ejYQreA4IWyAXZM2zVrf5DKbK7qNzntawvLqGfjyQlgBDhPwiybMK
qnwhjP6CAskshlMzsFzv0a2krVLrf+PrgfNCLolmA2B61McarFKoxUKK4cNAIhiM+6zWL+1QaIiM
0N4v8MpPUtXztwepj2PC8N0Q6yGJY6CBhalOix1nsQJ5JeH7SvHWvgWQuyuq5szYQ0i2P1vdgb39
fVDd9mMupmog2RwSU6F+rO8SgJyz0vlKA12NVzlfDTJRKPTOK2jp2kKTmsg4Po2XIEND8O+8i0NL
OvkQdCAhcrABEg6Iq/GbAo8pMHLYzpq0joylnaZNoW6/M8zbNrGYKTmw+uZhYMU1W0qQW/K2VRba
uTMpq8ln0Dpx1zCWCXm8oRfFU2xH/jZuyFvOHqN3+JAlJ7jKEuGk9uAJXVoKyNodUkt+1fZtKRV2
zf7ArA6t9ppQ4O3lsIO+aUDZkjsKI7u6yrEBu3vzBk7DQfc2HnQK/IlT/pT0mu5i2WAyse91diOP
npGtBIWENndjBbKeVJS//A4tur2rETSkiGVIwjHp32SzZG0jz8+aSFAhtglgIQ8LG8UzPYLkMywk
nzY48AHEZfE6VLaVtKKywUriF6piielVN158zzH7IZS3Blv3LenMNlCu2DSzqDDd0zX16WfCddlP
rkqzjYp7pBwzsu6VF2bRPJ2WnrPpkMM/sTWIxaKg9ZcUV/cVD8Kvhs0WJZE36OZALm4oz+aTlWl0
Z4rm3f2gWSsfvjhaBFxejs9bekTkLfeenlN360W2pUT0LiF8KXVH2kIyJ9RbEhVCY+S34oNZ4Uqx
yUP96GmsmzvZD8jEObJfrfsYLq2mtAE7vcGikZdXJXtWf8PgNBAukWbyo8XFF3m7gaD/zE4b8fxN
YOuMF/QRCyB299Nia2EFYDL4yK7Lxwrr4nDsWkDpfAzO4ZeqM+xbZqBisdcYwtV2lzC4uW04ou0b
kVMb1/mio+zmJmEcD7FUeU8VQx2C4aHiqG3R5fjoimG1tMJqSveBMwpney+LB8e7cxRgRi2mmcCJ
1SmPKkesxOMuIbdwBc2aohLp2KauLH4lDmdH80qN39Cd+oDdyos1g/aD5UJPU2af2kDKIPNZ5Pfk
SnRAmaebm3DcPUEquJspBa6e6KWDCee4hsKM3jjLlD9lJDfTY47slis144VnrsvD9nDskQ8QrxRw
7Q3LHnyks1RNx2moJN4tqOKxCGgxEzifU2/kRn8E6v4UpmpfJhEogACf/RiAqEEbzznn0k6SgsSY
ma0mI8V9U2YfC4tp8A6jc2P4FSwg0yRmD+bZ0Buaqu+4vR6bZs5+r1pAT48uttfvXfMNGpggiNjb
+VYy4n/pBkRUuNsN+/Be6W/C4A0uoQRheHZPGU6nvNCDW4ZbkBN4KpkZGALVABsl39uMYTRX1nor
9wRN/y9Zc9mPZCiCzDzvnOenBkjHbxKzrwKov6xvsTcz8vKBPOsGnYwPySxX04iQjErDAJ1Cmpqu
hNCZshjNOS0pM3tVzKQTeNs8N7ygEiP93wCpNB6e7kE6OG7KCatWvTfsvP8NihmbmVsQt6K/LFfQ
5QU9nVAy40aIsHqyIlyr+fh5ovRDxv/0hxdDEWgqQGbxcThXjVxAXy03Jts+LfT6JnrgWbYWUEHz
9OX2EZvZXdlF8djHA374VpSePENUnd2IlTpqezWzJwWSSH+Eg6YZ135ptiIrl/YBAwwcZB1eBXzn
OgVjQrtBqH6y/VL6n9TwqGsQwZ0dqKP/QPav/b5WPQqK5Rr1FbOpgTE/VJW7K7VP2WhFl4fluLSE
SANrlJ5KZjFYUjITy8rLpJ62uOh2R2ZTwDZK2uI/ECgj0m5TAIjNIwG9ggUax/LdlN9u+he5YQ+h
yNMIgiIA8gTvOJSqGS3sLFQR1hCz6wnRxi4gc4TcK13r8QVJMh1wrc9DryQHlWgA3+7gsRL/mJzC
BWhSXD/v9S0j8i8TQE2uSP2yUsg37FZeqnIWL34r5o0gwhFU+nDBqXc2VAw0IOkaqq+KVkehxS6o
zfCt/4zPHIaoUGPwE0YZly/KijxE0KMQORlc5JEbgu7bUFRobuW1lr7hz3X16AIIh96CejlB2Gal
H7H6BcgDK0qFsMuefkR4+3me9AsGnOL19KO7P5LzNre/svS0r50dS92Tse66f4G3hFSi3fU5ey0r
iCEnYUls5TtDmmPEfvpftJ5QjbU2w6ILB0P9daR6Nc1RM0uCs5PcJwpVFZSAbFW1DHXEw/KXnMdu
DTAGQhBdsDmExgG3m0bKdzcDdq8na1//BJqenKFDIQBHnhZsrKecbbEPJf1fyYOiTtFIi5zrviQa
FtU/kInyWgK2AiMQNbbXKBG/rS0TuzaxypnCqGoLKsGbX3ByAZDAeb/CLzGiwWvwKtn6qax0VjbM
VCjBjDsfgDF9NCg3lofIoot1ITf8fv1R9IbcWyv/7W6wcLXXeH2/0gu+DP0ufqaqJKS3AmXarjpx
ACP0SaWrv2qVmiJHWWaaGe+iBYOXQfCoP6ZT3weodLimIP6QIB0SrA3Gl6PrWlff086LTo83oFQz
Z/toTZnyv0biFwyULe7K+HdkhwnF13/QL3ep/bcJ4rTrB7/oPehzvIBa+PJp3BUYYMpcVdBPPNHd
tmpDFShyF4KSi79iEiwNXKD6qKllrqDI3r1OhhP1p84WFK+m+VRH5pF3sXG4/zR4Uc+f1xClfC3L
gOvLMuhY8abeHq2xJmSmfrLvMnCYD2E7bMXW01m4HfzyMKsRAToxh9VZvG1uNWH24J685d/AsoOB
YvriDc6EysGZpCsaVLu2jDKRB36EdAqQZCHOAhvYwgO1rxlFIil1mNEmwkLhSVv6iGDbMEfYhvmw
3hY80/yALQYoxE0s/FRpM0fVolLSwPZyHkQZmsxuwP3JfD/o2OCoVdcB5pdmn+79/3ZR3DdCl3oz
gti112cIfPFv8w5flRF7l5JzK+yQFESZyZiMh+MSwGYXFK4Elr3GmXi4yGNmL3BoeEavyicBjAq1
BYH0b9idcOTtpyBBvdE38VMYnzWIZSuagmpG0ZKAUHuL4JizQa4mAo70z77F4M2ROjq5PKuFSqPw
CD8vp9w26pZLomIPqHVbVRbwwL7LeJH0yA+T78Ss7iWePWMVzeSXrBuWuRNw6Q0qIaFudvtbHuci
Zj9rxz0xnjOQTF7Dn0EPH5Nf2Z8qgvlQAT2JXsPMx0PIovQpormJdFBnK+JCkhJ2ZsaexJhCO4Y/
d7o40QFX7toILxZuy8YNG6EmjRRtaXi2iez5irTsitTfx2J1eZyiAQhbMNucQfO7iMv8SmHcrDAZ
p3SmWZHlipjnmV5GCZa+6fD0toxWy8ueWZMCDMVbo9t6hXy85PuRIux2iSlxe/+gG2H+CrpNn1bW
l12R8iA6tDQgfqXerSQIKtmbSDgSEHiwz2/6Cm7BGkHCu+Id3zYG/0SILfy4BSA5LGNIROpX1Dg9
S10KGN1Fd8JzCAlpwODG5y49pb7D3bRIrA41HreAsHs7yBQs6wKR1n2996Mihj68oBzwuWI8RSJB
i8XLhi1g+7wTmfBOEzo2g23E+hEuhPM5h5wWyJC8ekDiAoKQIrUfdWwqMD51D1m6xEP0690qzFvX
/KbcS7Sgg3PEFp1vSWhKKHFQwsebTtuu7syc3z3bIaCqPtTRsYtxiUuQLNdohbjexONjb/Q2ZxpZ
bqbLOhYyrA+lDbOgZbvE51lJW8ubKOPsiYx5ftc8kTfZPr5imn5j85izTPhsQ/sYoNPm53BPJIZa
i/XH6gYEeGfR1S+5R1mP7Oyn6/Qxfv/p4IsiGuIFYG00+OkXhmnyUr/VS1KBypCdqImfyOBzciyK
qrCKWPeDzMQ+joD42u0MHU2+3IY+UoRfq53UWFJvcOxb+73tHGAlbwPTdhjFLDKMzxkogRMrzHTh
8dB1Eg/J9G9pc20TSzgs9ojwWuAWjJ4iMU9VIFcHrP8rdMgbToTLxvJv1WPRBnDlfxqOzXQevV8W
FvOXGcQHK8VJwIkgw7W/CsIpjgV9JNZhc083Qb/VS8DouWPpEpmuk+UlElTn3ytt9dYPO2t2wouk
taeaWrryKgBSA4Gd4qEpGoQRjFt9y54i4M9Q2ECT2B28AdgYh51v6SDWm2tEuIUnNlOzhOhwpoMC
SNdf1O/iCZVV53GqbIBFoeq2k+gzrtY4ziuaPmqogBiV3wqDO0YuigzWvXlJskk5A4BRdY3Oo359
FgVU0VddeOli/iOB3CWg0EIK9S7AAVQIdyrC+5aHUy9Xd56GVeyrI/93OPGrNiFHIBqWRHQgHNMK
F0z1zH/ufzMy1l89+8rVB0nCqzWy04TiqPBJ515tJrvokvLqocJWvcTqjzkKM0uplcPBnUeBf6TI
QagsrHYXD4bipDQT3b6mXUSpYZzyGG1WZ+YFmT2NKI6bhmRAFzTCtdBSry8VFg8jFXllgq7hh0Db
sKmWgKkpkM5K+MDEKGItDfG1xywM6lIdR7FvO7Sp/3GrFlOFXS1bB3reELbUcquoXV1zZcdr05ta
eTfLJZBTKy3JqKLX6w6TysiHWTR9sD5cQOfLSgjswa3CXmCD5WA2XrhSX5n0xQkkXn7DgSXg5ykH
8nLnKrCswjf8XGtiaV9avfttDy9DS5txyUohRnSvaJfgoUmkyddhAlRuel6OloxRiwxvIbPlatdY
B+BU9dLWpOTc75Ej5BXwINvkQxUY7PxA7jLsmmKDHqdh0K2dZTEaDcxX5d/AE7BV5cWlPhzs3Zmc
8LfjtV8AMhjgJMTzyVKZF1WMbb4wX+eply/WhFq8T0Eq3EW9KNCTXAkxSee/U9fIjsUaUIIYv5fA
d3UN14abVtMZzxu8Z7K9MpyRdI9kZ4Vn+1reAxODySolHoQ+nlynogG66MIun2OwiL4wPIBR+Jbm
mGHt7PWXVA4RFYBtK66Ix8qq+xMK/vteT1BFc6QBAhcmmsHTJSASA6EvX40CBvQc22/OR5ra4wWG
ynor5yWwbX7aDOR4S2SKv/3A3agcyNFrPcF5nyl+R3bwo+0fdttinYtldQ+963IbcY6urBGcvcbo
oO1OS8CPr0L3dOVEjWv66KqS8xeF5YO7XlkZHhmIvqfTRZnzNL9+TmG3eNffJ12atFe3fZuQ6UmE
LcLgnoqzf0P6LboCM6XFqoIqoLNVG7CfzvaoA/UexYIDpg3oUe+mBmEO6peEMMvw8l9Se226VL2x
xGA7idwWwMaNOA5mFTMN4olpOwpkyimetsjxnF+c7NJZ26RzsJSnmA2Ypv0bDc2XzrT7VAJTHTeQ
OiQpqjhRZ011HCE0vvJLg8a21HlJUIVVxgIhcpB4pbywEC0j1GMVFeJ+yUDHe2im9XwIG7SYlu11
ZgT/Jgy7/dWLD4lBNrMB2FuYw0Wg/rnbhAkT71mhyrOMes0t07y0A6XzlCaJ4wTURIHbHAdbDPeg
7JXpqBLiFj1tQMPhb8IGvGNdnyye/BXi+rfCVpnFDKFKRJQnRAtLPqvgN2IdbPXmoky9KmHx1JfH
M8J0+yP4hvey7oBNvos++KC9ZdBvIqsu6VMDPSMBaEGuhbNZYFiDqOJj+AvVZtEELPEREOxwcDTK
bBkr7w5IUaOIcM0Q1wpP7eixtFlIrW2HjeuMyqwhILvoeIGE5zsQLU9qNJLgGpqe8aDUS5oEKhSP
/AAOd58uSptTxnOaVFAuqZUI9VmHVFQKBBlOOiwVK5YAbjOAzMpeCJVjjO/RCCCqp2/24A2EkRM3
6cd/SzBK2njyykJcUkf/u9yk/Z0VExf8vpRP/WFbPGYKiEmJ3ToR/awzFLoMgs+01dRwLF2DqHln
qo+4S3m9bF/w2I86g3CG5qiKvamN8Aw7bdM1xbB6nOYy9PxMln93ynKDdvrF+LAQl1CtiDBk9EjU
3dXL/FuW+OGEZy1o+Jow3uT4RAriIkVUHkWO5I2ibOaNC2F1PHOFwAwfUfyS9PrxbsYQAYeJrfGO
Iu7vSRZEYFtqTolWjtbSN9ceIdR/+djc14bJV24xQtEbkspADmVtzYElfnCaZ1gMmkUFWSt35Aay
MtNwfaiBUM5n6ZreIhpUwbNvaSmIKbnqe2hVgNU4u3yFPa+B9LHWhxzWPuUh57E33krJyfH1jLk+
kVmmd7d+gw0x7m9vjTpePlMLkAguISsJc2ui10DxTVdnMBw78Cjj6NmuXBQK2JkY6R+6rNVpGdM5
e9Qpt8YoA3ci4hHzVK94VASqtvPxApJGgCbuTV8DJ1UFSOihlj/u/QfXpXd66uCu8ESUogSJ1X+u
3hdP7zgnvSLyaHR1rilmCbbANp3kX1dVLUYsVBmoz0wqLoJpAnImk4H5YD84QQ8+7bSi6uni4x0X
1aDJ5r1meAO6mQYWarsVobGHP4TTt/2U6cTRGPk9c26mqr3RYMAsPxz7mEOHzqPo43BjU3MR9I3N
TQF2WJI2v+1TF62RGrPqC53l6CRKWuksSbyX4uiP/Gb9XsGYqhSOzMr1tdkGBN137BdIaMBp+Knz
BIMqYpBHi0/0Sk1Rt7DioR0yGqfcTL0hvi62OwMDV/jFvu1UpsARpgG1xDoPBkJFKaP/SP/xXdGd
/YeTB/ADgrFNig4Q3WvLYpDDdy/+shF6FQ/7V4cZgyOsWUeueXOmwNsegYo8Utq6pdNoKPNS4njz
y8V/RAib/WES0ND49W3iscnP+6EwwqYGX0L03XF265JLMohFz0+NCZRWN5M1u0GRJsnzDNZhApPN
y20R3YEUfS+9t2WYNjZ3cVCtmbHHgvk8WWQwjgZcBBucHUVjF3+x2Nok4XauA2f2Ex0UebJwdq9N
4bkSoY3kc35gMpWJmLD3Gecd6NTAdqbAFUAETPgkfx1He2q7cLuVMW06ka8rXN65lyc+9IrXL9LM
pnvKrIUOhvgjbGHXh9a/+zBgQ86JUTiojhxHEa1aqWxfdqZxJkEfXfGBTPDPh9gzHtn+WHB80D47
X02xwSMqg0OlKq2zPs7J4UHxK6zY1v1OuSjqAHjf3gHo6azGSTpu6sjq30fdN3nEcjtH56xNtIMf
4m9hCyPZSDzqMpjP5IJlcUINhLdXckhfXyfi9y29cupmSpBzTndTJr3gBFzaTupBru8vjvn+cmiF
18/XPzyVrF41kX/XO6/0LZAJfnHep4kSCbamZIpFaBDU/xBYTPQsrjvITzIQPP4EJJbs2RhNdFpz
UOYPw4fs8c+o7pqWlnHR/F9FO1c+6RNloJTRqZsizmXQJW7vJs2/wKIIUY0aJ6HKrXx1qJ10rIjP
Hcf3zLrrCkaU0bnyfFxORMoPchiNGwh3SUOyV/Y99bm1efadeIjqOMiK0mUUrT6dX9LmiH4YkfYY
JqIEopq7GiWNICWZsUF70/NPIcbDHtbmJ70ZXPzA0UUJ+eIFRIjYRPFaRw2AearVNWlzcNmAKLfG
0KEVMzQJzyWygVvyNMVJGpVUKtD+9O7/zGBSqgQkiO3xb5afTWnFrarE3Fi76DmbgyzJCNp4x1HB
hckpQ5D0M74xgMUFm1UTWQLLgTzZMWrco/OF3b2TBcSIQugrK64jMEwk+Gpj4SPj3siXTuAXnfok
d364lsBZW936dQvWJ8BBISLlpxwRMky0ezW17+zaII0iGp9IKgvWnFnEpvcd5Lr10q/au83O2sgI
r3hpV1wlORYJRi5CIzvVfubA1nSo/8pc8aF5IstOE2PrKDadh+CzWW6Eo2C29XPm1uZeBMYZ7y31
7JDx+odKdrfx1gLkORvlPQZ95GcHnZIWPyZcQW0J+DtvD5bFwKLHl3k0ZSoVkCafrKuc7xUXjjxO
TBkKFU2xQQ2koPOOIWq1sakpuXe+/q0vx1IGj4FPrZbMoyPbpzgPmQ5qANr+f29attDopbesj9hs
e7565wrFmyerzE3WfVFcO3ivUs5kj79fJY6q5wR4CEOxliqC31TLnGNfbu4bDyEAHuW07iyI44RB
sBcHrgrqR9cxVOf1qSaNdAu2shIt8slXQPSHKD8V5Co3eTV74igyJ0p349aZzabbkWocmGlH1d3r
ldsQyo6KYhYRG3EeuWzKQxQUHVwGKf9lubCm0vjmgjOtK09wz8RyAkXidpRtK4iXvqZ53o4UHEW4
uoxsWixBLS+fGhLitLs/AvoXM/NaWLkPn1g3Y7YWjMp2a9grY1OgJpEA7bsEcTvRQIQaiwRF/jOz
QgCCUKKC6UYudzuFdQ/Uj/2ZZu6V+iqCtNppxXyYkitR+1aAS+eBUH0gSlDd5JdxWonBeGFqDf/5
LK8GqmCBj876xdnvGbTBCu8lyW1oEUUFoTRAEI0u2jft/EZMrNsMRuInro/135mykCthwDnuY3PC
vnFOwppCxYrLeNXSTGd5vB5KrOELwBZFXdlzTq/ZYukPQ3cbQsjtuqFagFwIU6D7CzF57EjHht7K
KBaRGiJBzavGQIqWwiB7Ihp9OQzniIlrdlEawSbrETdip3JAaqQt40q7Fw5j84I3ENv9hPNL/kg8
12yqd86LOoSGqdwxIAbzCxvJIuuueFdSmXguNLYQu4vnTXun+zQeDErgCmIjM2Xq4KKedTChrT5R
4ZX7Pa0btWiv1QCKEJBMBD5UAOG45gc0dsBgYLVZ3k0vwfsV65MA2d6DTojVmtWOfbAF2nsZYR8w
PCmrr/X2+cMsw4LZcanDzmJKUeVcwYxHSe4D97FP/I7g1it7p7NAaYfWwS/uLJcpTJ0UK2Nz8s3q
cDET/AnJn/He2i/cja03nVBGSlFyVulpcPk3DhYGL+Rncwl7LpR1CabYY9HWBru/5GZsrpjK9SFZ
uzbAWgtCz5qRQXVjp8UZnhEhroyyGYZmWV4O53C4tApWP1np78z4RsDwshib5IpJHObuJff95ODv
8doDCXoi0ewiJjl6butQxkjYEv6rLMMtufUvzqwcMg7qBqOLg/X2dhinczqd6AGRqw6rWrJILa4i
aNHxe5h8hg0QclDO0s0D72zh3rwP+T7xHYU/GdnkA//3jrKDF2pEfU5C/ZrGYsEl3CbTSVqMFiun
GKFTkNl0cKBG5yufmyDFIPk4EaSzVMIZ7bqgTDwuZc+xLd0i81po59YtWi/6QNp8ZPi3xv5Qce0E
141Wpix2vr38bZgF1SDfXgT5Pk7F8m99gKDojALO+s05Y8e5Lw3Ff5N+wBMKNBABIoOsv/FWpT3L
HY/FrWT4HPOtMqmKWiKPi3s88Ro3fpN8VHrXvWkOOmLKLFrqBa6lJkWu22dlZm5LjjIJkjE7L88A
eV+kFi1WzTfXObh4Fu2wEEgNzzMzwT7PGnUd9i+eGWpGlwvMBeQKL3PdROYeR1KQXu6PGWhjdxbk
+iEUWYmH5HuYxc2FrQHTfT/B/gf4cXc+LW4BQ3OtROQd0UJfU0DEMgnWxfElb5L6d6oBR0hYdD/p
O99d5WKPOjdSu3RvaAZB1ToGS3jbYcSBZ67EUF1z4hVZO4Jb660h/fBzp12ortD6HYMYkfiNJCmZ
3ZgC734rAI/b7Coh2FUpBqGhqdKJDvu0OYy1MNNYKW0H1UcqPAj6oSMAviLvF3juHrsgrLqi4rSV
/QYoiheZ2AOxOU8D8QUCmajgNImogCWoQZ8GZTWPtHA5fXGW+zm3fIVdQFffCtiIZUcy9lLw/SIk
23RDL4LMK9nmPlinCF399TQlIeN0TNpOW6hHLEwtLX8xIryeGk0+bfwO9RBINosZymLVMXNh7xPT
EFVgascZU6eOpTCuVCJ1/RE3efJ9wF9BtfUzFK/vO4njCm86fw/bFl5/Tipf0+NxhM5AY/p7KARN
nKTdONNS5W/OLIHk1sH08rJFnzWM7smXRDaxgzHTn5nvQ0rdKLBHbuFZC0mW2zOJD8JY0vA0uvuz
byks8gJnGxjIHhDWYpLXUw8OtscFESlAw6zqbKZJjyS5uaH+pYJG5r2MwudQvwIsvfrp6nhmt7oD
jH1Z+8FFyZOeyPKU80t7csYZYe5jzb2CTZ8jASj3FAi4sl0UqkstZCOQjJyOt3y0j3Ec/22vRGBk
UQ10wFKlQ09NCBEwt4QwGQrrntmg0Ajr8vzZIfZm4fFCvu/zYJx5qFuRobli2D41X1CyrTNmUBx5
mZV3eH2ZDmuKh54YdljkTE0fiu4/fbClW7ObJPQ/0BAwNtWQNsSvLxxDagU74AOBqSNbqyG5D+Cc
aDCYvUh124I4mz/9NsAp4G1ng2WHPlBOTe1jL2WsbP5srjE6CJo9lLLpb3Sx1+vNGMwyrSc+hRVE
N1jCp5eRDAfz/MZMeCedgxfcUZdaVt+P2w1qSyN0MD7hpHZqhUKwZKPlWWHlLYUl+Zd5/Z/IhGgg
7PvmFjTNL4MCMUMQU9/CJ4BVO41TQG169ytLUKcTkkmCGuEm2TkQRlcxSNFOXbmRniv+4ok+oc+b
5pkpEZ29BwWSgx8EvC/RX2aYp3QFpus84uV4Qd942AnuoDeOWEcPghXKVjlOv5eOVBnLUXZs99Dk
IuE16QK8WBEh9QUJzDmgCvV3RQXsGOPdMC/0mWNUWYjd9lyOCGcwQBHaxXR27WfTLyMP9itlqY/N
zGMMBFvXupdZ1lFaLL7hcJ+CJH+o/+S2hc0okKVagIxF86LX/2ZUHbWac2IpdVXDTOVwhQnx0qNy
NAfO/KA6s1Q+Vn8bES+/aEPv9j4mW1+hsUbvkkI4oCrOa4CSfA6+Uf58l50p1Y85u/Bi67uXJBa+
sOQCPwX00kdtFMgteo3FJaf9lkUo9j8jbVx6ZR+IihH4Jo7Pf4OGznfmUiVJ6IYX8YzRbiS18e/0
mrlpSrgyGt2kBJObnbsJ3w66TeJq5CIQ55LHwypOdUWUJGqiWaMXg9pwug4oxyG+arv7vQudwnyG
oEMPzsD28XaBsd2WR8Uf15c0a/wcv9v25Rtef922BjilbWa44xMBtpbTk10aNFlQkVbs3ypiwf82
PbqP0yGoCnLOsVlMw164r/LjV5eT9LZEKiL09MHCtbiG8SicKziWILj9RH+nzsRZ6CQCSF4lvd0Y
vOr8T7ro67hFqWyY3K5tZgCY1TWMzgP88jNOiIXfBUZpeDjy7t4Fsk3kRanxRXGV/iPN7OsaEmPC
YOny3xF0Gru26IyF+9x+0m8AYfrVpy26e057p3GZBPa6VulLA8gZ1vk+6LOnvUrk27SpEGlM8AIu
CwDopOVv9cNYNxfsHssI2lJaeUgFINxJzds97T+Z19v9yAdHU1G+FizkAvi0Zzmb2MoC1X8+ZC1Y
dv1bUubycTdNH4GVHQYknWHEXXP84DnmEkrqq57OSgntLera50ZnPXLn0JiqWtX8CTCdfyg9Rvzf
cSYD6PeCGpzRfQ6NodnN/Bhr6KnY8s0sUQMWmZzqkQiKYskMT8QhniEECAOEtZFMIj0PTBljjDnD
uPSUxpTNNuKy0+Z59OTT9lH61um9VOSO8tl3/lp6GKhSD2cLOTohKLf2NeUORwwY8vRG9JHCwM9Z
QNgZ4iggL95zbCLwJ2sxKiVHSkYZZUOY1td+64sBWXEA3R8hdE7ILPJFS61imapTim3n7ZplvPN+
IBVoZybaGRjX45jvrW1XW8x7AC0+HJLQo9YnbWIJs5bY5LGZgPTUPlLGvQ8aazi9O1Qfz/jhAIX8
yeOnqOi8R5ab06z6sUPUgvYcDemvdpP+1/IHjgdvjjmukrntvCP7iyoXjoaTkSRzFOTiKCCiiZkL
2mc7PRSZYsnPN95BcDpeIUM8svMusQkTrboUy20PzN0Gt76lHiOc8yU1Ei6/OuqIqneH3k2PKQHd
1+4tLXdcbWv96B5tuD+iHaontD2pdZDT0WITTPVSW4/KYw6N/bC84yeC5W9A1vMkoM6jwJl8HKCI
1RE1/8RDrzZOWlL0EvtSOOrjR+HNoMvUFWlNMuT8P7FNRCpyR17yjbmdVK5E5mxAsONKH7L0g7b0
gG3du4Q7apWMDF6GGRzOvdtMvt37abe2zzqBIvL0YdCd9Q4HVwtL786WYsafe6/EhBtmFFigFOrl
g7RN7c3SoK5/LmGpgpQJ0dxq0IXu+f/cDO2p9j+TIbf/ulThNmvP18hdaX7x+Fa52m+Yzy3WJEnD
BsND92u8sWSih98q5il/aAHNrovAUDsVhE8aehYv1k5DuMUwh1gWeclQwSRmTUJdluVSjYraj3lT
JcT4kt6l+14uhONCAoS3/jcOMZahdEOmVBXel0mxgSZ2WcN7vUA4KHezlfuiYLkycGWgYSyXiS5z
5+IrJLNjS/xdT8iKMu/LBv1L/OxEsvr8sCEsjG+nEOl6TOI2520P09hLWOSw5YSkiVfsV2gcokho
+Ly0NYC9gSyk9suD4mapxx8fqKjo/BFu6DJvzAwjIDo/Ne+am/nIoPitNUFexcPVUsMJJ7s9SZc1
gT0OYbkI1FlbGFxbcmRsg5uyqRZ1QZxk7Py+XY2khveonsOvkyu3W+E1lFi+4h/i7+SmjaOpgZ7x
MGLp4AyS1xTi6GKygMrmbdEXN/mlcCADB8R4vFL476a+VQ6Q2qi9T0U5Egjw1Mds8xJajdaZ9um/
R6uA8qdP2eJNlFWwluo2C5v1Bgh1DzRMXvwb+jtN1i925I4n8YSS4hFoR130dYOCPMhZjkGVrHey
lQbSB4UEJ1XWcNhjTuPLmU3xeVZhTGDxvtNHx2d803RcocSt2GfHpT/VCGqgfeKkwKw+WhnJncs+
pd2mVla9QO8klEd4uDTDQ93IZy2KYZtCtMEzcEhUOuSlI4rf14q4w5BJdBq4hozuRmxnDcNQ5GAf
VvZ8S5A/4Bmd81wPB7Rin3kSYn266AxALv1SVf83iJJe92vM3C2iQSi1+KT0anOXSvBnR9yX4KkX
EmDExV5k7RpP/2BD0bbxHuxu2PofbxJcGkdhcmHuRhhUK6MOkOyj//qv2/TRDLEkAKxHEBJ/BnWz
iHIh1IRzFW/ksYnlr92l0DcPqeG9qhqfJsORUq4CrjZ41mETvOYQSrDv4IO6gT0nsz49upTq4S3L
W+7t4UTTPSZInSHN68sIiPSHZS7OqeT20QrRdzu9FdBhqB8rNnBeDTuWHbSuvfX2Y1KXg5uzPVR/
IKxUE5vSY1jEoSniMoLZTSK/YRDfRswCj60SXErdlRdwawsA8z/mhbdxSkLSpKirXvMJYt8jOo/7
W+t1lyPRPEOkqTvcRKKWmbo24N9arCwM807YT98M3bbq8GW0r95CkLq2V12fmvcvVcs1/iYoTYxH
e5LVa9l7+u/R/SiuT6BqeV0553F7bGMqv29i6HSPdr+CM4+7SW+A21IUOZfNshT6ZGcbYfOkIzjQ
Bb3uN/3Td+p9JL1nFT30xL2e28yAHkHFRJR9+dMVwkPuKdWaPzi84hOJCbf7fDKs5FvvjyHUId0e
CLaEoX36zT58g8Qtc8hiXOap4GP893rWWkyzA26C4oEWGK3vhh3dNTrLYkA3NFsZDP6pt2VZ9rbG
uKB9txCwbVbx2bL2QbZS00XVGPyUaQGwB2mxksEo7yF/VR7/u6nOLaSlTm3Wlau+6gyVBpsUBr7K
G3YI/zZ/MfmGipEozjlbhmqztouMrnnOW42UKAV92HN8YKDe/DLLl6q63rDnc2lIZ2n6W0wC8kyx
zeDJ2g9d23nTSPmHiFttWDJVmP1ddUGxD6tCkCFoGipMsGd7KxncQ3kc157iZXbzO3fw3q00hE0Y
ltKO/mauH+qkIWBT2giUNfwxHKDPdA57D3hQylhAdhsbeKXAZJSIXVgQ/aos06+TdnF4+YGH1cs6
unV7UVzFr5Pz5R404Xxl7Rzw+rc5adPYsuiS8bB1U81HZEZyAwQTrG92ei75/I2mG11ourC0gpv6
/+V5vqwKCjNID1rXav3v13MLN0mFDQnQYhNZApJbW4JiHFtJsQ0RZJ/l3djLdrcUEmZMx3ArNgc5
OQt7Wd/6FXbNgjZJ1WFhO0ouw1xnxuJgPngI/gXwejFR6/l5h7MFafC9HcNJOTv4tuSjPTVAwxCQ
rPw3J3F9EdXfaurW2kFaKLx5fRhOm3cQDYYybWAtbTmpLIcblpaz+9orC4qBiWM5Hp7IKZswwbtH
zSYJCOvoqX6dFzX84ozLQdh74+WpF9HNsyBqzmFIrgaI3KKVR2XLs50X9wEm0mMemfVAxG0/dyqR
H7uAYRrXUDlxMWKyn+277Ythf+0iFax7Mfp1yml+r3hDA9+2IPZuV6csmME7tNqREJk2DVaOdXeR
mztbjrPDX1as7oA5pEuYdBvH609rG/ABp0gQErgl8Eokg48/6DQSRBIrqQeXiYeQ5mXu2ZlhVP+2
z17iqkpSmQLNDm2Ahv3U2vH+7mK0uWfQAvBhIzCaTtTgHpdC+wZqHIkUqFpkU16+q1btl1Mfr1Do
jHfvPZRFqdzpNZ9keG2fg10dgvnczonJWIcRwUU3k35DnZYV/l1njM1pDWwQ9OwJ7fA8bxqpRB4b
zNTTp9qzfJmfQvmaJghT71tXC7x/URWMvizP5qZ8u1pYYbaw/9PNrbfBqTEfQhFtOLzKF4514I3X
JZUskpqvEFCj5eabscbGY2OIBW0OfFJyH43A9SRfXPY7+jzITATi6//cvm1ENorVMkXKWgMTgdqi
NdXAOSdmkvUcgN4OxPkXXe096AEaPvPuFaXcbZ6NCSxTov89gCtXiDGtZOuxbgCeoLErlB8+9zLa
Pcnvf8zxggPvFKQ12VLr9cqkThA65OfxpJD6vgXNT8c1hDEW8NAnvLlJdZkZLMY5+86LTDfoFG4E
TDRnvbeyT+UXL33tX+3z4rQ+Bt0sCQ3JglY387akVlM5bovBaP2W796UpfLgNSsOsyAAP+YX5c3W
1M8cP3GCQTV7mb4sTevkkDnNnB9nOxkD9gMvVl43ghWocC/XZCp40lRyXFJW/DOnpdg1SNRDoAi5
u5B3ThtR2Dj1sQTPN+r1w/dDIPChOlbn1Wn0RcRwsNIP/8uUW5W8iuvwQJUy0Ru3jiPpM/V1j8d3
rnVEP7PmAuwjA9yEuuJIIej85NcqJ+hu+aVDcvp4ZNzqaWxF8KS//SEQkMEcFKtqNKjmuvM/pgdt
ooXzVGZPPx6v+SeMmGCz99t/p2Ff3YNIRfkig89Rt6FItdvMO1KoI4I9ezvBKPDhSY3bTYVY4KcR
zkNhJZq54QhdgstrQN0PTFtkMxyWNTuaZdhl+5WVraRLsvlP6LVBwG4PYHtt5FMuN4Lzx1o+1xKQ
URL6RbtiMrx3n3H3SER/3L6kv0Ze/BUDPxIFL7EB0bOpNujkg5YpbCbXV1vGIfLZ3F2rDUAbekhj
mMOdGKlNeCyrWtzM+xLqYt6TM6rBNSFKKxE7Her3EODKH7dSYoD60bwvToMfqD3YKQHBk923+dWh
Umi8B21usOaFjvRBMjvf1tDU/h8vovqtrj5/9C6Rlvvk+mXG7SuWQOvOcGiaSOAupCBm9ZRoPbVb
NiZONBmDYMqTqvJNbnpLuD3S7VkcIU4LnjxZDZUw6Nx2L4mzFmJGocT5RZYRMiNvvw0kPCq/gCJp
vlzwxK3EIiX5USVh9/sCQCl8Qjs4Hsy3Rbe6NlHYpO5kJsBYxTKyZouXAlmz0U+msxVkO0c2TbQ9
W/jYG7g3VgauCpkPpSjmOJTBA9pX5kLPQW1yt3I4ATzp5ZjiKpYsTnaEfCPwcPxjC88Jvy68FG8U
f4Hq02MRtBlw9hNNFjPRm7q7qUGZC9/KoRgaC6QL5eAHeeQ71na+CCxDtMyMdYO3WXDNfyMvlJU1
kZB+mbCE/iMyStYPzXRShzFrAU+X4iRxBkUUWG64MQvqeU/+TxYd89bg8jGUmV1qb48W26GBQT9K
127TNIDpiDSw2MP/WUN0NCOwK75nk/rZrqVJkfoe+bov51KH4zpWOn3GppK3j3+FThySYbdekZvK
3978VRS4vmfsH5op/m1tx7CYzuUI5V00cR/mkB0lYs4UvFtWpxkmPSEkmz6tD9e5G7Bi6E2u6+tL
sFZeLYY8aYOzQbiwIG3yyXyTDeBqEjUcZwrevCQSSnNmwm9WpjwtyUbsQjLC5Cht1xBKymifzwzO
flMUacIqWiXvHH5xQsikzB2tf0S3ADQXawMXrnb+H9sqcz4HNGDhYaDSKWTWAlLuxN3MxO/kcGcU
P6SEkDEs30bYCrLtgY0F9RLh5Pg0D04WgG9jqrhDFALdGEUt8xJe5PCVItFCs+vRyv/GD+M85sWU
81Zt8f5elMdarFWCnuOOgyey252cGHiwaZ4pyA76axMpkX/UHjm8jbB6gNWE8ZuH/C0HDm5VgRMB
lTyOLqaa2JoDUmn9qN1Zvi4aWtXFqdEo6gluxeGLdQnbKx0D7kzLvYvRMmX9hWSN8uibUYfFmSAl
Dk+q+4MSjaDbmgYpQrMx7MyCFP4n0cDUmUHVJo4PszVQQ/t/QHcmAZ5WKbTIJf64VRzdhHUvIsms
AetP3glsgQTLokD5n93rFWNXs5Yo8NFLmwRrMShJ6oVVU64J8btgzCfKbNQtKeyLIUI2vllzypFX
KLwg6r6ExSuWBzUWvrDpwK0sUhAZ8AQ3k/DLM7YUozM5Xz3O02wSEh7r6lwhcciBFvgdllIQ5dBG
iuPk7tctQR0mgUKmKyLH8pxDyM+uc82vyoIagGXhuWjl52gDY9TjI5aK4csoOxAOjbDbQJfdtM0G
4xF3+Soq5vaLtq62MqTvFtfX3k9mCThc6rSbopKK6g3hsooScGojHt6sFCNp4smhT7Pdv84P4SHf
CANVSyB5qLJmzdaYQmBrsiw+za22fIyuAJfnaAg1BcL+kgE7eucn1/5xuyirBZ0WcrHob1W/q0cq
ms1w0jLzpZ8r8/RKpRQI0ueH7wznvavAjYQzJpchEE3RS0C1IEiU4vIfjdrbWG448Ynlb3gJm518
zVexYSr8YKWscnVJMlg3FbHHhyHQFkf0U7jSsHew/+IPR45RYy9zu2g4ciVMd7ODiKY7SiSZm7jD
naJsRyut5ETZBpBx/thACt8tvwjExVr4s8LnqUGyoeJiQ4H8eFmmx/NX8Si9enKGzC+iUaPDrhxm
wP3BVZWNZpdM2vwb04duu7T7IImdH5p1fCmliM4rk5XmhSLBkEENZl2mxueSlmHPYRMus7Iw6Y4P
vtRY2TIu3kJfjwYS8kUvuUreDt8kB+G9KEByKPsP/RlGn64NGtXeBMFHW6K8w9z+vZic5iYP7pMA
uJ5MTuI1XalL5VcyOuN0kntdnPUxcJ6os5px/8fyhbi/azyoCmMykTmz6/avE5GZduyqjnFDFCv6
HDISR3qUIIPmrUOeYwtUlDfU+qTNoSIxwDjFbnYVKDi2V8R6C7dWeyUKRWxVj94UaE3XqgKeo3/+
SECu+hV9xlAbgzVoj+zvLYnyvbnGg10I7ffHSvA4XJgqoSchJM9FEXgiMLnkeL9aZt69d6BnrmwU
Tg0eK2Gev1MO2AKbO5O7VjoQMG2jC/txr0dVAB+wFuhA4lM6jRdqiFhD8NZl/QoguteIEMLr1eAA
T/DaZmZg1sCqTD8HoM4ONnPPNC7w9fuc9H4JVkvgf9H/lGTo131u3MTfivSj9rcxNWOBA+aQWCQL
UDlUIAo0HQY9lmY6SzL0ySrfHR7V+ug5aDVIthuCAC5/DgUE6Qu/KSyOeYFfSTkJL2oDflFCzFE2
pFkuXZ/Jx+V7Cz2khGE3ezkQfymnuPmLIOPWTeZ8AIveylrcRili26h3IiMxCwjs+fYKh36ZqQm1
HNkZuP+n4nDRKabuoHGCVyDFO8rbYTV/+1BTqN3WGwmSlxxl69h79Kik8+8OsakpL+GblhWRBQIi
Ja9R5Sh8VDshk/9rN3tTFQ2G7Q291PG7Zrk/oMj8vOVttSb0mmnvzpe0ftoR7TlA1YgAR0/bl2uP
jBoFPDxHn5Sp6Y/BP5JxTz6PB3i2AwGPtKKqPHrLcf56WpLP2/2Tsi5JRkPQOeg7Ttv1cW3qXNk+
CttNF/95HNZDcOS+I8LjzTxniRNvSongdWKIw0bPw8lnrSsSAF650fLbelbMRPFz9zlYbV2sD+5s
XlSI11IWx8DntjWcT3URsf35RruSz7CFWrven2aNwewZyLb8n1njHGPq5+QVHtISp70srYwtxKlW
2zt1fK2cnR6YTx2gBYxZT1DlpR3s/JCiaHbshPEAgc52gukL4qGVfvpaj/S5iPCycQKDawHYCGUz
LZHAUNqv9LDf5wBXjwOjydApp3JSypOtB2bT70yskBLpJi2sIBk+9wfUCltPsvW4teSYH0cu9Yna
SdyKgdp11N8EMbMKYGSWXC5hfXNEOOO0dv97MdPHRlx0InA8RM4Fc9cVea3f0YtJ5kOBUntODdy8
T/c/kns9zq8cZF9R+63n1RPWCkbJTCXx/n2nGT2KVEzUposkRqaDjp8vJ1dv3aGRvFc6tAroh0cS
fBAZZgrfPS9SKEi+JHNzPkE26V87BdkX0hKjwZy6XB72I0EN+QfgSAdsdLLTK8CZLRzRFckbm/1d
7YTdT1Os4cheGBydFVcEZP2c7M2brEWerSwGoHwdCZmqCOpFvVP5kzTZe9I5nYGSjq00LGgViwh/
PQLileJzfK7u3784qN+8MvKvCsoI0TIDiYqk4RkXYdUWoxk0mpIaSFW3KUirqY08qa4CRYK/w9Af
YsjUrNhKyB8UU+pUTWprT3zMd5A/gzOydXPOzyj4wZzba/kH0EGt84gTYsNcimZYWSXsUuaNBt8K
qs3ydoA4qAS7zl+6lNet5mWIo1ENbKeFSIxZgDfq493d8m0J0fRMLxMWQ9irYxamDJlNf8sILqym
86V6dmLz4dJp9lBq2vbs+1P01p7J70HUuBk8C4o5pNRvTI5o14RZt8aDFK6jmcqjWdAuRWjljTAh
cmS+Z9iGDS3htn4+DzVcPuc5CUB4U79UTXA9I6GDCtUSkBAmLMZBQ0uAjKLBLPSzh9xCXPkZuvOm
lzUVnn2rSTT2WKeyYOHGWdnviXlzawSE4UD3MnEyUaqeG7ruVLxLapvuha8nYqOfEoXmY6Wnv5LN
XqqzF/HBZxWqLY/Pzu4hl/1MQi19lkARviDDPZK9DDipq414inkIozU7kJBWRO2V2ioXNYGBKKB0
A4L3tM18q8GBC5fi4CQ544DAbPH1adxV1H1nLshS6J6sFUdEc16nl/6urmzXxvAVzJ84aprDcX0y
TFYNdljx2GZaCorV+6N9LHI7kgMGUWSwTb8vA/+kdzgEtfy4aLH85YxkBd69JMF00EPib6ZSWNbB
zQ58aShphadHQMYD76KahLdt7LRhOm082nGCnsVX5GOTp12ZpV0pMvWbSxz+Dzs8A9sMtKdPev0z
k3QNoxi08tol6qanygyvL+H/F0P1yQa16CjXaAqm5XzaWVJDWO5Jc+D1Y76cmJOevC6Yzs+2l3kM
EspEy1vyoWCrbqVOVgkkfcCcqPnB3qjSinXUjGhSKqBgB6kptwaWC48PB/p7Hkba/b49pp6AeADC
cZeVS1g+dzZKrCeQWc/qbQUB0NetQPAa02pFjKgenxekBEI8fTTcwqWEZOUC9T2cpEu9yEBhN63V
mf4NDSGHECwT4uRBi4sWafwd2KVAkhUp62BAcNQ6NLMin7hjic+zWF6Qd7j8LL/OezpQiR9dZoBM
MyLb4TFlPHZIe8c1MTK9wK4FwL6XKurcJX3dyrZ2KZpE0Ss0KTfGaw334OqDsS7P28tqxcbd1Vwk
D5+FB/Gmu3Yit8BMe89949hufl5YwF8YV5qRzNRN3IY5ewiriFqoeV9IsKbyEOYsVhqlZuZJIehT
rFyYO/i6sqz5E11mTQOElTOcNWlwCqSn3FhzUiaAvoF07hk+WgWL1bXUJ9oI9FaqGOmVyUkmndU1
M+l5hLELmTVjT1FDj/HB3addKJo0smuL28lL4auuYicgUUFaXTDFKxzeB6e68uvx2ti/SHbeguGl
bvdDVdDSx6zwUAvRGqloKbVTXV8UGNXnjfQPir50r2roryGXSNvrKGYbZQQVr95dJAoeheC8ktdt
oK0986DBPoTd0M4HAiH02Z0OPsLhsDPP0Y9TuufGxwmmXGrUHBRg/ivc76KU/eplPMj3/hoLOAtu
/e5oXRw9SUBNUNDr4MqF/imi7L6JRVbhw6GO4OErzyPVrnwZl3GbB28J3wF9hDFg0sTE4mlhSocm
Vijvar3k98bT1oRKkuJuJFmZ0/6meriqU04d6VdSJ8TzC6o4PSgKialXJbAYEeCcQ0NAj/L0Kw27
DcWOppTzFIrwzc8T+mdWmPNqEPxeRLyuGEUnuzhiCngbvJU+37t2/+ceSNWgqY60kHSi9wxAdbgv
qPRhxdONRc4ekqgLP2sQ+8E1TM+wFiYZYO2TVeLawZrZd2gkavPsQbvtYi4ix6fI4Kyr+TXA0fSk
2JRD4HGeuUPNUiPV6OLEEReZo0R1S9Fw/7m+I34/VHGnxo4Em9zCvwUx6jGQ8m54YL7qoFn9+C5a
qOaI/4R0e8g0VWHWCy61n3b0ptxMRqZdEtRjTOZXMNa9QU7QYami/IGe359YFgJASTs0dsK4T4XW
ToxRijKHqKrhs45ERVkmNHt3ymtc+elKbStudzCqecYbCYP1DQ+NtiS40t2SyYzGHuaFe8dpWCEy
ft5l7ljkJasznvAK6Tw12SaX85mcdsWkFN1zb458YsRvO4N7IScxWi8xOeVbtWc2bQkg4e967THb
HYlAHTUOyMvGw4xnRetPPgFOa0D0VvAKWmXfwcP5XdCowyVe2YOpeyCX7eOuwV+NODy/SLBQK/RK
2SfIVjL6TaFaFnNf9IuhUP0jk38+TrxFZIWm+PQASx//Oq+FS1KFCV/kw4lGbDQ8Sn/NeMDrdJkm
9otgLkY/kEn52CIpCnHU5S4YlR7Qgh9dxmdWg6dSKuA3e+p9ZcA/0sZpCWDTGhXH9mm40S9OCn7n
457g6uG57RmRe4LnTE3VVb9XdEtuPYKOGKIIQmDdt28tOHWnWRouKa83RH9MJXkN+fnwGSsA1I/y
7qmhPRKWFeYR0HP0vNMiEpWyUn0v4rfP7+CIoWEU/08YxMPg9DOnVgURrRHorA73pQ7czXaVaIWy
+ZmOGvV14PNV48Brh/hEH5P/Pv2eAm98H0vjc5JWt51V9Fl9qJCUUDrUNlEZ5MYiyfK7JUbV1vci
iX8BX4fsoSoGAg==
`protect end_protected

