

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ccgvBbguTrezyShnY9xAW/HpaGeHavwBvTfth+93Y2So8ZQVvgUaGmPkMA5fupJiO60pXuATtAgR
h6fHFSlc+g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
q4mKJUn84pqRLnyNSp5FvZDsBC3tA27R9Ty7vHTKlyEMNGOZCiZKb8HmbV2J3iuouo7BLqG2431m
CkY32t8fXZuC+q7cAsEXi1a4FeGBeUQ9IkCw51p3xhD/0s8BtrXsNEynK9BdveFoMVLoaDg7n19e
KYJAj3ZkAhhhnRFDyh8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VaYuuvS79Fphv7xg+4ZYMYQvh7CgVaooUisLN2Jpuk38UGwaE5li6PU5RNeTg4DqMBbQC2DH23Q/
MLhoUSWplGEhhCewZqBPfycFcl9K9pMica2Fay4TUTw6LpMhH7HajNNBJnLPejvhGmq0KlU9xPG0
IYtnuZ7KJeAv4uW5ECo68HgpMJ39vU9CjmQdjAOY7jgfrux/5fIaIqU3VgFpIEQCWZbFLdNV89ur
IZUpDvDDzGfRNpWdsaG8Qid8h/KXTlckOrVnUb7uMr6UyJi6rUrbsSC/9iOtXEIdLjbvys0Ra03v
lAKHHp8AMG6juVMuNGzgrVibWRGvAPuh160BgQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
txQTkR4itWkUxsisvv0qMJHQd8t+rcZaRcaCQftW0a445QfH1Ev7+7RACB3OKyadbprV9zGHPuZR
GNZt9meLSv4Xk60uC29jkYfq8RnEhhi6/qKxv6Bg7+OTUXnFzdXrB9tpU8muxBJtUdM0x6NfqjKY
lCYWycdkiTsKGS9yKo7iy7gKS6p3LopW4jol+sl/pvgWuw9aQG/bhkQ0DtZvR+noYTOSj14/MS+b
eDyc2hFUyUUkH4Q1ixrbanfT76InfmBaHzkrMA96ulADkY/IdEVOU26NNUOt5gpf6KBe5PNKyPac
4qTagIHF+iT5AKGBBmw7pPnp98SpvtvCxJqmVw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aW08EHu6MAGRN8QehR/ru5yNHkBlO3jDuIf1S7SFu0Fbj1b+YJ6ZbwTiujjEwj7Iy5S60LK3EgmR
qIW6iq7htJ1vYKzy9DYRANRGrd03BSLbHqlZ5azoECROxMxtZaeNVzLOUmb1SGpT4gc0LXy8AjNa
JapHsLf+JnwY7W4K9omf4PgkJIrLijg03DivKjmYCiFi9HtaSReCv40J1Lf1wElKuGxz5HXCq7g5
Y7C0F68PBaiOL1bXR/5LOBTdwns4krzkwm5eMgU+niuOqxdn1Ml0rD4tUbjIswk1rtBPkhn5K33K
3v8NnbGycg8l1j2ezDxpjM7XEgHVMB4RiZKUYQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
j7a2SWmYcxwtgVQAUHJ9nHI/0GY4I0MuZC03yIoH9RaBnUKXD90qoVwIKhwQT46xdfjSnlII3RIq
7XCVCtav6NqVkfrydLzRUtJkopQWkenHheg//WoTlYzUfPjKFth6jyMob6fTAYGFZ4hvQNKNqFTH
/Ar4HCoXm6ejIkBdm68=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hhKugNyI+Cd8n65fCkDMxK5a0oXLa0EiQ3+awjJ7cSLS6gtwUx2/hbPP29mX8ImEFlULydcBan3d
1JBelzw4s7lytLYSWhqvjIDzR4dXho6V+mvt3oCM4RBSywBLIvJ8xaSwKdRuSBK4l6Lp54RUckvX
1pUj6MpFAFmunraHKY93l9WUekDALrWtNUqllJ0WXuD+PNY8S9YknlA7k0zGkQgDO7yfVlRYHGZQ
rqhEjAOzbKvfRPdWjJpE83Fub6itAKaPtLiuzVy1DxMTeD8MIFriCX7MBj4cLL7DULVax2gw8oNH
+fmh7rmvnZrlt/U2wY4DJDjbGqCBk6HmtlqN9g==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
cEbyGTjjFU1sV8+iGdkdt/bxOdaSbx3sxU0x+KbZbSoHlLNKQn4kkSjAwpxXEXwp47hIRL8dTRg5
F3kv/cRMUIVipZPndplQQYB2JcTC5hZVOdL8UNM0edjyAF7CaNd/Ig+uAjshEsslv1xrHZweKYz7
ZUlxy4M+1QwiBGTZSHRDUosbheIdKJP2meL7NI2VBAFeX9xnc5C526AWmlbEyjfUIGyqyKDNKyiL
Gl7pcqcBdhTZMdPq0zLQCkuC/vQR33AeGb1ebou0+DrIh1EKiRmPte3/Sqpv87bV86C5I+LiXGcI
L0Eja0Oi9Xncsyoc6U3cyMcbLKBhb5ZevHd6Esj81X4wu3+iKtij8qvQQAFieoXbWMyPqyae7CYg
Owc/v/2usvVnpkcbWeAfxTp422cG/LUipCSTG67uLnrIs8W6euF/4mORsPxCksqh7b0UhPmTYUkX
cNdnFSxtHxvJMXlB4W4Ytem628Iit3is1iP4tb9NR52C6312TstxkkAO8tEAxgEV9Ft3EbknQOeW
iTmXSaXBHZ8M0jalutxy5k9e1cxDW3KVumcSFYyNlwv7B5/SXrKTNa9JJJw97VoSQr0UBUP1TUt2
BH9X/skE1ytnUBC/RMSW49On9Imb75er33d4xcF/LuJpoFRjllcbZLaYolU3nFMM1mMyrwbNLcRu
NUmBZlXDCSJ5oSysqzqe5+dfbDIGodlpKgEbM3f1BwUuMPzqqWM/ObE1gRCdlXD2QFGvqAs+nhQX
kxtGFB4Z9hYmowfcuPNR2J9S+/eevTCMc58qh5owU+e2NUObKUY3eQaezESeKBMJKLjOFB99R6I7
d7n9//L9cyZwLZ6Gymwc5MHkchFwpaYrDHepdEw9neHq2zt/oMm7+pX6Zdr0Jv41C4neKGdDoRGV
5+bLDCnJ3pPEZS5ucPQdIXfK2NCM3GYnGO4TlP+Zfq3NwWl13hezbWX14zBE9UBhO5eL3EBiybtp
r9igMlAPJaj9AADkJ0OEh9NszkwJO10n4Quxkz1OOiCcNIQRaSwi4PvgCT3rcBAk4QyvUz132RAK
OsJr/DUPKsqyOEeQjYf0D5b1fSkxbcnngJvTpo0A1ANbQPPwYBrRzIW1AXROIT16j7XepOauzUFI
S7PlZVpgZsly7RZELuVWmUEh1se4BkiX1JpzIS47fE5A4DZDpQ7hLNZyreYrVHOBmEn0aHRPChJ8
d+u9NwjDgTviUoCKC0C5v+suEW0fqzl8ocm3yucL0hCBTEAb3vUtnQFOqzO8WER7U8ngzU9g8OI4
kw/rxCbKm5UHs+x13E9VFPmfuqH9iUm2ynmyNVbI/n62mWsYe8JcGN1JoLVagBEnQzB1G+/9PU/N
CpgdnpdvgIkQIq4IUX7CNYOcU/dflqLb+Vbvddx8cZv5yor+5TJgIQ1Vg3WfOegf8m+1+faOW6io
xzNUKd0iKms3BpG4ArK+kR864EaXGYRTju3zeDYmfryDzNRszm+o0tAJL+2PQG6Zr+n9yyIfOOC/
D/Cny3uVD2a5RodSvgVz+NlmcRWF/fHGLUyfc/qG3Ka/ZVXzjr2qGmK74fOZwbdhDwAvKCvU4XPp
p+rYuavRv5DOr31+FJJugRTXVnybpM51hOnp5uhvnnpRGaPxUfbHria3Kzck1mXYkJCadC/tNVXa
fU0HK9DEskK038S/MwODch4BVlF16RagtLOpZW69PeVyFPiDHnmnvvZEMlJoixp+OwCZzuwrjsbr
T4cYrcJILYP2LpgHLZFB/p70KVaSdRQ/ZAKCO5wbtpp0l5N9OggXz7JyPzMievZCdcwwubSJe2Dz
XUY1uAGsylBuEPgkThwyrH8S2HE7ULfJv0jjoQz8H/W2wTH1jNXLJww9qlu280WNzRs2XbA6fZSu
vzYsviXVAfnJwVjLvIrKOODR5UMX/dHXZt0DgPGKIRM5AwFb9+MDCWj/Xx8k9I7h52K36vAu9ec1
eYEIhngsYIm7yAlhSHIIKY/GlRFAYbOrgnyogZxjXx8wbBEXgPYku5KiBUYj6MQe8Sutyc/aSkGc
+x92Zy2Y3IKK7v7fvEQSqbJFU9MPDNSnuTMz8oy4p+YSB9bkj6rzL1z8ER7eX5dbc7I4gAAqWWFu
0x/zTN6HqSuGKcaaLNn6Aldswob0Y3tYsv8xfS/7ejQiPiCZ9m9oUCMSB7XMqvsag65kIEsg6nrH
t9jRCLu7GRrNKrEIzoXdSGBL7FeujHVue8+MxeOBhwYJQTK9m/ClShnVhdF9M413wa6XJJEozGgj
iAmijZV29Hj44K/tBZ18j3NJQRcBT9odBDYe7FyF52mGVNBn802FTyBeFvXngOhoBLx0xfEwmyEy
umdAfJ+28LXv9PEp/S46UmsYpDw+fDZ1BQKHZaFsThKsqBFS7y3zl1r4pD/mthn8/PQdLgphFhUq
qeKcKmasbPe5w02bC+sm0pG1U1Z9oc5IT8a7p/sWyqYxYMbCzekBVY031+P1+C3fPOQgyg5Ix9sQ
AlT64El+O5jwIDJ9o1jA+0AkB6oTKJK3V64GC2bke5qzp2asAuM3ULY3XU3+j5SLaGd6jTaLJGQk
UZpOoHQhWXYPajujhMH8ga0mVxnjrZYP2RRiHrMqtGiEmKC9phxQBnucfIR6cEjDpIS3QVGSMQQB
qEjEfpOKj8/AOflRFRukNMiH+5sd1N0fz+iJgya6DKQx128GD4qYypQ1amA0ySTkQw4ouxclQLGb
eemBQSgcucfwuo2S8K6CchHfLTrL6FhqmvsYZzYNH9lmIP2rjEq6AAddNWPRIKfGwdUFVr6Maw3G
b28QnNb8M7Y17DvhnTyOuA6z/HFjPGtPLxlWd9mEVX3HqTYEMTVWCnWc8vP6wU0LlT2sfnDUDgl2
QwzvvLgpIfnhn0io0MC7ZvOVfPUbtGnyETb3ONrrFV7sepqUKMGSciilo2GWVLjzlZ7LOFCLPWoH
U0bIDyTCd0X+1hliJssVZ30036oRaLQvtjq52xRiaUVjBh4GiQe9+C8nWiIawTJWZonFMv/o/gFn
M7pDVn3SdvO8P+OOphteMQr4bnyHhFwiRvGSwvq+hf2dijGt6kkWmlsVCLdVV5JGMZ+B1sxLzzXN
eSdIwU5zWhKTpl1583aGTeqb+WZBwBktzGn+Y4Wgdi/FbAoIS7yMRf7DzV1zABKPfJBLcfUdGKpD
JpRe1nwpyEO8hTIrtCATOdoewnp3q619/249QXiPvVnqMcUeMCxGp9cddaUBl6Jq3zWrvOJyCKSm
D3InQ/Qf6w2GtGQQy8U8GvAMNtFIIc/8MRIymAjVh/mwweRxXOHEl1zwhWWCbjD9y1fslwUMc0Zh
XNmjtJsh0l9KQmU45iE0aip6TipWycweiZkc+OVOyjnudGQHi6b6CSl0D52mSkWuU8w22S6VxzSE
t7yaCVicMnes77VGMaSHNnkHdKAvAsK6+WBNsb10q0Hg02PdLBPDnT3VKaoZWaFRYaVnaUJBG4ai
SBU7qmtMOOiq9kh8MjQ49agHd/PXiFqB1wlEr9ndurf5JJy/K+j9Upw7x9vTAEotHsideWOEo4X2
JJ6YePFp3Y8ycWY+pBZ7SiijnCUPDR92MaQ+2v33dcSz2/ILeyAsWF9V9jgUzNPkUzpl7qOYVA1q
9guAc4SZl5PEBeUdjKUxPNyM6YCF4AIDCVX135f08DS9LgaI1I6KNYfKiXsjGLg67rSrVxLbnDlk
o676CSK9jmwje85RJM20YQfswGNCLL1W+1/Y7CntIiGV9rzTZ0IESH3HSUR/SfGnvlKNWfb3YiNF
VTM5G0wfjU88xJhrqNrmmnRvG1CfZpLI7mTsEsQSJ1DwO8lRO4qzvng1LUe3uu399RWzxPIFKT9/
e0+uh+BxaIiHt7DH3ylv7E4kEJ9IK5OtpnIH7eD/t2nrB4iMJYnf8SzQNAVAiFwHFo+AF50iU99H
kHxfJo/9r3IrZEhEXqIT6nudmYT4ddaiyg3D7MJu9/V02WJ1vdhIJY8vonKCvyOM7Zp4ZHZzVNdI
zhkAmbymi1xjh5Ov+u8Oz0koIFecE4GkIOPLXtNeGel54uigtBE4w2BHs0XfD6R9Ho3kXRMa7asF
uTZcn/Jguu+8zCaZernNHZwYlmcGNQvNqCXyyUcnz1iAfv30JGAf0AbLewOjspHaRUsivFxt83AB
YmSkSOXkgqmJTifOWBRjZv2JRnpwgt+6JIgnQEKdWyu2ZJirVm9ErC0kTXt7uA/2T7zO1yUxsVbG
6tMOrQcLoUFj7OuFyBZ6doclwsFTdO1GvBdyqwC5h7a1Il36h3DfsWgPH+cfi0ghfGSJOpxG4pJ0
7lA5VyKlygG6snl7WcqS82FD+KCg+smxxVL3u+Rf2GehORwIFyN/lHB76mnsupl981djZXm+lbs3
cLBVKGEK9CAdUmo/GWEcKYG9N9OusYsCf3Oz3rZsrnA8qAp0Z000Tub5mQ3Q8CGjfxQhfCN+V0W2
8VIHpFXDJxWN59WgGMoh9X+AcbrgKLfVFYroMMpJ1z8HUtcZTEiAIfc8hGdztnh2vZy3eDjQBiGm
BlTlGnkH2PhzaKmNI9G0wKXOClZgAP59zBMedp5TjcDFUywOamaiD/WeC+RTzJUrLsj55WdghMZF
Mpjef72QPvS2ii1mk4LBpg8OBWpKA1CdSnxNvZvHSlqVGdrb8XHuJhwfbUyIKdZSPSKYImQXK4OU
OY8EV8vB7BZ06j1ESoDGD8LW+FrYHJLUdfszMmG5gS+BB6ZU+LjOp3iXMhl2qcyQM4dkSupoia8D
nyDrrUIjkH3mEkoQT9vnke8/iWk8BlAASOFcCslsC58QZqKeDeFyamar63/VuvuTec8hcbXmz7gz
1TPqhjeIEcYWbwTO7mn4Cdk/vyVZHp4VMY8IXBh4xlYJHXjRZNqgdODfWbC8b501FzURhPuPArSM
PUnDitPrtRw1km5HzNkUY4WJIYXrAUIEar7m3i8G4Gx0UOZfGN94L1rcunWSso6gu+NvXVFHqIxE
2ndFVFm5gUGyDY/pUSCo+LIoz9pJFjX40vV6Rae6GpTxpozd3tdhhGI1rK8B099jRjr8DxfYOpXh
qtnMH1i1uzkn2SYmMNO+uprEQ9v+bz7bG7MFXuhtnoTkkaKGjgkCkPzd+0/N9B1PNJc5iO1EgEUw
wI6nDXK0YZMoBtey4lwOeW11A9ihBVKBZBjw4h19IgFmpuzBtApQ8rSDvPa40Moztl2b0lgYF37Q
PDMdyw2C+lj/1nvmj+myPqk3BKV4kOtBNgnlFa9/+N9aiC8RqOSAUjoibRr/WYZsfaQjOIdPDOSZ
FHlnoSheqytz//oWTXcL4SUjsW7FuBRR3VY0tlQzBFc7iXtTildIey5sFMtbQoqvJiHddpt6WjKf
kdRluC/Unps2234vSHLvje8yCt4yC7b2YeKn/hQi3HQhngzQOZchAUmZAz3GvobmfDByw1Nt9ifO
csQilWqQjffwKHWZojDBU+D+OeUGIhePZVjg0UVYGUcqD6YVHup24ppNW7a4nEIrSndLplbAN0xP
tnzLHD05WN8qgaIgxltBx0PjxSPZ/1316hs9YzTYJ1cHqF1g7yHVE9uIxeSD9DWS3Ek7fJZci9NE
gTV6bCSaR5LWm0hhL0KKexHRQCzpmatHV2TKhpY2gFnAPv0F88SHEQDksPnkBZoraD9RFvzbGk4o
kaw4cF+z/kW4w1W5uuJ6DhcKAqN8waQENqdSAqaJyosaa8Gb9dSXYILMwADPcXSSchNfX9CmzAKn
Wscfj9tET5s7N/8VpASvY8nwFW+hYak/lmNOGAEZhp/bZ8krZYMB/HfLepaJRlLiGjqzoyQy/6VN
UiftXFOftEXGVoi4D7rwnHiaTkexEo/h5eR1ENGvwZjyRj1oZbjRSoBVJBXmM6CnvVgv9JssP88X
eOlJ8REAwgpA0LhIQHx25LI9skhkyORSVa/LrgfGyvwEc6dJDFMM1DHH5Fka8vvysesLNwY8141G
OFt1vbd7TIetIjHCseWnuWPGO4fK8wzxDQiDpNKizKOtcwq7fewFY0DJvQwIFfLPyj0EBkFglBL7
JX7DL9Sg44NwUE0if/GUg9m9LksCAK2AZTo+GTwMS62Y46oOHYpTCxXIkSZ4Ojs9EnLTfPl+0swn
rmGKTA3xO8+/YnNNamXJ5JmLn/VCP3kLltF2RodY7XtxoZzfB4RWubBm2selzv7DRb6K/843zLB4
kAP7aYcPVIL3C9RDRZlRuJbopluBqMujR9BolTlBHP3WvQc8ZpfJr4n/9G8a+V1zEM38N/ukMFRy
X3Se5mvnca6ci4YjhjbY5pOZWyuePdstAG4V8Wr2xJflKSL+sVTywxCk1IdLiEIrbOUl55aotXnp
5Sxs0/F7nudn2JOOOCiDOOLLnDWUm8x5gbe3w8t7GSQkEh0/hbOugSis35kKyMToSvY/XOcnItw8
hJs1JqC2ncPBpaQ9yT1dRcSi7kqztPI0Hilylgvw9pcQ6chzbGBQpDcsBUOi76KVzqm2inIfmGNf
fYxHKgWHVVnWwdDuiw+7y7lX0FjcYrPKlOPV3R1TlVWH9bpBgvPqEaids4ilz6Urw5sEErIHF2pI
d5vjR1d4R6Z0BLoC5thD0HbkmHcQ5EtxZsvpPrNkYc7gYEiJ6Q5oElNiBk9nswQAE7C/1NVobSRe
7Yi1RT5tLumtzsJDCnjheD+jq169e3TW0cU/hHlJeQ1f5iSQsKndx1lkMlsaftWmX5NcgUjDxw3F
Utjvns9q6zjputfX9n4GmGAOy+sCkIQ1jutNnLcTi08r5Fl5XESkpTujfm/poDbv0bRp/m/mqVaP
D/2GvhdJagvZNKZMsac5Bkd1v3NW6uLbTi3LNs2W78+6cLTQED/sGaAakIL5QZULYXALdBDUWCcR
WoPT/JstxhKz12mv2ZAMyxHIIGQ8bZ53zgOk0oFZWVa4N9vjVSeLiVNpDEUbFhP4l0d7V6kcyYRc
8CyTgBTR8zY5KglEqlJTAYW1cnD6sQ5ctEBUEyMZ5lVj1o8F1/CmPKunTQsnniJ468g5iOpXXSlc
jHkM/Ah8YkpH/nd8po6mtuOcRAFwVame5TBLul7j11bHpjgfH2evwIlT49oQ/A+JMwUadK7vJoVB
m0k5+rrXuEMhexDD03BPZswIfX5BlwHolceA143FVxFQW5UqCCciu064CSwdRtYfG0OKaexx2h86
nwbqy/ArBgmlHBVPuij1aQA2qWk5G0yBNE+vBHR3kHxFDNyJ7Y/Ac8mEtwFH0F/lYaPreoyVo6UQ
GXwPAM4/GeBT6/6UoSBSdNkjd8HnITLsdBDnJeRZ1OUp93Txz2zOu5EqlJ/h+v++dohmf5nYwwkp
l4iRUT+5j0OAOD6DXELnd4d/PY1tkCzlos5gm68LZ1PbrRnM65Dg3ZnGVgVwASP0r5ol3IDSV5fU
pWBc9Tm51wWfvemTZvLGiiuIapK1XQskjxlO3JTesSccjae3buaU9W6vePSQYoXi/C+vIhM+XIMy
B0YYmJpNrqUlU7S1CdBBBQYYEpGvlicdMfHJBHUrHFw301v6b98NPpyGE91KQfui6WQGrCbcz3bF
Hls6vqpAEHhsMPERaqiA2PBQVNRLTyR4ebF9o1/fhahRiygAK9e68flWx+bBdcEMPAsl2Z2fFcbH
GpFmbEEEhkiHM29xa16mn+85tgfjhF5FoMSz9fJKaIxqgMNYg5UN19JgBah/MgQnE4PdL/004qBP
Ie7Z3UWHF2r5r4tWQVvcbUGR0XF0TEdHScKm9U7sgQH73+ixDWNvPn4Nn0yu4EjZMXEd4EclQxRa
vRVGcovK0ikl3ecdBVQwp31a+JJQQXSaQIAoxlQSMgmoRrtBf96f3dX3yynAJgYuMuj3/XUyWpJ5
hfGTuvtlhMuXBJVW9uVKXtcM4YljFjNqdJ0pmlvvBJiPrs+V3vxnnk5MAb8iyaZgMdkVxYCC+qPa
2+umJY+Qd4fM+BOhcuaNurBNx3yW3tkZeYVlBaXwotsNneWZRbe4aPBez5fqyYRn7N5qYTup4f9p
9j6RsbRmFHycHahNHIBvzXX8sxXNjdU9z3u169EQh8B27N25+oXawjV4DI1PZpUCeCmSM/Tg0u7N
tWNQ60jIyTWpvvcb0aGTD23uud4Yydfh4QURLp5qiqH6/JB7dIuEeWPYRRCMQVsjTduvmpMEX+d9
ifta8mnuruip2EkvNOmgKy23yMVrVf1WRqQHSsFIfJe0uh6M7blxnMoJGRoNBu/fBmkUYc4cCtID
36uNdnCTsFZxqMs1N1fziomMIDgtaN3DLzVXFB3AWpFaHMUL4p/Sl/g3Z0rYhMm8F9/8pqV+4wWZ
mr/b3sj7PQKmauLg6sqReWCTBmWsi8lZHm/RU8+n/fwGJndZgmCxjXPSHjjzqDlwxZRBnLUUuu6/
lpX7qht2duV9jUxGPwXYlt2fSwSvZTc+oTKAdUHAAr/IE9r0Nn/nGh8CRVUJgfsLslI3kwCYW3uY
zVaccZybq1c32M+v1b8rr6yv6C/evU4+USninEULtso9ljDjyzDRXilxWlRSX3ScJ+dFIg9Yc8DR
FTRmpOcOFtc/qExka3ktYCEyu3Rn2PpKfa+7yntTcwg0JUTVFmiWK53WEmisB6Ju9GNeAVfo2Y4U
ybIor9nXhH0iLd+LuTCNYyceXU3aBd0YdDxHpvEIe5STI3zoBxHn046/IibsSKC+0K4JbG7GCh4M
PCbHLZO7TPn95d9dLUcOefpb6l2yRroxrUBbYnfrNN7/MOUFvMkB44Y0rsExkldqZUn68/Vn2oGO
SnhqJMixa/pqiyPvQUTGuirfxwuGWWQxMP9Ntf23WFpitoU/bReGDGXd+jNFCMrp9+BVKSJId31L
RoyyAO/GHicaTgceAiWrVoG6JZFIBgpL1+wFpgILiE96H/EAVONqfX6Rnj10ZakY076wzmXXqIJj
VLsHTIrAtxQj+7aakTgXN0J8+8z5GmXYhcZA7OZE2Ttp3NGpWEcXx/6XywdlS0dd8IJVUY0ll0Jg
Sv8A43lqWm1WEnq0h4cm7n6lnhBEkeeq4i4it82GZ8Dwjk3bMPv/MvCfjHh/hUkKdcYNA6Nd8NPT
8KqnJh6kWiDW3yXl4Tx+ZIb7g3ncZg6d41qtFQNogVOLc49pkFVi7hXRe0bdzUO23JRu8oqDoXfa
9Yr5xuW83R6k7qXp1AKm8E+N0bS7X6TIKHaCvtlAGcGkelCbTN/6chwsbUuB1XV2pNCTZMSI3DUy
/as6nTZofsozI8IWpj7pBnKuPNtVgzBSNnfnfOICvpG5sLiksbXNoxsTQ62O6IiGgmJajfLDU3de
EEhiSXbgLyv9a3IZfUWA8owYvW4FaQ+AsapgiRIjz5Jj8nW89DI2PC/c1yR1xr/tqw0gcHHHVIBZ
9wxmR+9OlWBXg57z3A8qMshuf8xCwazt0aoOvuXSxQOjfsA6t7G5qKOwQrvHowBN/YjIJ0Pqedgo
/s/BRcD8i1o4NaugAYLvvkXKuU2pOR0nY/KAGsU9deRNLqQcYBxtQLS1o0dKK+BilxXKb+ua2tcI
A27lVfJnbKliofD+YU90DowGGuBTKpOm4fpsaHKr5+wRvF7oAg0NhbLtXGc6d2YMxFdVFJeenMIb
wWjPfjswRLZy7VmVud6TXUtAxqx4r1prgtN7AFYl0+TsFjScu8o+dik4of7Zl55V2lpFg2ApCUql
92DL/rltS3Pi1LvF+bOK/ZXTexGSgy0PW7MUagEZMPe2IKVgSm3YU2EnpS4DR4nhHg5/HZ2LXoYY
7m2EuqtzeoBP+PE1q8Q8kMHEr+vv6cCpN8l7eA93rbbJpiUKRpPmn/GduaLOUvnwXiFdc9e1jbLF
SYagmy9loJaZSpDPZTaIuKDeaVKlVJIWZh6miDT3fwUuSm8AogwaufDethMNAVN0kXKNtmmNfOlH
IxU0P7kfJrntnYNYb9fzpbjnAOStYJ3OQXHK7xC6ZuKpwz3E4cRygkuf2Qfv9A+efc1V787KKvIt
Seoph/NGYGy0Td6YRaeokNUIg4+jiycMAOMIFNOPNdINWKvDOvj9x86QUDwv70LYx/Ka4CdxiEk8
jQ+NJEM2mSGVK9AloKV0fcK/mGMux4LRZ3ysjsQr2V+zfCZDurGs/zqHDDuK/IOH89RCttgcoxGo
0LUP8gFe6W6RGIx+hTFRXmemV5xN/KtQuUwdIPp5pSqnG8yiEiIgxyzvnHDx6c/nu4ly45mcTzqX
shZXLcv/0hpcd6eg5WTSgqsFTiqEZSP2RasSaS9C17ljNm5Syo9YJMvI1t9ixiQXNQntk3WaJ3lP
/h7JJe0QF8LlZYQBsYbIWm1Nvdo+AkDivil3PYMSgShI2lcmpRcHx9Ah3O16QLhbFQMuu0j2eevI
qErnNPFcc5JFQOB1e+fRM7+Je8k1ZC8EaLcTMiBPbtz5CDOFiCO3pbtxQkIwaiUW67zLGgZJmk5L
2NAklgTxgaC+6j7O7dLEWZRIDJ26mtATZiozfMUakfquNX0UVQz+9kKDP20INmnCJbOYSOLmi/HJ
cqsGR8buFpY5djQJKWXxJcZ+r2F1Nk9StM3VI/9zpt+oAZeYj2tpxuZ1YHeLgIUd03dyMxpUZj6Z
jC2tLO1mJYoFoxZ46Qm9qKWMa7fuQVO98PBwc/rL/to1Ie3p3YWjqxGy5Y47FjQetKK6ukQ4lIet
sKQ+zAkIMgR6WA7E57o41VmA+FOqEf45rkNRUCX0h33PWsGrga5P53cypnrxCoQEZFENE8BP13sq
XeCGzWIW1xhOfBiDSzUUfFqy0Lz7ttHcvlrcKZkyZZxtoel0wXDWKT86opeopgq6gcSY3PKNcZc+
nwc4TTck18aR+EqTKOY5iqhxUD1lMILOeERuibL5idNWq/IR1EwDPXtn2BQCWk+t78iguxXJ5xlD
Ajxm3XYr+QJpp2GxqGHglxgW7Fx3TEyJQBIjiGeJ+B9mTX4FfI3iWPDg4hK+bFyJQus9/MIICnjo
iKxar3EZ/tMcTMZEm9wTm6nC33jmbJWNyokjnrKHWm13RMJ+yiNQN2P+phxE+WIekXZj21/Mscxn
C5u9KmDhGwLxyhjTeBNO7m2/UrqHmJTaooUqa5jpXG71rgDQX3HyPnQmNLvl+A+Wsx+Sdx2GuHU4
Uk+DPTXyob9ZPWjAkUGqwm3xAckCC71jUVBfEnMxap/QB9u55gXzbDvINtDK2J/E/gBoOlTIDi1j
wrhzIGF2Qt9PR9VN4FjUncUbc1arwskUCOarslb62xalvtAxBOYHQh+RbbzR/wT3CNNOXB1jdGcl
JcuwHab9GIM9ori5YZSdMSnXY3Bcqhj5rvnCFXC6y4PddRpi9DrUgS60RiE6cuGUiSX+gz8jK0oH
P0nXVDg1J6eP1x1VNEUwHFTNfWZIQqXqDGXVyfM1t38znQ00Q14v9vTOmQuBm8Qx2Ca8V6YdkEsq
KK6QzEEsy7QOHH3sfbnUdmL2MdZkhyJ61WkcJ+N80qxCojy/BQGJybiL8BsIHlAyQTNe2+BlJdyx
1wDwwkFm/mGn2lvX8VlX1Q8qsLFtcNh56mg6xCPov90T6l7oGrJEVwZ9SuutmpzpJ7ZJSHuz798c
e5iBN86FqjbqDxrQuYJIhK8pZMYxTF480/BbRrArd1UMV0Uvv8Dsts2/yWYSYiZQAIDrMEYbumr+
4wb5GfybP3IwWC4FUEalEqb/k1f88hE3lJBzR0Yk7rYwS9iG/8vyIouEY6SOIcQVVWGvN2DXBgKh
yQgaY3RUKFrt2GVPp3M7boJiO0s+Cy7fPP/fPVve0r3WQ3h1/wGwnPT/Htymo1VyLMwh4NC0lVcV
//c2A23bDdl5nW+4ZrQDDUagxAjr1bflbLyUIdCCRFiS+L/YqWnnyFXhWYzsC+mvdp2KyuKXRYa4
Z3MJwTgSm43mUxA+85UmSrP7M1dKkW9PbmScvKwyuGTG1eZqjV/Su0kYoQ3xUZm/K3Y7GMD/xVj6
hi3d0o55qTfVvg46uJgXY3vYZq9M/FyTvm5OwXLbiptdGhtGkUdsWSi/Uvlv+iFhQB+8d35Xwkgg
8DWNgshTUkxe+FOSsC065s6ewlK18N9fC7yvtg0jUqGXsF+E95zmBKHLAlfG5k1ZFKJk611S3kXq
HWQtFM+Pjmhj0smirFg6SRcPidPmxQY0J42zKKZrkMsnXSDode7tMaZerv16YlxaEnfkmylXbMwY
jqBZY4jFPH9YVLvMfsLPThGiiiD+DbhJtkcKE3EuFy17YdZj8OmckuqnIwm/7NVpzMb1h1W598wL
qtdcFPP1RjDWapy1BGk2u645DaDFGhB0LvwxLJUFW/C9QviwKQU7jVALQyrvdEdmkk0F7Je+Qv/j
8ypzEpPksJWX+9gfQ2h/r4mBSbOXWkL3XatEErxrmjfstdrPX6cKhxDXPYBkMZVQP3VQzDrbV6vB
gNbzLWnDkpkezEmOmA6Bp49g4izdfSxSTROIj3MHt30He7tPmvBiJa5IESU0KTpSWyVmI4MQaj28
1clWurBkC+fDVqtUx/bho3Hm+zVzOA0ublHc+yOUb9VrxW+YRaGVJKtGiH6M7aZhg86Wm1amelOS
YfvdZrA+4frGBiP6vVW72nQMSo12Ll89PfIDInzo+8b3xSkScigCKt5bPOVCqF6Vek9MgNQ+1ejq
3u60axMzyjXDW7eMcH8FgOEgbiw6KvUFAwbKO+89qOuyjBEK8/kCapET9/tkV394rDHL237A9nMr
EmPsJcPexMlcShHF4bZERhqX/MZ/dtrQLtPZLHqcm75DKeKPN1qgo5kjII6hmQwqM+SBlGreSr4l
QAF7C3qilx+Kzq64FsOlkDXjdjIdEpTcKiJG59CTp3Xgq9lla/1rYTP5gjvAvWZwKSekfiSXfUwL
nLVtHTVHqPUSeXAA09mgMJnQ5D30206sGghRVC8jDuBpGoFeyZadvL72w0TOKQ2LDPv/9ViXnqMu
hnyxU1mV/0TzEZ8wFRaic8tlBDsuyMA0frOHJ96MT3tzOLGP8VzYH6ifzAVOEVQnx6718cLTf2BW
b0DsVqCPVbT4szywCbHubg2mUvbuNppWMYhCHYSmJQwWdbSkTGnzo7T+dgJaLCKsb9A7bablOW/r
hM+32spqfFRupqZFZwv/L502lTnmK1mx8ATfQbZ0zI1qM2P0+/Mv/ExUn3gUBOK8N49YrUsLaKu5
Q6i5lzKKDldKIHcq14VWX4G8wzip92WB7S1qQIi76Mk3qy62T6+vgrfl5mj9Qo9OmRn+Lp0389zj
IZV3nW1c177yOcBnPEBV/cpMnX5d6A4bM1gyKbbAdGlwsDSw1lWQVbrH0qyfZmxgvxJI9rc2Nz59
nU7Y7qAY9bOH6Ie51Tkz+hZOKt+nhIHX9Ut7Ib+5JgAyUTdixjFTqvFK62kk1hkqstGK9SLek/lT
ohFBt26us/X6Ale/mUtmNaS+6ez0whvVo890S0uVguB1o+LHa5rulNkoZ27g1XYjYw8bvIruRXZh
hdRACyCC7eshA8lS0Em7SB8Xmwv+0BmNJB2w+q+XJfVhONNDuqY+8TwT9nerSfY7SwT/c4h0OaXt
KFB5st9wUa/PbnAg+f0Bwa2T4YMa7EswGd+5oZeQL0AsUv5w5/wuKuyN0Dor5BbzCl5RVY5r8Dwg
EIQ8TiGxHLyIqZr9TMZq2Ef7JQtlo8tmR4XfAi3Hoo+IQSLTWLDZuqtbBmkNPfBrax0qLBFLGn+1
ZDjbmh5RSVSwfxRi7fwqi1YI/5MPciF2q9gql9GKV3S0TnWsIA8i+4l0YvmNCHC/nlFXLpkEGMOT
VlAKJXoqUxr8OXl1IIszls3WDxwzy1b4mxQP3KIObtJdAW7Zr2MyPwrdP7QT6wvaI3VEbGiqkeZ2
XWXTlI6W6jc6d+Swv6RIxkR7E1H0cxnJRnITujFJtKdrRGXnWJx/aDTn0HgQMmI7yAAhLSjSwynS
A50SzhJfA2LCnibQkK6FPKjk0rspQgjPBRSlnn3pLRPBeC+CK7kSKd3JbJAZdL0nYZYoUMxpAQdo
5MU09U5LTcKa9XMTJygFUFtYDiSdsllKsM2Pm/HGsV0nqFNPWrdoi3c8XwtJH/HjqquZNumzlldX
O0hLVnASn0vxrK5M6V39Cy+LJYUme/TO/TaOM3pYTfpXlVJkUqIgvYyZ6m9fYzobBItzPiEcGtm4
kIbelna6PZ1cd5XDHetd4wNrdDmbwNVBqWo3Vr8dc/YikY+4/pE8f/SAuHkxN/UdMh4Sm8wHLDbZ
AIEl8hnxaJ9QxGO/sTMPDNHDQscMQJzNI6USZiz+Qto5KnLjVX0iEA4I+kXde/A5nN9pV48CVgiJ
Nz18OJAphKbn90MsqHd49U13StTqb7x01tXidblmjrkt3sIbfglyPRhSrCPGmcoiGfYj5c2UlttG
RlS05+CcQJT/l8y9wxLh7M7CdJbfJwiJMmpxKKCOrd3EsLPbMo7NOUlXx6875YxJZ6XK9e7buji1
lhwc4t9ISYQWNDZ6pgcs2nGZQgt3N550/8jVlA+3XHw+PrPEYDG29Iy7+S9PO2EqYdVN4nvmHxrg
5BeSR6xVm2yPf6aHbp9LCvCRcGv8A5jVcD5SBa2iAW8A7dz+GKO82fKhYK5Huln2PMkWicO/cTdu
f8tf4WRyTwAq3QPVb67Bu+MZVm4Yp4JsCWdfvfus5FoaoF9Wu9Xb3aE4m0IitZy4xDi4UC753LYh
p1EcaeAHjLmqdpUsgR1qFrh88nNKxjKGmSxGCoJ9N5FTfHFV8usr625pQm+IlrUwB2TtE/fuOeFq
TGHJVCELDWlE6Jvjn8YvuGux1mnhYPR53O+looe7SPldoL3d0eHijN/Uq5lr12uFpc1ZCJwgDtXk
Gf6tFnWLGMySseBd8Wg3xFQQ2o0QyVriYkAvT/JZTIS7Pjqy0VKb3+AdsTyygEfY6rddJ8oo4J24
jzP0aAka/5Do+fDvMcOxzcUkQpYNBCI2Zl4yIPzkbmKZFhfTDj0AIepykOCR85lbzD7e74H+oBqe
w5qyAxFE9Ed6o+CsLt3vdugmmLbvWBLWGlyZ7mQO27AEBTKKjvx9h/7bnfMQuzr6YSDgPMRMq2Ph
Ptgn6qfq4R0utk/2AfSBzmWXaVlgTKI1ORj4f5V9jExCUTqAgND/7N2pdVDlIX0v/nBpPp/gLclG
ReZDdbMnXQAWXXRKqcG7Y0J4njnSS8wzEjy5cfBXPYqudlrcS94eAJgVdd+jP8PQ+SEmv63H/yE4
skkeFmxftfkKjIkRbAtyoe9MT6sgyk6D7nYKMq5X7U5gxicZNrGKFLFB7kS4RuXouKP6Vq++7gP+
dYtBc8ufae2G9XpVHNJg6HxOJCueEzNjQt/o6El6VB8okzEp3yTHlKnKfdY8lkpKrnfEcTKS9IOV
MAi+8jwiZxGK/F0uQWPc4sAoIPupyHG2BTnfja82hJy2AuA7lSvH+krcaiLuBexISn1hRkzeb3zY
GRYx60EcdKHHqyqjTOP6ijcVRnS4vb9Ufows7AI/mNxH7puptzUVjSefS3by+1sLidoIoG5I359u
HM4crYfE7Z4sFkgwd6FYfIcm5EaFpqdP0GoBXGqOopNu4BlJTDYVdxi7Mue/kE7yrWV14xuGQvwO
FGbiLxXWmULhi7ZiGNvgCmBduW3WPeSGzuJm2HfkNMiIG4gLOmNHZHcCwozb1a4Mj2uN94Y1lD91
/NiYYRPemhhCfExaFBhyzZmo/3bZqI+gG6X2DyztIG+UYf7njylaZ/Fgg7F9BZt1E2mjZmKEvbOD
uMf9aLLxeVtFWBkyNkXiTAJ7rmVEcjpqJkPPy49jLOrGYKcxJeOBprGfvArP8mIE/BUR6tck7+Cv
5hY6eUFB79vBJtqMvwR+28DEa/JHpTV1ja4DhA8fUGKrNa9AUFqT9XwEArkk39960XQHNwieE+lU
I6vjBgou6U/Ky1nyHuQA2CL4vsHIG0vCn/w7k1LjAq5uPQ/Juutw9aqsSExZD7MTHs7DZRedkcWv
P9KLMqfdi/d+nelub6NCrGFu5deS52stJ38Nus5p58yLR0o4LSBu7ZMIHwYm2RKbfNP7ydEqPbxZ
POvd9V5JPsRgKHjUhelgW7XtvJUECeK8bVpFziEtoUX0GSz9lnJ+ilmfOCiTyvg7d4kT8/EpZozp
YOFli/wz4m1EOM7DTA8lkWoo9A9GgFVGBVoAlhV/ZAtv8738YYITEyi4EMDw5Np32U01Zuode2xN
6sI8hVv3HBWaj+xaj0fRlf3qyuCdoOKBHN5eIm55jJcy6U3Gwr+G95RI5LuWciWExih+U9MsxVht
SDz2JhL+6tzPm23InZUqwqUmCUNazLW6IR6B614dMXqVA8EHAU1rLUX3I0DJo8mGZhzcS6Q3lIOL
kxu2QGX59mhX47xzq594Kkxg1acpJh4zYYAwcEpWVKRbxhc1SO3Y7FzjBQj0UTvRkUI3e2MlN4pX
qpswYYnwmXlfCpSJOCvrdWctqWEW1o39TVFrTpuc8bfaxEQ3YR9QUQRf2q/syGDAXBxc0cNPEqnd
T/uSPNTV8wZo8hgp+ENbYktLq0MvHC/Yctav7Hn6DI9vojgaiEKEjZ26s1F5y2upS4r6Cs5Ufe3z
AgPHGqF9KoWpDQ6YPXw3jaG1QyY/x9ArkIqGR8J/W0Ut9cRSVDVrm/51NVe52OBA2oBrez9g8omH
QzZU0e0EWuAMZi+o4trn5/B5/90fuEkLPeB1CzCgZ8HeNvT/7AxHE/f1BCDTH+HIsspDpLmTJU1t
Fwy85FWFZUkUIYucPNNdu70ZuBX+9OK+tph6RJ+Aod34n5R1kUbq+7t4OLoQ70qx0whE2zhoqTxj
ZKSnRIA0CKoTCzD5FbnH9Sp4NZLP1tP52Ln86bFglc+k3SXuzCEiAOt7uRtxR69bZcWd2NkXkapk
y0a1zpm+lJp+xSWKSUz/wmmoo0fYr/tm3SvrvGvGvx9CWYuMkoR2uQfWHcXJRGEhJHV4xYlbYek2
cnhspKEbbc0ErXGY0PS/cj2f27pdFlwvi7nkx4KQsiScXYHY49vIhfLMy0HpMwZrv00fRG6yqfA6
bh8ETq1ax6OYDB4hehR9bJXR+sIM+8XkYjAeZWcduYd/KNHX41sjfkmEnzy9J9SsS0PcqSK49lCe
uUcP6+mxVcRPo+B6yyxzJnzPxh1yF66Z9d2tGwkXFZTB49gWNGyR4oLrYM74ob2hoMNHVH1Z7iM9
120qC7wp0CZDJvpVfIOMUlQ4x3STNtNDwm13qVsm3fIfaMYDHLlvWrFhEXCB0ps7SopKGd9aDvvt
dknIurLHUUvPEKp9bnO2zxAUW5MbSWCS/XiXLI4E9soxTc+11gjPawHjpM798kL4dUUj4BZmsKBG
AjNWA4Pql5AVficJ3qFm1UZ21TQNh6bwbPwThyglaNPlt99dPBZi9dxhdrv1+U3eOGyjD51AwQ0w
s27iEcPDqdO7LN42N/1KQfI/ZeHsdjsRmBKpujO7YNkfxpaOHHbnyL6m5WzbIrtQBmxdODDtAblH
Nh4Tpng5UysaAtSYXbD+b/49+y7EyATqoDs+OZ5I7tFor3D9vR4NIxpzMhfX1g7laVLoHq1ijRsI
ur+7eq+obppS++et6Bcyo/XbEyk22/OFWIPiYVVOAS1/1+V3l3XtyKxVyBQFfE2z3zwbBaY35wKS
3UFG3id/4aC8uK0+tAV6YMX/xuZwtHJ/u47cJu9ggsWrFwSBP/SLS/ILieowXFx6QKLv8IdK/+iA
3q5V5e7u/IHzm9KXw15KaFCTAU9fMXEIERWvmbgQ9TrrrqQqEQsa2kEVK/AH/zoCaykNVYzO7zRa
4I/FIhs6ehxCfzYM9WK+5OVifbjMG1cxQjVfUR8mDBF16n/7/oTJdK/KfatsTWhk2sOqMElTxmBP
NwSrOjuQIAK47b20+9xJAk+3u/SJiS9iXCHXdNI5GffUn2ZC25iTob2CLaYmyjWgk6h4YRJ1/xYC
SnUbOsLWPfKsb1zqxmq0pENQ/o9aZ04ckl8QZ76IAdsJmpfTNY/jIM3EqZI6OOa/SU57iPz28e1v
X0kDb8WS5r5wwjsSJlS12A/FrjSpp0dR7Y0nVfyRvddHJjvBuFavqJpUxS9qsXyjBRvXgqptsrtv
Qw81vohhEmntlu7EK4C20fmkafM0t5UMuLj1W7G68J/NTq+RfZuNZ551JRWsqBieB3V93lhsdkzU
eYkx0fizQVTpXtBKqq20qM2hC0yaunn3d8pxysKA3iPUNJeEApjkLYa1RLlyBMKh32aVOl2xGnVD
2YLEkpC90wgViaNDD+F3AygCBTd3W1VZRfQf9B/UZ8TW4KYnEwWD52H4AXVFyMdA++8NZk8WQgDn
nB6fhZwjXwNcJOltMmXiqYOS5NNzfTxBqeVnm5zLnyaBfaV+5hUN9U0+9wL38lRiP34hPIoNlJTO
uYoGWhgQl1Tt9oZGW9VgASeF5G5Z5UZNM31+gyjqP/NmRV7Ycmp1kIRdkPzsb8Tyq8Rmouz8guZf
TA4WmR8/ZxaNpQw5OJbJKqk4Qvgp27SLzYw5XEvfWHGMI4WXsGspeFV7uTUpM4xeeF5DmPaZWisN
kutCbw8O3Iz4OXLklmD8AotYeehJSd8FkAeHQO+TggxuYIOTN9FcA8TrxeyZMio2Ap9IRcxz0dcZ
qG/wkwA/rfUteip7hFDU/aJ3LSfA/KCkHZwVBoGR1YBkJGqGcDc7ao4rqM+76bNB4rHottu+Xdct
N0e9fNMOcuo/Jpx7o/68NrhxrReZ4DfUAOwCywI0jDdwdcXQmAoaq+cmDKKOeOenok1VBMv0Z+Ik
n2rf2HFxx63cvKGxKCLMi8/AcytTS05RRfFOvJObyPoRVX9WD0KDmFutrdJV/lE/BoITLUEj+VLK
IVOpa2ex9I1utt/WiqYf9iAA9aaeZ7DhUEUz78jA/ObPSeBl2niuwAroRJO596BSPQe62Ne4Ftnm
2IPCWFFvFRCcuBw4KfxbDbfr0GQem3vAvZkcC+r4aciBX8CuUAJGMnb907Jm4PghzhMigisD58Jh
SM57jjI8oHXGkyWZjzeBpACInop6XSdiyYea12dLKpIYdMklQsBGhfB9H5HQBqnckJEFYCrBdtHk
pWwQCTcXWexEJyL6DpFO4Trz294PF6PJmnKGZZ1ujWl9AN2nxcXttKVqczmCaOcOso/bpPwBXYL8
IN9Hwf3qrBSdBu+XfxOOGbNVeatiA+qtN3DCF4NWmHdNufUBWA7WjNPXSHMQUw7BG9hdfOn/9VpS
4xCed5U/ufrcOeIAEQQpccWk7KZfmkmP2m0g21ujkayi4goTfvU9Ewf7p7CoUSsdJYh3Wc9ls4R1
Kjba1IS8hpLA/LHW4X5Gxyqn6U/uv2+FMgBi2jlG1O0k6ZFxz0sngSOW+kijXa2hPJlrkRuEubzu
nFDiez5ekxDek68adxndhfHtqritPtRCDlvBbfo08wdVacHeo3/HSsSTM0+CoXQqNgHlPXMoXivC
qzQysNiQzWIOiAFJ9ERgQYuRU7QY8GP8hJKCriS3PbIp5c9Tb9i4oLGRLrJ8rnPc32MtXu0NCfIK
SlMon2MTuXfsrr9rVZ1UOE+r1VjoelmTSO/10gb1IaKP8NocjKLjfRpilWag6xJx/905UqOxPqmy
ynGckTHI3UAUF2I1snpPpfs7O8GlebfGgkzW1sPFmod9VmpTKAMbC1qBCAkGiCp2vHNlac7hVfr7
pwwUFQolDw+XPqqPbRYVImbC0iM/TsQ9VbWRIfG3XX993m1gJsVl6ZCD16rIKBw42JZaGEL89bUR
RAVcVSIw8SXG6GP5CpNvgUDGjYTjlKIx9BwC20hFK2NvW1qLjjIozAEqq7jomFos+8W7XuQ7LrWW
yJwgX9wOfbj1Wf2Rg7X89d5RNWO2sfGtdvsBx4ySo+S4KY9yj6K0wx8L4RPgNs0jnoz5rn/yeOWL
IBPZ4ZT5ARiLsl5+nPtjQ9LuBwfl/kDrfcM1N2xKR6MKQp5yPWqXkM6/+40fOmwvP95vm+oQ4N5p
RbQsoREfj0gOQvfCFopG/FBxU+nuKgvT4cXgvwStDMTdA67PkRIaoh9MeQGsdszaJoD1OZ5gWQIq
7yEp7MyRUMZly5pJpPcGx/hkZ7fASAiSyWpG+c6/gyaYS6+uMelAId8ugEWB8/jmzLKqw2XNcNO1
UopAAfDJIAIunYI6BEwauMHMM8uUEHgg9aCZjkMD4vAWB+SUbHEwo3YUmLjYec6tMHQwwvE6zCTr
BVEU5GPpYQQFehsdHDojVW9YrS1VJiD+VuAsbL0030/SCRpttmmkuGEXN9x+aJzKiMf+dMfIRHbm
uriqapTHkkUrIUOH3tRzjp5tI9E+gvMefEuiXPq2LCZQ/nQhkn2oYBsFJE6FIBD16hXa0IMi6wDv
GjAl3pgce5Lqid01JQ1W24fx01DTXEqkOzLKr0KfLyWlzwZ3sgG+neKBuok81/Hi8/sw/9xmFDZ1
QU+PbuQ4KYSp0h14V3Ub61fe6RSVFbZ2+Uee2AOFf0lolAu4Luh5o+ZFIRbPP+fLTyhG85VWukFL
s+DA1J1gwg7rW/UFoyvrZL1Q0JcM6QHOXuEUmRn9QVbNZNQHfpPcvmcsbYYuX8XBOGNAb8mG98s9
0KoDB2ezMxuqR2T+XmubGS299Pz850QBJOe0Fy8wyT26/wdmoNSwNWIj769F3THQ172903Kz2fQ6
RBi5kvM8L9RO8qvPWPhWRYMWEM3iGJJQc3fnIJUtjd1pTyYQ8iphX2fIDNiVHFiOMs9Fe6s+lqqV
NAbK3Y2kHY76vTnMfNPsI7LnD2VOl1APJ9WCNnTX7j8LIBKrIKyIxl72+rfDLktfSZzb6SpMSUO7
Raw2x8fWqOXnX2N8qWoqolEaW9lkXMA2McSRwJ86b8q2e1KEsaq1iwxuXTJ10831so89RArs7amg
VwV7TVXUoBOkKR25GG0R9A3zw4Z4wygxyjLCEOzstbVmaxudXxe2a3p4YuYEj7H0PKz37u6Ce3kJ
eKbPItdFvnrMWfckm0c7V6UTt8bFdNX5ezfdeGFzlC483jW3vf/FguMIVMgnLsClqT71OCmv6o4U
blZ48uDV/xs8bve1mOS3I5HwIXYUGX+XTz9eE9Ag7neGUjPNk9md/uIDrlgL8THxa2rPI+erDnhw
eFHwjn59RRXpc+ogPOqyUphXrnG87Q3JHIIR0wppDSCZ/oGKjDn0/egfCgn1NADAtZN4+pPzzlWF
ne+9bCW9vPXzdIVOngQ0rpWfrU81kbNMFC8cKevJzfNYObvNgQOTKKdN6D9oZn5v6vBckwwE7KvC
KwkHs95HU274UtZqsqFq9obPVcPmXb/Ji3imJ7+wBABD6LN+nTmhBuHodYPNZlkzKF6qwm4wzrOc
uhMXfkLsDxyonJZ02RCu8zrKJwwWyfm9aVfFrPnBwW7+4VngWCPua1jFE897mArlcpSY7av++fne
Z8GCjkq/uLlSHm5oHkPvpF5bfDcwv1sGNI2kvPFRyKlkmxMK9V1cQ2MkQ4vyuGhaxPcJG8UQ/m5+
9PNJJWltZmw4YO7lP8B+zIK2oLfY5/cDjKqC75RyOQd/l7X6Kt9Yos8q4IFKa2l3/zF1jWZoPHqG
eLTFXLG7FAF5kP//VyDetyoizPua5uOJJIRXU7E+KowwzpIVdFUfTt3Ocv18Bsjd8EOyQgPiNhJl
P0bhDNjIYB2bHth7E4J1dl6N/BFV/KrgXt5B57YQ7Vq9Q0erOOyIPxEzDNlNBiu93AQmySREbYWN
hrJrRAHAV2MPdKlslR3BdeWaK2MXgwiDpiRmIPc4TFAo9LECCQCvareqojVk8jwhJZirwEf5Q/tv
Ja82243SJ8ww/0e42I6iT+/ztIeTTPnLM087ZviGfftqOenJXNw56f2H2vFGthIao1PWWBLuJIxE
XKhYJ3ko4ZuPF4MYxcxXa+bXDvzQcZAAxUX9rA8E/Az5Kgb5ZbAYR0H/yQqu+uLPgyaY+OMDNVtN
76qpxBJZwPC5JzN+FViytEHvVa0Xv3YXD6aQlmgfoMNumiXx7NhbHyCtMeMdl75dT8drrSNLqkPP
O13BIvQcEvW+/mHT71CEiU8xQ8Rk9r7qPh1NPqk03XhuPAZPgyQaHU7INAiIH8caA5VGR3d88LRm
KW6e/dSnbl9XgsHvF667hXtAq9L/UNCCWNQTq3kHiZvVQvTtQFTZR+fvGkh7vK5+3SThTZ/NQzG/
3sGeJv2OqSERfmELQTKXfX07pyoPwNvz1rD5O2abhTnz4VW/8z9tHJm7uyWw8J2RFJUWbr1hd3iL
IH7QzsLbk99egnFHZI8hN2EEQBYZj1bg8GyAyFx763vaSWP/nZo6GjRfHFln5J5aGg2eFk3ha/vM
BdxpPvOtNhC3J9WkCLltKZddhj3/gqSgR+RhYrzsjJjMU7pAUO78YPYCQv4s3I2TL/8asAGxzhGx
02bHTMNCkh/DazPZppm58HQf7FRs9eYBu1gaV9uFDVlEfEfsXUEEYDu6LFmtEtokp8veEhlGfpIf
GQx3U6WLeH9D4C6ILOo1xnMoWYCc8baIVT9QZxAGOUfjq4kMSr5SUhTGkA2HoAbg7vc4MW9srvgD
VQsFmnlJceGDQpGqahTbEkhFs2mIBFwm0I3igiqZJfCzpu/O38c3ieDJdwN/P82lx9yk3Bm5dOz/
K5r6hmGbM5yvTgDJcypc5Zvcf8ZtdDLX1x3UvVZBRLFEg2p+3H3jgbdWqcAHDqoLZpCikGBH/R0O
6ZNqm6YzFJs6rgew5UvK4XvnEwxRorWYfvHm+lDUT9JC9MK8iGXs1IWbvz6GCgueA6CaRWTkUS1S
5O25QwNxlcTRvkWZJbl+cjbSTt98I3mpOpGCHadn0v4fWN/oXoxeCRbsDGQqCBKf/OSxp8imhbqv
O1olfCIrt6utjrnKITuiDBlRc8Whkksjmqpl2Aul+DUwLBM67gAvb4eIT5AyARIFEfskMcE+yONa
SR6i2qL0AIZfhPJ1voZ2KaXFbqI44VnlXlvVt3akZSriYUNSl6LuZSflhqJcTW+W2XFKEXeWHNLF
D8I9II1sRc/lEeON14cRXKvt822TQ7wrqEy+5yEXAPionTvsaHD7Q/94xTAsE306dDHjyWkXUbny
E0ORUlR4DqrOhTa3lEYXGWr+pB/uBCHW24xR8e5gUe/JyMaHXXn+Nh/nVEhGGhQcJZdfaEvdxQWC
AUzfbbxbRHsVoZEnBf22ZOcX4TBH0jn1nsGDwkZH5W2dcqMTvtOVuoKuH3havPhqcQ9w/4pd1bhw
ITsMVBBwywsM9zlqx2PE+ib8JiYs1im/Jxql/iH+oyQ11Aww9h25J/C12B7AX/CVZoccPF92MUc/
lKNIb35vaCXEjIL8cDXZ3jUuH5V1FRxdTfhiSIAvEpE1DibjwE3AyiaC91LUiIyTMSy8HZ2PNBVm
4WU8VK0hm+i3+EDAXvgF3Y84fm37RjbQ2N7sdJyTzEoBetasITWfPx/NJJAUBSQf/itdedetpZp6
lu2YBrTQ5m3OGNUuMC0THZh7dsYcP5u4VbUV7bproqAmH48BccBoAIYikgoskRJlT15FVKU+CGXX
w3UYI8P2aE5zHGXYLIAry4CnhdALRT4oDgKNwuOpVLtZo1H8+SS/9rHlroTYqzpDz4FO+8g0eODC
8qSMpvX0wPC2jMYpyFNTiaUXylkcJFo2ncFqrPvrImKaXMu4IMciPM6I6VhPfueCG9qzk5mwWMIZ
bOyAAVfzZUjgyYAKX7Saj2Hey7otgwav0Hv3m+veDgjhmPeqSFku/yp5qul1ppQzOaj5qAMFbcPp
aIQloF6NDGjsqkgHHWR4vbCHOD3YeuCK4KjbXaJ7tT1sU40FyuA18YGiNbIJrk12aPDJTgZumkk/
PqOzUTJYDvA0AOweBdiQMpfffOjN0sHzmewV1xJ8+Nwlr5ZInGwAeQ5SOGKaKi+VEYUXPhIohHzM
rpUVdr9qdFnh7NrEtc21LG0YVkUKxjc70pjWShkQZE0Jb6j5gAzoTwcFs0rZQgAL6Wje5Qr18vTN
W5hnb04jbT4vDwYOorlFRaNGmLU1dD9CUaXlsQFJhfE5lUd9Y+WD2WF3uWGlJ2qyiV7pWvRWvChy
PdKaD6tJSBqHoPX3aoQ93NMzpq9rO7bnsYnIwNtYDHPXfhXdM0BibTQY3Lu53s0X7kKt7xPpjDxD
cRkESYhVkLtcY7SHxp87COaca+CCttrd8ca5C/J51T+gLqJaHz7pHs1XsNlZ1ShHeoI293yrYnso
HfV1eGdFzuwzfzbjRWd0xseQZqysMicHsi8U1Xxe2Wcyivo83Ukc1/A3ylXcx/k9SK3lznO0C5bq
zUoEn9P5jh/tJYEI6eYMkBfx/C+Vtsn0NjdFGYMFuiW0/ohOcVfQfbIZC93/P/tmw3GPqeysofRl
93t/VNIw7V2G2q1Kg52IeFMA5uFB2djnTAZpVz47ayvMbjzqGUURfTi8SVTegMQyVWRpBLWMdRGM
BTSTehtHVm4hl+h878J+8RklfcR6Ba18A49eS2bpO3RzUtSjq/+i3YHIyN8e51RXCw4AHZnwBNSX
cKbrFawBvGab0UaM6F6lOLB7gyTL/bVqehROnXRY9pmxq8IDeogJm/MuJimZnTFUsdic4PycCqwQ
ZGyianqT0/NGXcvBUfGnhAKGtmLtYzNYj1nSsA/T+nPHkgEBETCROVQgoFtf+P/is2LNRb3Onwyy
KUwa/gmwDY6MLmcuxc33f/LMOA32pOMMK/OyA9mtQ+rwpMLzhKmIgngCsnD3HTULDxd4UE5B7nOV
j71MJ+4HTucw0Wdit0YyOjGre8sHGSXHRMgD/heoHi7r3YoRYDv5xXRgfj0aLMM5B5CDqW1mlW8w
3rUPm6M6za+NYL807JCY7phDDFmyeJTDA0iB8QmDyE5ZW9Rj6jj4TeoRVMoNJDJ5IwQJH2jJPyn7
LGSDPOKixkFD/XHK8wZtBVXdxLTUvPb8BcjtJJe3hEZw8jZdBcEZ4e63l7vTrpClsH4VbjkUXPft
H8Cg9tNq/y8iWHN0e5aUUsY9jOoNbIt4EuF6Xp8Bg4eEyZYC/wUw5iuzrZyollqedwrIWn8+JIiu
zIt1Mm0oVYyyMgnlhuY3o8CZ31aHzW+MCDB1v9bba4QANbIVrnxLWPZTsDltCsTpAXfjtrTKIT1l
WhTMlrv/0IGkQr7XQc82/Spdzd4Dgmd7jTRt/Leh35B8KNFP73F33XtzUs/+BMkzdVALDbtgNWrw
qhLtLZRGh8sH9JCk0TV6Fb8LuVAKOv2ucZ3Fj3hGif2hltZksYRK7rQLKT9Zlpwrfdl+scAAKkNl
f6p1zA4rglEVKOpKQklOGgd/zgYW+nyLndWbUs2nvoQ/clXsytlnC7tamQdUZlKdpDUVXORPmsTq
P7Q8nFm9hnBsMB6WUz0sosAiJ47sz97VNUVVfv9YiYIyguNZY7ljpHlPPcvhKC9CPPZCTKdJN5QZ
KHtoSkSoFfU96R8XBZrnGX/PtQjLzpX6wSq1GLxTq7AZTqt9/4tPxMlXKwd3zBE2A+gaiuT6Rxqi
8Hz4Qc0Zb7/rscmfoDlA5fcoRGXHE+WXXMCG4SU4JHtc1prcw6x35IRae1+BcvtjGfCwnYiPiA6j
o5bOfvONM2lnDuUM8bThO01UGy3wQugYd/o6tQuW4nbnEWbn1EmQ6a4gEuIsg5VJPYcn2vOJ7w8R
ZXHEvAnbne46zT4vmGKprxYq9ZL68OO2wzeYb7caZm1PZFlI3kw4Ds6y+AfJO82JhRdxqneMJdgD
+sYem1f2ynWwT+45g6RepdH/b9ExlkxFgwZ02dCVDJ8XLvv18etYDt0V9rO4OUL9rhnA1KVxGCUc
MlZBox9XQ/66bp4O8HC18QP/ZP32h6dDQUR7XKlZgjUgkSBgFEyzj/zybuMfbu8pxOF4k4WRIcLU
OoHYcjWfNKBW7W0JrFfU3o2+nUvO3KAM1R3DTjasF1+9RggGAyhJjDsbjipe8oJK1xYKRLPZmAKS
GtXFj/pKLmSZoRjbrNZzipfAkxad48L369DTt4/7vLiMRiu7NzqyvCmCXarXUbV8ww59snRGBIGn
AZ2/OFP/Q134ZXRVI8R5se8LK7kf9ixbHuVa+FUYz4GXxb6GE9hryUlsaIQSiCSZBBrwF2ouhaIZ
U4XrH0hzc8UoaZcwbZDK26Rw7eQ/OWLBP3a+SahvYs670zM06/I72GiUO85+IKCRE+Q4hDduayNe
q057We3+bnPhhsmrVYLoULzZC0lUGBRw1LEV3V8V7ZmFMbehJ4X/KHSdiQyw6k/UnF6tqsSAD8hB
D81edLVmMRancMzjeA8zUBbtqscO3gXhnAno5E56fchG8vl8XJ3yFMmj+oWFo4wIDAfPlUQKk/4w
jqHWN0LI4r+zokGtOTDRR9y4QPeEDeFueFHFpr6Arlr14y/PQRvlGwi2lqLYMle+UqaxMV862W80
3lS9rgPm7Bp90Hetr4Bcyfy3HzYX6SnNDIhtmtY4s25AHX6Hy2T2j/aeC8zce3xjjnuvDL2dsROB
KFIGWFU47w2tjOgIMQoeCGpvDT2IbFYPr2O2f/7nzzP93l66BKPg4zTFG0uHghAGoPKRmp8ilUC+
rcWCPvzWIp1A0M/YDcnB+q4HsRuR9BPtlSIsO775JGIduaEKCmeWCu8cgaWIQBTnAXvkZ0WCUso3
c1nT5TiBM7RpmPKNHbNHqsdEcv6ddQ8J3CS2N1TDTlKu+Hdf+cUB8rPO8UU8BujXmoGOBXKvPvUh
4NvMj6KzzA==
`protect end_protected

