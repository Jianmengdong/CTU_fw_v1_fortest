-------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 3.6
--  \   \         Application : 7 Series FPGAs Transceivers Wizard
--  /   /         Filename : gtwizard_0_multi_gt.vhd
-- /___/   /\     
-- \   \  /  \ 
--  \___\/\___\
--
--
-- Module gtwizard_0_multi_gt (a Multi GT Wrapper)
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;


--***************************** Entity Declaration ****************************

entity gtwizard_0_multi_gt is
generic
(

    -- Simulation attributes
    EXAMPLE_SIMULATION             : integer  := 0;      -- Set to 1 for simulation
    WRAPPER_SIM_GTRESET_SPEEDUP    : string   := "FALSE" -- Set to "TRUE" to speed up sim reset
);
port
(
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT0  (X0Y4)
    --____________________________CHANNEL PORTS________________________________
    GT0_DRP_BUSY_OUT                        : out  std_logic; 
 GT0_RXPMARESETDONE_OUT  : out  std_logic;
 GT0_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt0_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt0_drpclk_in                           : in   std_logic;
    gt0_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt0_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt0_drpen_in                            : in   std_logic;
    gt0_drprdy_out                          : out  std_logic;
    gt0_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt0_eyescanreset_in                     : in   std_logic;
    gt0_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt0_eyescandataerror_out                : out  std_logic;
    gt0_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt0_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt0_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt0_rxusrclk_in                         : in   std_logic;
    gt0_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt0_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt0_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt0_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt0_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt0_rxdlyen_in                          : in   std_logic;
    gt0_rxdlysreset_in                      : in   std_logic;
    gt0_rxdlysresetdone_out                 : out  std_logic;
    gt0_rxphalign_in                        : in   std_logic;
    gt0_rxphaligndone_out                   : out  std_logic;
    gt0_rxphalignen_in                      : in   std_logic;
    gt0_rxphdlyreset_in                     : in   std_logic;
    gt0_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt0_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    gt0_rxsyncallin_in                      : in   std_logic;
    gt0_rxsyncdone_out                      : out  std_logic;
    gt0_rxsyncin_in                         : in   std_logic;
    gt0_rxsyncmode_in                       : in   std_logic;
    gt0_rxsyncout_out                       : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt0_rxbyteisaligned_out                 : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt0_rxlpmhfhold_in                      : in   std_logic;
    gt0_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt0_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt0_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt0_rxoutclk_out                        : out  std_logic;
    gt0_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt0_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt0_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt0_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt0_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt0_gttxreset_in                        : in   std_logic;
    gt0_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt0_txusrclk_in                         : in   std_logic;
    gt0_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt0_txdlyen_in                          : in   std_logic;
    gt0_txdlysreset_in                      : in   std_logic;
    gt0_txdlysresetdone_out                 : out  std_logic;
    gt0_txphalign_in                        : in   std_logic;
    gt0_txphaligndone_out                   : out  std_logic;
    gt0_txphalignen_in                      : in   std_logic;
    gt0_txphdlyreset_in                     : in   std_logic;
    gt0_txphinit_in                         : in   std_logic;
    gt0_txphinitdone_out                    : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt0_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt0_gthtxn_out                          : out  std_logic;
    gt0_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt0_txoutclk_out                        : out  std_logic;
    gt0_txoutclkfabric_out                  : out  std_logic;
    gt0_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt0_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt0_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT1  (X0Y5)
    --____________________________CHANNEL PORTS________________________________
    GT1_DRP_BUSY_OUT                        : out  std_logic; 
 GT1_RXPMARESETDONE_OUT  : out  std_logic;
 GT1_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt1_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt1_drpclk_in                           : in   std_logic;
    gt1_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt1_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt1_drpen_in                            : in   std_logic;
    gt1_drprdy_out                          : out  std_logic;
    gt1_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt1_eyescanreset_in                     : in   std_logic;
    gt1_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt1_eyescandataerror_out                : out  std_logic;
    gt1_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt1_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt1_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt1_rxusrclk_in                         : in   std_logic;
    gt1_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt1_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt1_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt1_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt1_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt1_rxdlyen_in                          : in   std_logic;
    gt1_rxdlysreset_in                      : in   std_logic;
    gt1_rxdlysresetdone_out                 : out  std_logic;
    gt1_rxphalign_in                        : in   std_logic;
    gt1_rxphaligndone_out                   : out  std_logic;
    gt1_rxphalignen_in                      : in   std_logic;
    gt1_rxphdlyreset_in                     : in   std_logic;
    gt1_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt1_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    gt1_rxsyncallin_in                      : in   std_logic;
    gt1_rxsyncdone_out                      : out  std_logic;
    gt1_rxsyncin_in                         : in   std_logic;
    gt1_rxsyncmode_in                       : in   std_logic;
    gt1_rxsyncout_out                       : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt1_rxbyteisaligned_out                 : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt1_rxlpmhfhold_in                      : in   std_logic;
    gt1_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt1_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt1_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt1_rxoutclk_out                        : out  std_logic;
    gt1_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt1_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt1_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt1_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt1_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt1_gttxreset_in                        : in   std_logic;
    gt1_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt1_txusrclk_in                         : in   std_logic;
    gt1_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt1_txdlyen_in                          : in   std_logic;
    gt1_txdlysreset_in                      : in   std_logic;
    gt1_txdlysresetdone_out                 : out  std_logic;
    gt1_txphalign_in                        : in   std_logic;
    gt1_txphaligndone_out                   : out  std_logic;
    gt1_txphalignen_in                      : in   std_logic;
    gt1_txphdlyreset_in                     : in   std_logic;
    gt1_txphinit_in                         : in   std_logic;
    gt1_txphinitdone_out                    : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt1_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt1_gthtxn_out                          : out  std_logic;
    gt1_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt1_txoutclk_out                        : out  std_logic;
    gt1_txoutclkfabric_out                  : out  std_logic;
    gt1_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt1_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt1_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT2  (X0Y6)
    --____________________________CHANNEL PORTS________________________________
    GT2_DRP_BUSY_OUT                        : out  std_logic; 
 GT2_RXPMARESETDONE_OUT  : out  std_logic;
 GT2_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt2_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt2_drpclk_in                           : in   std_logic;
    gt2_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt2_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt2_drpen_in                            : in   std_logic;
    gt2_drprdy_out                          : out  std_logic;
    gt2_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt2_eyescanreset_in                     : in   std_logic;
    gt2_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt2_eyescandataerror_out                : out  std_logic;
    gt2_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt2_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt2_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt2_rxusrclk_in                         : in   std_logic;
    gt2_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt2_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt2_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt2_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt2_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt2_rxdlyen_in                          : in   std_logic;
    gt2_rxdlysreset_in                      : in   std_logic;
    gt2_rxdlysresetdone_out                 : out  std_logic;
    gt2_rxphalign_in                        : in   std_logic;
    gt2_rxphaligndone_out                   : out  std_logic;
    gt2_rxphalignen_in                      : in   std_logic;
    gt2_rxphdlyreset_in                     : in   std_logic;
    gt2_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt2_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    gt2_rxsyncallin_in                      : in   std_logic;
    gt2_rxsyncdone_out                      : out  std_logic;
    gt2_rxsyncin_in                         : in   std_logic;
    gt2_rxsyncmode_in                       : in   std_logic;
    gt2_rxsyncout_out                       : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt2_rxbyteisaligned_out                 : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt2_rxlpmhfhold_in                      : in   std_logic;
    gt2_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt2_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt2_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt2_rxoutclk_out                        : out  std_logic;
    gt2_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt2_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt2_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt2_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt2_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt2_gttxreset_in                        : in   std_logic;
    gt2_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt2_txusrclk_in                         : in   std_logic;
    gt2_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt2_txdlyen_in                          : in   std_logic;
    gt2_txdlysreset_in                      : in   std_logic;
    gt2_txdlysresetdone_out                 : out  std_logic;
    gt2_txphalign_in                        : in   std_logic;
    gt2_txphaligndone_out                   : out  std_logic;
    gt2_txphalignen_in                      : in   std_logic;
    gt2_txphdlyreset_in                     : in   std_logic;
    gt2_txphinit_in                         : in   std_logic;
    gt2_txphinitdone_out                    : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt2_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt2_gthtxn_out                          : out  std_logic;
    gt2_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt2_txoutclk_out                        : out  std_logic;
    gt2_txoutclkfabric_out                  : out  std_logic;
    gt2_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt2_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt2_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT3  (X0Y7)
    --____________________________CHANNEL PORTS________________________________
    GT3_DRP_BUSY_OUT                        : out  std_logic; 
 GT3_RXPMARESETDONE_OUT  : out  std_logic;
 GT3_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt3_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt3_drpclk_in                           : in   std_logic;
    gt3_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt3_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt3_drpen_in                            : in   std_logic;
    gt3_drprdy_out                          : out  std_logic;
    gt3_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt3_eyescanreset_in                     : in   std_logic;
    gt3_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt3_eyescandataerror_out                : out  std_logic;
    gt3_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt3_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt3_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt3_rxusrclk_in                         : in   std_logic;
    gt3_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt3_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt3_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt3_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt3_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt3_rxdlyen_in                          : in   std_logic;
    gt3_rxdlysreset_in                      : in   std_logic;
    gt3_rxdlysresetdone_out                 : out  std_logic;
    gt3_rxphalign_in                        : in   std_logic;
    gt3_rxphaligndone_out                   : out  std_logic;
    gt3_rxphalignen_in                      : in   std_logic;
    gt3_rxphdlyreset_in                     : in   std_logic;
    gt3_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt3_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    gt3_rxsyncallin_in                      : in   std_logic;
    gt3_rxsyncdone_out                      : out  std_logic;
    gt3_rxsyncin_in                         : in   std_logic;
    gt3_rxsyncmode_in                       : in   std_logic;
    gt3_rxsyncout_out                       : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt3_rxbyteisaligned_out                 : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt3_rxlpmhfhold_in                      : in   std_logic;
    gt3_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt3_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt3_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt3_rxoutclk_out                        : out  std_logic;
    gt3_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt3_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt3_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt3_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt3_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt3_gttxreset_in                        : in   std_logic;
    gt3_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt3_txusrclk_in                         : in   std_logic;
    gt3_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt3_txdlyen_in                          : in   std_logic;
    gt3_txdlysreset_in                      : in   std_logic;
    gt3_txdlysresetdone_out                 : out  std_logic;
    gt3_txphalign_in                        : in   std_logic;
    gt3_txphaligndone_out                   : out  std_logic;
    gt3_txphalignen_in                      : in   std_logic;
    gt3_txphdlyreset_in                     : in   std_logic;
    gt3_txphinit_in                         : in   std_logic;
    gt3_txphinitdone_out                    : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt3_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt3_gthtxn_out                          : out  std_logic;
    gt3_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt3_txoutclk_out                        : out  std_logic;
    gt3_txoutclkfabric_out                  : out  std_logic;
    gt3_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt3_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt3_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT4  (X0Y8)
    --____________________________CHANNEL PORTS________________________________
    GT4_DRP_BUSY_OUT                        : out  std_logic; 
 GT4_RXPMARESETDONE_OUT  : out  std_logic;
 GT4_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt4_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt4_drpclk_in                           : in   std_logic;
    gt4_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt4_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt4_drpen_in                            : in   std_logic;
    gt4_drprdy_out                          : out  std_logic;
    gt4_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt4_eyescanreset_in                     : in   std_logic;
    gt4_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt4_eyescandataerror_out                : out  std_logic;
    gt4_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt4_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt4_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt4_rxusrclk_in                         : in   std_logic;
    gt4_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt4_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt4_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt4_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt4_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt4_rxdlyen_in                          : in   std_logic;
    gt4_rxdlysreset_in                      : in   std_logic;
    gt4_rxdlysresetdone_out                 : out  std_logic;
    gt4_rxphalign_in                        : in   std_logic;
    gt4_rxphaligndone_out                   : out  std_logic;
    gt4_rxphalignen_in                      : in   std_logic;
    gt4_rxphdlyreset_in                     : in   std_logic;
    gt4_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt4_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    gt4_rxsyncallin_in                      : in   std_logic;
    gt4_rxsyncdone_out                      : out  std_logic;
    gt4_rxsyncin_in                         : in   std_logic;
    gt4_rxsyncmode_in                       : in   std_logic;
    gt4_rxsyncout_out                       : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt4_rxbyteisaligned_out                 : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt4_rxlpmhfhold_in                      : in   std_logic;
    gt4_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt4_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt4_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt4_rxoutclk_out                        : out  std_logic;
    gt4_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt4_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt4_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt4_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt4_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt4_gttxreset_in                        : in   std_logic;
    gt4_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt4_txusrclk_in                         : in   std_logic;
    gt4_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt4_txdlyen_in                          : in   std_logic;
    gt4_txdlysreset_in                      : in   std_logic;
    gt4_txdlysresetdone_out                 : out  std_logic;
    gt4_txphalign_in                        : in   std_logic;
    gt4_txphaligndone_out                   : out  std_logic;
    gt4_txphalignen_in                      : in   std_logic;
    gt4_txphdlyreset_in                     : in   std_logic;
    gt4_txphinit_in                         : in   std_logic;
    gt4_txphinitdone_out                    : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt4_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt4_gthtxn_out                          : out  std_logic;
    gt4_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt4_txoutclk_out                        : out  std_logic;
    gt4_txoutclkfabric_out                  : out  std_logic;
    gt4_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt4_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt4_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT5  (X0Y9)
    --____________________________CHANNEL PORTS________________________________
    GT5_DRP_BUSY_OUT                        : out  std_logic; 
 GT5_RXPMARESETDONE_OUT  : out  std_logic;
 GT5_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt5_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt5_drpclk_in                           : in   std_logic;
    gt5_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt5_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt5_drpen_in                            : in   std_logic;
    gt5_drprdy_out                          : out  std_logic;
    gt5_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt5_eyescanreset_in                     : in   std_logic;
    gt5_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt5_eyescandataerror_out                : out  std_logic;
    gt5_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt5_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt5_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt5_rxusrclk_in                         : in   std_logic;
    gt5_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt5_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt5_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt5_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt5_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt5_rxdlyen_in                          : in   std_logic;
    gt5_rxdlysreset_in                      : in   std_logic;
    gt5_rxdlysresetdone_out                 : out  std_logic;
    gt5_rxphalign_in                        : in   std_logic;
    gt5_rxphaligndone_out                   : out  std_logic;
    gt5_rxphalignen_in                      : in   std_logic;
    gt5_rxphdlyreset_in                     : in   std_logic;
    gt5_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt5_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    gt5_rxsyncallin_in                      : in   std_logic;
    gt5_rxsyncdone_out                      : out  std_logic;
    gt5_rxsyncin_in                         : in   std_logic;
    gt5_rxsyncmode_in                       : in   std_logic;
    gt5_rxsyncout_out                       : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt5_rxbyteisaligned_out                 : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt5_rxlpmhfhold_in                      : in   std_logic;
    gt5_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt5_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt5_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt5_rxoutclk_out                        : out  std_logic;
    gt5_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt5_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt5_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt5_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt5_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt5_gttxreset_in                        : in   std_logic;
    gt5_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt5_txusrclk_in                         : in   std_logic;
    gt5_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt5_txdlyen_in                          : in   std_logic;
    gt5_txdlysreset_in                      : in   std_logic;
    gt5_txdlysresetdone_out                 : out  std_logic;
    gt5_txphalign_in                        : in   std_logic;
    gt5_txphaligndone_out                   : out  std_logic;
    gt5_txphalignen_in                      : in   std_logic;
    gt5_txphdlyreset_in                     : in   std_logic;
    gt5_txphinit_in                         : in   std_logic;
    gt5_txphinitdone_out                    : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt5_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt5_gthtxn_out                          : out  std_logic;
    gt5_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt5_txoutclk_out                        : out  std_logic;
    gt5_txoutclkfabric_out                  : out  std_logic;
    gt5_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt5_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt5_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT6  (X0Y10)
    --____________________________CHANNEL PORTS________________________________
    GT6_DRP_BUSY_OUT                        : out  std_logic; 
 GT6_RXPMARESETDONE_OUT  : out  std_logic;
 GT6_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt6_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt6_drpclk_in                           : in   std_logic;
    gt6_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt6_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt6_drpen_in                            : in   std_logic;
    gt6_drprdy_out                          : out  std_logic;
    gt6_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt6_eyescanreset_in                     : in   std_logic;
    gt6_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt6_eyescandataerror_out                : out  std_logic;
    gt6_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt6_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt6_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt6_rxusrclk_in                         : in   std_logic;
    gt6_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt6_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt6_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt6_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt6_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt6_rxdlyen_in                          : in   std_logic;
    gt6_rxdlysreset_in                      : in   std_logic;
    gt6_rxdlysresetdone_out                 : out  std_logic;
    gt6_rxphalign_in                        : in   std_logic;
    gt6_rxphaligndone_out                   : out  std_logic;
    gt6_rxphalignen_in                      : in   std_logic;
    gt6_rxphdlyreset_in                     : in   std_logic;
    gt6_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt6_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    gt6_rxsyncallin_in                      : in   std_logic;
    gt6_rxsyncdone_out                      : out  std_logic;
    gt6_rxsyncin_in                         : in   std_logic;
    gt6_rxsyncmode_in                       : in   std_logic;
    gt6_rxsyncout_out                       : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt6_rxbyteisaligned_out                 : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt6_rxlpmhfhold_in                      : in   std_logic;
    gt6_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt6_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt6_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt6_rxoutclk_out                        : out  std_logic;
    gt6_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt6_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt6_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt6_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt6_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt6_gttxreset_in                        : in   std_logic;
    gt6_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt6_txusrclk_in                         : in   std_logic;
    gt6_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt6_txdlyen_in                          : in   std_logic;
    gt6_txdlysreset_in                      : in   std_logic;
    gt6_txdlysresetdone_out                 : out  std_logic;
    gt6_txphalign_in                        : in   std_logic;
    gt6_txphaligndone_out                   : out  std_logic;
    gt6_txphalignen_in                      : in   std_logic;
    gt6_txphdlyreset_in                     : in   std_logic;
    gt6_txphinit_in                         : in   std_logic;
    gt6_txphinitdone_out                    : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt6_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt6_gthtxn_out                          : out  std_logic;
    gt6_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt6_txoutclk_out                        : out  std_logic;
    gt6_txoutclkfabric_out                  : out  std_logic;
    gt6_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt6_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt6_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT7  (X0Y11)
    --____________________________CHANNEL PORTS________________________________
    GT7_DRP_BUSY_OUT                        : out  std_logic; 
 GT7_RXPMARESETDONE_OUT  : out  std_logic;
 GT7_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt7_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt7_drpclk_in                           : in   std_logic;
    gt7_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt7_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt7_drpen_in                            : in   std_logic;
    gt7_drprdy_out                          : out  std_logic;
    gt7_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt7_eyescanreset_in                     : in   std_logic;
    gt7_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt7_eyescandataerror_out                : out  std_logic;
    gt7_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt7_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt7_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt7_rxusrclk_in                         : in   std_logic;
    gt7_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt7_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt7_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt7_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt7_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt7_rxdlyen_in                          : in   std_logic;
    gt7_rxdlysreset_in                      : in   std_logic;
    gt7_rxdlysresetdone_out                 : out  std_logic;
    gt7_rxphalign_in                        : in   std_logic;
    gt7_rxphaligndone_out                   : out  std_logic;
    gt7_rxphalignen_in                      : in   std_logic;
    gt7_rxphdlyreset_in                     : in   std_logic;
    gt7_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt7_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    gt7_rxsyncallin_in                      : in   std_logic;
    gt7_rxsyncdone_out                      : out  std_logic;
    gt7_rxsyncin_in                         : in   std_logic;
    gt7_rxsyncmode_in                       : in   std_logic;
    gt7_rxsyncout_out                       : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt7_rxbyteisaligned_out                 : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt7_rxlpmhfhold_in                      : in   std_logic;
    gt7_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt7_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt7_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt7_rxoutclk_out                        : out  std_logic;
    gt7_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt7_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt7_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt7_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt7_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt7_gttxreset_in                        : in   std_logic;
    gt7_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt7_txusrclk_in                         : in   std_logic;
    gt7_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt7_txdlyen_in                          : in   std_logic;
    gt7_txdlysreset_in                      : in   std_logic;
    gt7_txdlysresetdone_out                 : out  std_logic;
    gt7_txphalign_in                        : in   std_logic;
    gt7_txphaligndone_out                   : out  std_logic;
    gt7_txphalignen_in                      : in   std_logic;
    gt7_txphdlyreset_in                     : in   std_logic;
    gt7_txphinit_in                         : in   std_logic;
    gt7_txphinitdone_out                    : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt7_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt7_gthtxn_out                          : out  std_logic;
    gt7_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt7_txoutclk_out                        : out  std_logic;
    gt7_txoutclkfabric_out                  : out  std_logic;
    gt7_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt7_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt7_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT8  (X0Y12)
    --____________________________CHANNEL PORTS________________________________
    GT8_DRP_BUSY_OUT                        : out  std_logic; 
 GT8_RXPMARESETDONE_OUT  : out  std_logic;
 GT8_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt8_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt8_drpclk_in                           : in   std_logic;
    gt8_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt8_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt8_drpen_in                            : in   std_logic;
    gt8_drprdy_out                          : out  std_logic;
    gt8_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt8_eyescanreset_in                     : in   std_logic;
    gt8_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt8_eyescandataerror_out                : out  std_logic;
    gt8_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt8_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt8_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt8_rxusrclk_in                         : in   std_logic;
    gt8_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt8_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt8_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt8_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt8_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt8_rxdlyen_in                          : in   std_logic;
    gt8_rxdlysreset_in                      : in   std_logic;
    gt8_rxdlysresetdone_out                 : out  std_logic;
    gt8_rxphalign_in                        : in   std_logic;
    gt8_rxphaligndone_out                   : out  std_logic;
    gt8_rxphalignen_in                      : in   std_logic;
    gt8_rxphdlyreset_in                     : in   std_logic;
    gt8_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt8_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    gt8_rxsyncallin_in                      : in   std_logic;
    gt8_rxsyncdone_out                      : out  std_logic;
    gt8_rxsyncin_in                         : in   std_logic;
    gt8_rxsyncmode_in                       : in   std_logic;
    gt8_rxsyncout_out                       : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt8_rxbyteisaligned_out                 : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt8_rxlpmhfhold_in                      : in   std_logic;
    gt8_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt8_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt8_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt8_rxoutclk_out                        : out  std_logic;
    gt8_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt8_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt8_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt8_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt8_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt8_gttxreset_in                        : in   std_logic;
    gt8_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt8_txusrclk_in                         : in   std_logic;
    gt8_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt8_txdlyen_in                          : in   std_logic;
    gt8_txdlysreset_in                      : in   std_logic;
    gt8_txdlysresetdone_out                 : out  std_logic;
    gt8_txphalign_in                        : in   std_logic;
    gt8_txphaligndone_out                   : out  std_logic;
    gt8_txphalignen_in                      : in   std_logic;
    gt8_txphdlyreset_in                     : in   std_logic;
    gt8_txphinit_in                         : in   std_logic;
    gt8_txphinitdone_out                    : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt8_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt8_gthtxn_out                          : out  std_logic;
    gt8_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt8_txoutclk_out                        : out  std_logic;
    gt8_txoutclkfabric_out                  : out  std_logic;
    gt8_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt8_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt8_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT9  (X0Y13)
    --____________________________CHANNEL PORTS________________________________
    GT9_DRP_BUSY_OUT                        : out  std_logic; 
 GT9_RXPMARESETDONE_OUT  : out  std_logic;
 GT9_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt9_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt9_drpclk_in                           : in   std_logic;
    gt9_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt9_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt9_drpen_in                            : in   std_logic;
    gt9_drprdy_out                          : out  std_logic;
    gt9_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt9_eyescanreset_in                     : in   std_logic;
    gt9_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt9_eyescandataerror_out                : out  std_logic;
    gt9_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt9_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt9_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt9_rxusrclk_in                         : in   std_logic;
    gt9_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt9_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt9_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt9_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt9_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt9_rxdlyen_in                          : in   std_logic;
    gt9_rxdlysreset_in                      : in   std_logic;
    gt9_rxdlysresetdone_out                 : out  std_logic;
    gt9_rxphalign_in                        : in   std_logic;
    gt9_rxphaligndone_out                   : out  std_logic;
    gt9_rxphalignen_in                      : in   std_logic;
    gt9_rxphdlyreset_in                     : in   std_logic;
    gt9_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt9_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    gt9_rxsyncallin_in                      : in   std_logic;
    gt9_rxsyncdone_out                      : out  std_logic;
    gt9_rxsyncin_in                         : in   std_logic;
    gt9_rxsyncmode_in                       : in   std_logic;
    gt9_rxsyncout_out                       : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt9_rxbyteisaligned_out                 : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt9_rxlpmhfhold_in                      : in   std_logic;
    gt9_rxlpmlfhold_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt9_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt9_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt9_rxoutclk_out                        : out  std_logic;
    gt9_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt9_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt9_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt9_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt9_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt9_gttxreset_in                        : in   std_logic;
    gt9_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt9_txusrclk_in                         : in   std_logic;
    gt9_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt9_txdlyen_in                          : in   std_logic;
    gt9_txdlysreset_in                      : in   std_logic;
    gt9_txdlysresetdone_out                 : out  std_logic;
    gt9_txphalign_in                        : in   std_logic;
    gt9_txphaligndone_out                   : out  std_logic;
    gt9_txphalignen_in                      : in   std_logic;
    gt9_txphdlyreset_in                     : in   std_logic;
    gt9_txphinit_in                         : in   std_logic;
    gt9_txphinitdone_out                    : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt9_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt9_gthtxn_out                          : out  std_logic;
    gt9_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt9_txoutclk_out                        : out  std_logic;
    gt9_txoutclkfabric_out                  : out  std_logic;
    gt9_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt9_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt9_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT10  (X0Y14)
    --____________________________CHANNEL PORTS________________________________
    GT10_DRP_BUSY_OUT                        : out  std_logic; 
 GT10_RXPMARESETDONE_OUT  : out  std_logic;
 GT10_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt10_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt10_drpclk_in                          : in   std_logic;
    gt10_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt10_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt10_drpen_in                           : in   std_logic;
    gt10_drprdy_out                         : out  std_logic;
    gt10_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt10_eyescanreset_in                    : in   std_logic;
    gt10_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt10_eyescandataerror_out               : out  std_logic;
    gt10_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt10_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt10_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt10_rxusrclk_in                        : in   std_logic;
    gt10_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt10_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt10_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt10_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt10_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt10_rxdlyen_in                         : in   std_logic;
    gt10_rxdlysreset_in                     : in   std_logic;
    gt10_rxdlysresetdone_out                : out  std_logic;
    gt10_rxphalign_in                       : in   std_logic;
    gt10_rxphaligndone_out                  : out  std_logic;
    gt10_rxphalignen_in                     : in   std_logic;
    gt10_rxphdlyreset_in                    : in   std_logic;
    gt10_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt10_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt10_rxsyncallin_in                     : in   std_logic;
    gt10_rxsyncdone_out                     : out  std_logic;
    gt10_rxsyncin_in                        : in   std_logic;
    gt10_rxsyncmode_in                      : in   std_logic;
    gt10_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt10_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt10_rxlpmhfhold_in                     : in   std_logic;
    gt10_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt10_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt10_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt10_rxoutclk_out                       : out  std_logic;
    gt10_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt10_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt10_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt10_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt10_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt10_gttxreset_in                       : in   std_logic;
    gt10_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt10_txusrclk_in                        : in   std_logic;
    gt10_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt10_txdlyen_in                         : in   std_logic;
    gt10_txdlysreset_in                     : in   std_logic;
    gt10_txdlysresetdone_out                : out  std_logic;
    gt10_txphalign_in                       : in   std_logic;
    gt10_txphaligndone_out                  : out  std_logic;
    gt10_txphalignen_in                     : in   std_logic;
    gt10_txphdlyreset_in                    : in   std_logic;
    gt10_txphinit_in                        : in   std_logic;
    gt10_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt10_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt10_gthtxn_out                         : out  std_logic;
    gt10_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt10_txoutclk_out                       : out  std_logic;
    gt10_txoutclkfabric_out                 : out  std_logic;
    gt10_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt10_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt10_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT11  (X0Y15)
    --____________________________CHANNEL PORTS________________________________
    GT11_DRP_BUSY_OUT                        : out  std_logic; 
 GT11_RXPMARESETDONE_OUT  : out  std_logic;
 GT11_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt11_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt11_drpclk_in                          : in   std_logic;
    gt11_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt11_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt11_drpen_in                           : in   std_logic;
    gt11_drprdy_out                         : out  std_logic;
    gt11_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt11_eyescanreset_in                    : in   std_logic;
    gt11_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt11_eyescandataerror_out               : out  std_logic;
    gt11_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt11_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt11_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt11_rxusrclk_in                        : in   std_logic;
    gt11_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt11_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt11_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt11_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt11_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt11_rxdlyen_in                         : in   std_logic;
    gt11_rxdlysreset_in                     : in   std_logic;
    gt11_rxdlysresetdone_out                : out  std_logic;
    gt11_rxphalign_in                       : in   std_logic;
    gt11_rxphaligndone_out                  : out  std_logic;
    gt11_rxphalignen_in                     : in   std_logic;
    gt11_rxphdlyreset_in                    : in   std_logic;
    gt11_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt11_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt11_rxsyncallin_in                     : in   std_logic;
    gt11_rxsyncdone_out                     : out  std_logic;
    gt11_rxsyncin_in                        : in   std_logic;
    gt11_rxsyncmode_in                      : in   std_logic;
    gt11_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt11_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt11_rxlpmhfhold_in                     : in   std_logic;
    gt11_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt11_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt11_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt11_rxoutclk_out                       : out  std_logic;
    gt11_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt11_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt11_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt11_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt11_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt11_gttxreset_in                       : in   std_logic;
    gt11_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt11_txusrclk_in                        : in   std_logic;
    gt11_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt11_txdlyen_in                         : in   std_logic;
    gt11_txdlysreset_in                     : in   std_logic;
    gt11_txdlysresetdone_out                : out  std_logic;
    gt11_txphalign_in                       : in   std_logic;
    gt11_txphaligndone_out                  : out  std_logic;
    gt11_txphalignen_in                     : in   std_logic;
    gt11_txphdlyreset_in                    : in   std_logic;
    gt11_txphinit_in                        : in   std_logic;
    gt11_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt11_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt11_gthtxn_out                         : out  std_logic;
    gt11_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt11_txoutclk_out                       : out  std_logic;
    gt11_txoutclkfabric_out                 : out  std_logic;
    gt11_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt11_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt11_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT12  (X0Y16)
    --____________________________CHANNEL PORTS________________________________
    GT12_DRP_BUSY_OUT                        : out  std_logic; 
 GT12_RXPMARESETDONE_OUT  : out  std_logic;
 GT12_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt12_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt12_drpclk_in                          : in   std_logic;
    gt12_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt12_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt12_drpen_in                           : in   std_logic;
    gt12_drprdy_out                         : out  std_logic;
    gt12_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt12_eyescanreset_in                    : in   std_logic;
    gt12_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt12_eyescandataerror_out               : out  std_logic;
    gt12_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt12_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt12_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt12_rxusrclk_in                        : in   std_logic;
    gt12_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt12_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt12_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt12_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt12_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt12_rxdlyen_in                         : in   std_logic;
    gt12_rxdlysreset_in                     : in   std_logic;
    gt12_rxdlysresetdone_out                : out  std_logic;
    gt12_rxphalign_in                       : in   std_logic;
    gt12_rxphaligndone_out                  : out  std_logic;
    gt12_rxphalignen_in                     : in   std_logic;
    gt12_rxphdlyreset_in                    : in   std_logic;
    gt12_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt12_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt12_rxsyncallin_in                     : in   std_logic;
    gt12_rxsyncdone_out                     : out  std_logic;
    gt12_rxsyncin_in                        : in   std_logic;
    gt12_rxsyncmode_in                      : in   std_logic;
    gt12_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt12_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt12_rxlpmhfhold_in                     : in   std_logic;
    gt12_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt12_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt12_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt12_rxoutclk_out                       : out  std_logic;
    gt12_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt12_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt12_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt12_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt12_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt12_gttxreset_in                       : in   std_logic;
    gt12_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt12_txusrclk_in                        : in   std_logic;
    gt12_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt12_txdlyen_in                         : in   std_logic;
    gt12_txdlysreset_in                     : in   std_logic;
    gt12_txdlysresetdone_out                : out  std_logic;
    gt12_txphalign_in                       : in   std_logic;
    gt12_txphaligndone_out                  : out  std_logic;
    gt12_txphalignen_in                     : in   std_logic;
    gt12_txphdlyreset_in                    : in   std_logic;
    gt12_txphinit_in                        : in   std_logic;
    gt12_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt12_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt12_gthtxn_out                         : out  std_logic;
    gt12_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt12_txoutclk_out                       : out  std_logic;
    gt12_txoutclkfabric_out                 : out  std_logic;
    gt12_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt12_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt12_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT13  (X0Y17)
    --____________________________CHANNEL PORTS________________________________
    GT13_DRP_BUSY_OUT                        : out  std_logic; 
 GT13_RXPMARESETDONE_OUT  : out  std_logic;
 GT13_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt13_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt13_drpclk_in                          : in   std_logic;
    gt13_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt13_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt13_drpen_in                           : in   std_logic;
    gt13_drprdy_out                         : out  std_logic;
    gt13_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt13_eyescanreset_in                    : in   std_logic;
    gt13_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt13_eyescandataerror_out               : out  std_logic;
    gt13_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt13_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt13_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt13_rxusrclk_in                        : in   std_logic;
    gt13_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt13_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt13_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt13_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt13_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt13_rxdlyen_in                         : in   std_logic;
    gt13_rxdlysreset_in                     : in   std_logic;
    gt13_rxdlysresetdone_out                : out  std_logic;
    gt13_rxphalign_in                       : in   std_logic;
    gt13_rxphaligndone_out                  : out  std_logic;
    gt13_rxphalignen_in                     : in   std_logic;
    gt13_rxphdlyreset_in                    : in   std_logic;
    gt13_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt13_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt13_rxsyncallin_in                     : in   std_logic;
    gt13_rxsyncdone_out                     : out  std_logic;
    gt13_rxsyncin_in                        : in   std_logic;
    gt13_rxsyncmode_in                      : in   std_logic;
    gt13_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt13_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt13_rxlpmhfhold_in                     : in   std_logic;
    gt13_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt13_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt13_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt13_rxoutclk_out                       : out  std_logic;
    gt13_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt13_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt13_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt13_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt13_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt13_gttxreset_in                       : in   std_logic;
    gt13_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt13_txusrclk_in                        : in   std_logic;
    gt13_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt13_txdlyen_in                         : in   std_logic;
    gt13_txdlysreset_in                     : in   std_logic;
    gt13_txdlysresetdone_out                : out  std_logic;
    gt13_txphalign_in                       : in   std_logic;
    gt13_txphaligndone_out                  : out  std_logic;
    gt13_txphalignen_in                     : in   std_logic;
    gt13_txphdlyreset_in                    : in   std_logic;
    gt13_txphinit_in                        : in   std_logic;
    gt13_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt13_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt13_gthtxn_out                         : out  std_logic;
    gt13_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt13_txoutclk_out                       : out  std_logic;
    gt13_txoutclkfabric_out                 : out  std_logic;
    gt13_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt13_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt13_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT14  (X0Y18)
    --____________________________CHANNEL PORTS________________________________
    GT14_DRP_BUSY_OUT                        : out  std_logic; 
 GT14_RXPMARESETDONE_OUT  : out  std_logic;
 GT14_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt14_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt14_drpclk_in                          : in   std_logic;
    gt14_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt14_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt14_drpen_in                           : in   std_logic;
    gt14_drprdy_out                         : out  std_logic;
    gt14_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt14_eyescanreset_in                    : in   std_logic;
    gt14_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt14_eyescandataerror_out               : out  std_logic;
    gt14_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt14_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt14_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt14_rxusrclk_in                        : in   std_logic;
    gt14_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt14_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt14_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt14_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt14_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt14_rxdlyen_in                         : in   std_logic;
    gt14_rxdlysreset_in                     : in   std_logic;
    gt14_rxdlysresetdone_out                : out  std_logic;
    gt14_rxphalign_in                       : in   std_logic;
    gt14_rxphaligndone_out                  : out  std_logic;
    gt14_rxphalignen_in                     : in   std_logic;
    gt14_rxphdlyreset_in                    : in   std_logic;
    gt14_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt14_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt14_rxsyncallin_in                     : in   std_logic;
    gt14_rxsyncdone_out                     : out  std_logic;
    gt14_rxsyncin_in                        : in   std_logic;
    gt14_rxsyncmode_in                      : in   std_logic;
    gt14_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt14_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt14_rxlpmhfhold_in                     : in   std_logic;
    gt14_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt14_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt14_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt14_rxoutclk_out                       : out  std_logic;
    gt14_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt14_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt14_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt14_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt14_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt14_gttxreset_in                       : in   std_logic;
    gt14_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt14_txusrclk_in                        : in   std_logic;
    gt14_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt14_txdlyen_in                         : in   std_logic;
    gt14_txdlysreset_in                     : in   std_logic;
    gt14_txdlysresetdone_out                : out  std_logic;
    gt14_txphalign_in                       : in   std_logic;
    gt14_txphaligndone_out                  : out  std_logic;
    gt14_txphalignen_in                     : in   std_logic;
    gt14_txphdlyreset_in                    : in   std_logic;
    gt14_txphinit_in                        : in   std_logic;
    gt14_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt14_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt14_gthtxn_out                         : out  std_logic;
    gt14_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt14_txoutclk_out                       : out  std_logic;
    gt14_txoutclkfabric_out                 : out  std_logic;
    gt14_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt14_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt14_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT15  (X0Y19)
    --____________________________CHANNEL PORTS________________________________
    GT15_DRP_BUSY_OUT                        : out  std_logic; 
 GT15_RXPMARESETDONE_OUT  : out  std_logic;
 GT15_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt15_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt15_drpclk_in                          : in   std_logic;
    gt15_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt15_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt15_drpen_in                           : in   std_logic;
    gt15_drprdy_out                         : out  std_logic;
    gt15_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt15_eyescanreset_in                    : in   std_logic;
    gt15_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt15_eyescandataerror_out               : out  std_logic;
    gt15_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt15_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt15_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt15_rxusrclk_in                        : in   std_logic;
    gt15_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt15_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt15_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt15_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt15_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt15_rxdlyen_in                         : in   std_logic;
    gt15_rxdlysreset_in                     : in   std_logic;
    gt15_rxdlysresetdone_out                : out  std_logic;
    gt15_rxphalign_in                       : in   std_logic;
    gt15_rxphaligndone_out                  : out  std_logic;
    gt15_rxphalignen_in                     : in   std_logic;
    gt15_rxphdlyreset_in                    : in   std_logic;
    gt15_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt15_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt15_rxsyncallin_in                     : in   std_logic;
    gt15_rxsyncdone_out                     : out  std_logic;
    gt15_rxsyncin_in                        : in   std_logic;
    gt15_rxsyncmode_in                      : in   std_logic;
    gt15_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt15_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt15_rxlpmhfhold_in                     : in   std_logic;
    gt15_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt15_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt15_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt15_rxoutclk_out                       : out  std_logic;
    gt15_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt15_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt15_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt15_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt15_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt15_gttxreset_in                       : in   std_logic;
    gt15_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt15_txusrclk_in                        : in   std_logic;
    gt15_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt15_txdlyen_in                         : in   std_logic;
    gt15_txdlysreset_in                     : in   std_logic;
    gt15_txdlysresetdone_out                : out  std_logic;
    gt15_txphalign_in                       : in   std_logic;
    gt15_txphaligndone_out                  : out  std_logic;
    gt15_txphalignen_in                     : in   std_logic;
    gt15_txphdlyreset_in                    : in   std_logic;
    gt15_txphinit_in                        : in   std_logic;
    gt15_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt15_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt15_gthtxn_out                         : out  std_logic;
    gt15_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt15_txoutclk_out                       : out  std_logic;
    gt15_txoutclkfabric_out                 : out  std_logic;
    gt15_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt15_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt15_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT16  (X0Y20)
    --____________________________CHANNEL PORTS________________________________
    GT16_DRP_BUSY_OUT                        : out  std_logic; 
 GT16_RXPMARESETDONE_OUT  : out  std_logic;
 GT16_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt16_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt16_drpclk_in                          : in   std_logic;
    gt16_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt16_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt16_drpen_in                           : in   std_logic;
    gt16_drprdy_out                         : out  std_logic;
    gt16_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt16_eyescanreset_in                    : in   std_logic;
    gt16_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt16_eyescandataerror_out               : out  std_logic;
    gt16_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt16_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt16_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt16_rxusrclk_in                        : in   std_logic;
    gt16_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt16_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt16_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt16_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt16_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt16_rxdlyen_in                         : in   std_logic;
    gt16_rxdlysreset_in                     : in   std_logic;
    gt16_rxdlysresetdone_out                : out  std_logic;
    gt16_rxphalign_in                       : in   std_logic;
    gt16_rxphaligndone_out                  : out  std_logic;
    gt16_rxphalignen_in                     : in   std_logic;
    gt16_rxphdlyreset_in                    : in   std_logic;
    gt16_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt16_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt16_rxsyncallin_in                     : in   std_logic;
    gt16_rxsyncdone_out                     : out  std_logic;
    gt16_rxsyncin_in                        : in   std_logic;
    gt16_rxsyncmode_in                      : in   std_logic;
    gt16_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt16_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt16_rxlpmhfhold_in                     : in   std_logic;
    gt16_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt16_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt16_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt16_rxoutclk_out                       : out  std_logic;
    gt16_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt16_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt16_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt16_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt16_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt16_gttxreset_in                       : in   std_logic;
    gt16_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt16_txusrclk_in                        : in   std_logic;
    gt16_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt16_txdlyen_in                         : in   std_logic;
    gt16_txdlysreset_in                     : in   std_logic;
    gt16_txdlysresetdone_out                : out  std_logic;
    gt16_txphalign_in                       : in   std_logic;
    gt16_txphaligndone_out                  : out  std_logic;
    gt16_txphalignen_in                     : in   std_logic;
    gt16_txphdlyreset_in                    : in   std_logic;
    gt16_txphinit_in                        : in   std_logic;
    gt16_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt16_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt16_gthtxn_out                         : out  std_logic;
    gt16_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt16_txoutclk_out                       : out  std_logic;
    gt16_txoutclkfabric_out                 : out  std_logic;
    gt16_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt16_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt16_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT17  (X0Y21)
    --____________________________CHANNEL PORTS________________________________
    GT17_DRP_BUSY_OUT                        : out  std_logic; 
 GT17_RXPMARESETDONE_OUT  : out  std_logic;
 GT17_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt17_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt17_drpclk_in                          : in   std_logic;
    gt17_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt17_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt17_drpen_in                           : in   std_logic;
    gt17_drprdy_out                         : out  std_logic;
    gt17_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt17_eyescanreset_in                    : in   std_logic;
    gt17_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt17_eyescandataerror_out               : out  std_logic;
    gt17_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt17_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt17_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt17_rxusrclk_in                        : in   std_logic;
    gt17_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt17_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt17_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt17_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt17_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt17_rxdlyen_in                         : in   std_logic;
    gt17_rxdlysreset_in                     : in   std_logic;
    gt17_rxdlysresetdone_out                : out  std_logic;
    gt17_rxphalign_in                       : in   std_logic;
    gt17_rxphaligndone_out                  : out  std_logic;
    gt17_rxphalignen_in                     : in   std_logic;
    gt17_rxphdlyreset_in                    : in   std_logic;
    gt17_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt17_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt17_rxsyncallin_in                     : in   std_logic;
    gt17_rxsyncdone_out                     : out  std_logic;
    gt17_rxsyncin_in                        : in   std_logic;
    gt17_rxsyncmode_in                      : in   std_logic;
    gt17_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt17_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt17_rxlpmhfhold_in                     : in   std_logic;
    gt17_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt17_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt17_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt17_rxoutclk_out                       : out  std_logic;
    gt17_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt17_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt17_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt17_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt17_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt17_gttxreset_in                       : in   std_logic;
    gt17_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt17_txusrclk_in                        : in   std_logic;
    gt17_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt17_txdlyen_in                         : in   std_logic;
    gt17_txdlysreset_in                     : in   std_logic;
    gt17_txdlysresetdone_out                : out  std_logic;
    gt17_txphalign_in                       : in   std_logic;
    gt17_txphaligndone_out                  : out  std_logic;
    gt17_txphalignen_in                     : in   std_logic;
    gt17_txphdlyreset_in                    : in   std_logic;
    gt17_txphinit_in                        : in   std_logic;
    gt17_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt17_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt17_gthtxn_out                         : out  std_logic;
    gt17_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt17_txoutclk_out                       : out  std_logic;
    gt17_txoutclkfabric_out                 : out  std_logic;
    gt17_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt17_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt17_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT18  (X0Y22)
    --____________________________CHANNEL PORTS________________________________
    GT18_DRP_BUSY_OUT                        : out  std_logic; 
 GT18_RXPMARESETDONE_OUT  : out  std_logic;
 GT18_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt18_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt18_drpclk_in                          : in   std_logic;
    gt18_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt18_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt18_drpen_in                           : in   std_logic;
    gt18_drprdy_out                         : out  std_logic;
    gt18_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt18_eyescanreset_in                    : in   std_logic;
    gt18_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt18_eyescandataerror_out               : out  std_logic;
    gt18_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt18_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt18_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt18_rxusrclk_in                        : in   std_logic;
    gt18_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt18_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt18_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt18_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt18_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt18_rxdlyen_in                         : in   std_logic;
    gt18_rxdlysreset_in                     : in   std_logic;
    gt18_rxdlysresetdone_out                : out  std_logic;
    gt18_rxphalign_in                       : in   std_logic;
    gt18_rxphaligndone_out                  : out  std_logic;
    gt18_rxphalignen_in                     : in   std_logic;
    gt18_rxphdlyreset_in                    : in   std_logic;
    gt18_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt18_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt18_rxsyncallin_in                     : in   std_logic;
    gt18_rxsyncdone_out                     : out  std_logic;
    gt18_rxsyncin_in                        : in   std_logic;
    gt18_rxsyncmode_in                      : in   std_logic;
    gt18_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt18_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt18_rxlpmhfhold_in                     : in   std_logic;
    gt18_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt18_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt18_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt18_rxoutclk_out                       : out  std_logic;
    gt18_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt18_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt18_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt18_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt18_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt18_gttxreset_in                       : in   std_logic;
    gt18_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt18_txusrclk_in                        : in   std_logic;
    gt18_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt18_txdlyen_in                         : in   std_logic;
    gt18_txdlysreset_in                     : in   std_logic;
    gt18_txdlysresetdone_out                : out  std_logic;
    gt18_txphalign_in                       : in   std_logic;
    gt18_txphaligndone_out                  : out  std_logic;
    gt18_txphalignen_in                     : in   std_logic;
    gt18_txphdlyreset_in                    : in   std_logic;
    gt18_txphinit_in                        : in   std_logic;
    gt18_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt18_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt18_gthtxn_out                         : out  std_logic;
    gt18_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt18_txoutclk_out                       : out  std_logic;
    gt18_txoutclkfabric_out                 : out  std_logic;
    gt18_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt18_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt18_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT19  (X0Y23)
    --____________________________CHANNEL PORTS________________________________
    GT19_DRP_BUSY_OUT                        : out  std_logic; 
 GT19_RXPMARESETDONE_OUT  : out  std_logic;
 GT19_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt19_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt19_drpclk_in                          : in   std_logic;
    gt19_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt19_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt19_drpen_in                           : in   std_logic;
    gt19_drprdy_out                         : out  std_logic;
    gt19_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt19_eyescanreset_in                    : in   std_logic;
    gt19_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt19_eyescandataerror_out               : out  std_logic;
    gt19_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt19_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt19_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt19_rxusrclk_in                        : in   std_logic;
    gt19_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt19_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt19_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt19_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt19_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt19_rxdlyen_in                         : in   std_logic;
    gt19_rxdlysreset_in                     : in   std_logic;
    gt19_rxdlysresetdone_out                : out  std_logic;
    gt19_rxphalign_in                       : in   std_logic;
    gt19_rxphaligndone_out                  : out  std_logic;
    gt19_rxphalignen_in                     : in   std_logic;
    gt19_rxphdlyreset_in                    : in   std_logic;
    gt19_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt19_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt19_rxsyncallin_in                     : in   std_logic;
    gt19_rxsyncdone_out                     : out  std_logic;
    gt19_rxsyncin_in                        : in   std_logic;
    gt19_rxsyncmode_in                      : in   std_logic;
    gt19_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt19_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt19_rxlpmhfhold_in                     : in   std_logic;
    gt19_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt19_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt19_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt19_rxoutclk_out                       : out  std_logic;
    gt19_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt19_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt19_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt19_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt19_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt19_gttxreset_in                       : in   std_logic;
    gt19_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt19_txusrclk_in                        : in   std_logic;
    gt19_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt19_txdlyen_in                         : in   std_logic;
    gt19_txdlysreset_in                     : in   std_logic;
    gt19_txdlysresetdone_out                : out  std_logic;
    gt19_txphalign_in                       : in   std_logic;
    gt19_txphaligndone_out                  : out  std_logic;
    gt19_txphalignen_in                     : in   std_logic;
    gt19_txphdlyreset_in                    : in   std_logic;
    gt19_txphinit_in                        : in   std_logic;
    gt19_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt19_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt19_gthtxn_out                         : out  std_logic;
    gt19_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt19_txoutclk_out                       : out  std_logic;
    gt19_txoutclkfabric_out                 : out  std_logic;
    gt19_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt19_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt19_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT20  (X0Y24)
    --____________________________CHANNEL PORTS________________________________
    GT20_DRP_BUSY_OUT                        : out  std_logic; 
 GT20_RXPMARESETDONE_OUT  : out  std_logic;
 GT20_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt20_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt20_drpclk_in                          : in   std_logic;
    gt20_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt20_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt20_drpen_in                           : in   std_logic;
    gt20_drprdy_out                         : out  std_logic;
    gt20_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt20_eyescanreset_in                    : in   std_logic;
    gt20_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt20_eyescandataerror_out               : out  std_logic;
    gt20_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt20_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt20_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt20_rxusrclk_in                        : in   std_logic;
    gt20_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt20_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt20_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt20_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt20_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt20_rxdlyen_in                         : in   std_logic;
    gt20_rxdlysreset_in                     : in   std_logic;
    gt20_rxdlysresetdone_out                : out  std_logic;
    gt20_rxphalign_in                       : in   std_logic;
    gt20_rxphaligndone_out                  : out  std_logic;
    gt20_rxphalignen_in                     : in   std_logic;
    gt20_rxphdlyreset_in                    : in   std_logic;
    gt20_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt20_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt20_rxsyncallin_in                     : in   std_logic;
    gt20_rxsyncdone_out                     : out  std_logic;
    gt20_rxsyncin_in                        : in   std_logic;
    gt20_rxsyncmode_in                      : in   std_logic;
    gt20_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt20_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt20_rxlpmhfhold_in                     : in   std_logic;
    gt20_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt20_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt20_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt20_rxoutclk_out                       : out  std_logic;
    gt20_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt20_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt20_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt20_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt20_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt20_gttxreset_in                       : in   std_logic;
    gt20_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt20_txusrclk_in                        : in   std_logic;
    gt20_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt20_txdlyen_in                         : in   std_logic;
    gt20_txdlysreset_in                     : in   std_logic;
    gt20_txdlysresetdone_out                : out  std_logic;
    gt20_txphalign_in                       : in   std_logic;
    gt20_txphaligndone_out                  : out  std_logic;
    gt20_txphalignen_in                     : in   std_logic;
    gt20_txphdlyreset_in                    : in   std_logic;
    gt20_txphinit_in                        : in   std_logic;
    gt20_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt20_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt20_gthtxn_out                         : out  std_logic;
    gt20_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt20_txoutclk_out                       : out  std_logic;
    gt20_txoutclkfabric_out                 : out  std_logic;
    gt20_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt20_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt20_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT21  (X0Y25)
    --____________________________CHANNEL PORTS________________________________
    GT21_DRP_BUSY_OUT                        : out  std_logic; 
 GT21_RXPMARESETDONE_OUT  : out  std_logic;
 GT21_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt21_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt21_drpclk_in                          : in   std_logic;
    gt21_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt21_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt21_drpen_in                           : in   std_logic;
    gt21_drprdy_out                         : out  std_logic;
    gt21_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt21_eyescanreset_in                    : in   std_logic;
    gt21_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt21_eyescandataerror_out               : out  std_logic;
    gt21_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt21_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt21_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt21_rxusrclk_in                        : in   std_logic;
    gt21_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt21_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt21_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt21_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt21_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt21_rxdlyen_in                         : in   std_logic;
    gt21_rxdlysreset_in                     : in   std_logic;
    gt21_rxdlysresetdone_out                : out  std_logic;
    gt21_rxphalign_in                       : in   std_logic;
    gt21_rxphaligndone_out                  : out  std_logic;
    gt21_rxphalignen_in                     : in   std_logic;
    gt21_rxphdlyreset_in                    : in   std_logic;
    gt21_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt21_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt21_rxsyncallin_in                     : in   std_logic;
    gt21_rxsyncdone_out                     : out  std_logic;
    gt21_rxsyncin_in                        : in   std_logic;
    gt21_rxsyncmode_in                      : in   std_logic;
    gt21_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt21_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt21_rxlpmhfhold_in                     : in   std_logic;
    gt21_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt21_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt21_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt21_rxoutclk_out                       : out  std_logic;
    gt21_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt21_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt21_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt21_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt21_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt21_gttxreset_in                       : in   std_logic;
    gt21_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt21_txusrclk_in                        : in   std_logic;
    gt21_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt21_txdlyen_in                         : in   std_logic;
    gt21_txdlysreset_in                     : in   std_logic;
    gt21_txdlysresetdone_out                : out  std_logic;
    gt21_txphalign_in                       : in   std_logic;
    gt21_txphaligndone_out                  : out  std_logic;
    gt21_txphalignen_in                     : in   std_logic;
    gt21_txphdlyreset_in                    : in   std_logic;
    gt21_txphinit_in                        : in   std_logic;
    gt21_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt21_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt21_gthtxn_out                         : out  std_logic;
    gt21_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt21_txoutclk_out                       : out  std_logic;
    gt21_txoutclkfabric_out                 : out  std_logic;
    gt21_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt21_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt21_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT22  (X0Y26)
    --____________________________CHANNEL PORTS________________________________
    GT22_DRP_BUSY_OUT                        : out  std_logic; 
 GT22_RXPMARESETDONE_OUT  : out  std_logic;
 GT22_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt22_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt22_drpclk_in                          : in   std_logic;
    gt22_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt22_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt22_drpen_in                           : in   std_logic;
    gt22_drprdy_out                         : out  std_logic;
    gt22_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt22_eyescanreset_in                    : in   std_logic;
    gt22_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt22_eyescandataerror_out               : out  std_logic;
    gt22_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt22_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt22_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt22_rxusrclk_in                        : in   std_logic;
    gt22_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt22_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt22_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt22_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt22_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt22_rxdlyen_in                         : in   std_logic;
    gt22_rxdlysreset_in                     : in   std_logic;
    gt22_rxdlysresetdone_out                : out  std_logic;
    gt22_rxphalign_in                       : in   std_logic;
    gt22_rxphaligndone_out                  : out  std_logic;
    gt22_rxphalignen_in                     : in   std_logic;
    gt22_rxphdlyreset_in                    : in   std_logic;
    gt22_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt22_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt22_rxsyncallin_in                     : in   std_logic;
    gt22_rxsyncdone_out                     : out  std_logic;
    gt22_rxsyncin_in                        : in   std_logic;
    gt22_rxsyncmode_in                      : in   std_logic;
    gt22_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt22_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt22_rxlpmhfhold_in                     : in   std_logic;
    gt22_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt22_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt22_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt22_rxoutclk_out                       : out  std_logic;
    gt22_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt22_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt22_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt22_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt22_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt22_gttxreset_in                       : in   std_logic;
    gt22_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt22_txusrclk_in                        : in   std_logic;
    gt22_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt22_txdlyen_in                         : in   std_logic;
    gt22_txdlysreset_in                     : in   std_logic;
    gt22_txdlysresetdone_out                : out  std_logic;
    gt22_txphalign_in                       : in   std_logic;
    gt22_txphaligndone_out                  : out  std_logic;
    gt22_txphalignen_in                     : in   std_logic;
    gt22_txphdlyreset_in                    : in   std_logic;
    gt22_txphinit_in                        : in   std_logic;
    gt22_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt22_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt22_gthtxn_out                         : out  std_logic;
    gt22_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt22_txoutclk_out                       : out  std_logic;
    gt22_txoutclkfabric_out                 : out  std_logic;
    gt22_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt22_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt22_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT23  (X0Y27)
    --____________________________CHANNEL PORTS________________________________
    GT23_DRP_BUSY_OUT                        : out  std_logic; 
 GT23_RXPMARESETDONE_OUT  : out  std_logic;
 GT23_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt23_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt23_drpclk_in                          : in   std_logic;
    gt23_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt23_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt23_drpen_in                           : in   std_logic;
    gt23_drprdy_out                         : out  std_logic;
    gt23_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt23_eyescanreset_in                    : in   std_logic;
    gt23_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt23_eyescandataerror_out               : out  std_logic;
    gt23_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt23_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt23_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt23_rxusrclk_in                        : in   std_logic;
    gt23_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt23_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt23_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt23_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt23_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt23_rxdlyen_in                         : in   std_logic;
    gt23_rxdlysreset_in                     : in   std_logic;
    gt23_rxdlysresetdone_out                : out  std_logic;
    gt23_rxphalign_in                       : in   std_logic;
    gt23_rxphaligndone_out                  : out  std_logic;
    gt23_rxphalignen_in                     : in   std_logic;
    gt23_rxphdlyreset_in                    : in   std_logic;
    gt23_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt23_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt23_rxsyncallin_in                     : in   std_logic;
    gt23_rxsyncdone_out                     : out  std_logic;
    gt23_rxsyncin_in                        : in   std_logic;
    gt23_rxsyncmode_in                      : in   std_logic;
    gt23_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt23_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt23_rxlpmhfhold_in                     : in   std_logic;
    gt23_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt23_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt23_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt23_rxoutclk_out                       : out  std_logic;
    gt23_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt23_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt23_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt23_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt23_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt23_gttxreset_in                       : in   std_logic;
    gt23_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt23_txusrclk_in                        : in   std_logic;
    gt23_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt23_txdlyen_in                         : in   std_logic;
    gt23_txdlysreset_in                     : in   std_logic;
    gt23_txdlysresetdone_out                : out  std_logic;
    gt23_txphalign_in                       : in   std_logic;
    gt23_txphaligndone_out                  : out  std_logic;
    gt23_txphalignen_in                     : in   std_logic;
    gt23_txphdlyreset_in                    : in   std_logic;
    gt23_txphinit_in                        : in   std_logic;
    gt23_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt23_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt23_gthtxn_out                         : out  std_logic;
    gt23_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt23_txoutclk_out                       : out  std_logic;
    gt23_txoutclkfabric_out                 : out  std_logic;
    gt23_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt23_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt23_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT24  (X0Y28)
    --____________________________CHANNEL PORTS________________________________
    GT24_DRP_BUSY_OUT                        : out  std_logic; 
 GT24_RXPMARESETDONE_OUT  : out  std_logic;
 GT24_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt24_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt24_drpclk_in                          : in   std_logic;
    gt24_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt24_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt24_drpen_in                           : in   std_logic;
    gt24_drprdy_out                         : out  std_logic;
    gt24_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt24_eyescanreset_in                    : in   std_logic;
    gt24_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt24_eyescandataerror_out               : out  std_logic;
    gt24_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt24_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt24_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt24_rxusrclk_in                        : in   std_logic;
    gt24_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt24_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt24_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt24_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt24_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt24_rxdlyen_in                         : in   std_logic;
    gt24_rxdlysreset_in                     : in   std_logic;
    gt24_rxdlysresetdone_out                : out  std_logic;
    gt24_rxphalign_in                       : in   std_logic;
    gt24_rxphaligndone_out                  : out  std_logic;
    gt24_rxphalignen_in                     : in   std_logic;
    gt24_rxphdlyreset_in                    : in   std_logic;
    gt24_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt24_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt24_rxsyncallin_in                     : in   std_logic;
    gt24_rxsyncdone_out                     : out  std_logic;
    gt24_rxsyncin_in                        : in   std_logic;
    gt24_rxsyncmode_in                      : in   std_logic;
    gt24_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt24_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt24_rxlpmhfhold_in                     : in   std_logic;
    gt24_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt24_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt24_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt24_rxoutclk_out                       : out  std_logic;
    gt24_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt24_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt24_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt24_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt24_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt24_gttxreset_in                       : in   std_logic;
    gt24_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt24_txusrclk_in                        : in   std_logic;
    gt24_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt24_txdlyen_in                         : in   std_logic;
    gt24_txdlysreset_in                     : in   std_logic;
    gt24_txdlysresetdone_out                : out  std_logic;
    gt24_txphalign_in                       : in   std_logic;
    gt24_txphaligndone_out                  : out  std_logic;
    gt24_txphalignen_in                     : in   std_logic;
    gt24_txphdlyreset_in                    : in   std_logic;
    gt24_txphinit_in                        : in   std_logic;
    gt24_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt24_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt24_gthtxn_out                         : out  std_logic;
    gt24_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt24_txoutclk_out                       : out  std_logic;
    gt24_txoutclkfabric_out                 : out  std_logic;
    gt24_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt24_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt24_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT25  (X0Y29)
    --____________________________CHANNEL PORTS________________________________
    GT25_DRP_BUSY_OUT                        : out  std_logic; 
 GT25_RXPMARESETDONE_OUT  : out  std_logic;
 GT25_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt25_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt25_drpclk_in                          : in   std_logic;
    gt25_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt25_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt25_drpen_in                           : in   std_logic;
    gt25_drprdy_out                         : out  std_logic;
    gt25_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt25_eyescanreset_in                    : in   std_logic;
    gt25_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt25_eyescandataerror_out               : out  std_logic;
    gt25_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt25_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt25_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt25_rxusrclk_in                        : in   std_logic;
    gt25_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt25_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt25_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt25_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt25_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt25_rxdlyen_in                         : in   std_logic;
    gt25_rxdlysreset_in                     : in   std_logic;
    gt25_rxdlysresetdone_out                : out  std_logic;
    gt25_rxphalign_in                       : in   std_logic;
    gt25_rxphaligndone_out                  : out  std_logic;
    gt25_rxphalignen_in                     : in   std_logic;
    gt25_rxphdlyreset_in                    : in   std_logic;
    gt25_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt25_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt25_rxsyncallin_in                     : in   std_logic;
    gt25_rxsyncdone_out                     : out  std_logic;
    gt25_rxsyncin_in                        : in   std_logic;
    gt25_rxsyncmode_in                      : in   std_logic;
    gt25_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt25_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt25_rxlpmhfhold_in                     : in   std_logic;
    gt25_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt25_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt25_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt25_rxoutclk_out                       : out  std_logic;
    gt25_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt25_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt25_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt25_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt25_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt25_gttxreset_in                       : in   std_logic;
    gt25_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt25_txusrclk_in                        : in   std_logic;
    gt25_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt25_txdlyen_in                         : in   std_logic;
    gt25_txdlysreset_in                     : in   std_logic;
    gt25_txdlysresetdone_out                : out  std_logic;
    gt25_txphalign_in                       : in   std_logic;
    gt25_txphaligndone_out                  : out  std_logic;
    gt25_txphalignen_in                     : in   std_logic;
    gt25_txphdlyreset_in                    : in   std_logic;
    gt25_txphinit_in                        : in   std_logic;
    gt25_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt25_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt25_gthtxn_out                         : out  std_logic;
    gt25_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt25_txoutclk_out                       : out  std_logic;
    gt25_txoutclkfabric_out                 : out  std_logic;
    gt25_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt25_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt25_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT26  (X0Y30)
    --____________________________CHANNEL PORTS________________________________
    GT26_DRP_BUSY_OUT                        : out  std_logic; 
 GT26_RXPMARESETDONE_OUT  : out  std_logic;
 GT26_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt26_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt26_drpclk_in                          : in   std_logic;
    gt26_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt26_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt26_drpen_in                           : in   std_logic;
    gt26_drprdy_out                         : out  std_logic;
    gt26_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt26_eyescanreset_in                    : in   std_logic;
    gt26_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt26_eyescandataerror_out               : out  std_logic;
    gt26_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt26_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt26_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt26_rxusrclk_in                        : in   std_logic;
    gt26_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt26_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt26_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt26_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt26_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt26_rxdlyen_in                         : in   std_logic;
    gt26_rxdlysreset_in                     : in   std_logic;
    gt26_rxdlysresetdone_out                : out  std_logic;
    gt26_rxphalign_in                       : in   std_logic;
    gt26_rxphaligndone_out                  : out  std_logic;
    gt26_rxphalignen_in                     : in   std_logic;
    gt26_rxphdlyreset_in                    : in   std_logic;
    gt26_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt26_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt26_rxsyncallin_in                     : in   std_logic;
    gt26_rxsyncdone_out                     : out  std_logic;
    gt26_rxsyncin_in                        : in   std_logic;
    gt26_rxsyncmode_in                      : in   std_logic;
    gt26_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt26_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt26_rxlpmhfhold_in                     : in   std_logic;
    gt26_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt26_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt26_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt26_rxoutclk_out                       : out  std_logic;
    gt26_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt26_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt26_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt26_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt26_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt26_gttxreset_in                       : in   std_logic;
    gt26_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt26_txusrclk_in                        : in   std_logic;
    gt26_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt26_txdlyen_in                         : in   std_logic;
    gt26_txdlysreset_in                     : in   std_logic;
    gt26_txdlysresetdone_out                : out  std_logic;
    gt26_txphalign_in                       : in   std_logic;
    gt26_txphaligndone_out                  : out  std_logic;
    gt26_txphalignen_in                     : in   std_logic;
    gt26_txphdlyreset_in                    : in   std_logic;
    gt26_txphinit_in                        : in   std_logic;
    gt26_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt26_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt26_gthtxn_out                         : out  std_logic;
    gt26_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt26_txoutclk_out                       : out  std_logic;
    gt26_txoutclkfabric_out                 : out  std_logic;
    gt26_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt26_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt26_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT27  (X0Y31)
    --____________________________CHANNEL PORTS________________________________
    GT27_DRP_BUSY_OUT                        : out  std_logic; 
 GT27_RXPMARESETDONE_OUT  : out  std_logic;
 GT27_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt27_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt27_drpclk_in                          : in   std_logic;
    gt27_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt27_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt27_drpen_in                           : in   std_logic;
    gt27_drprdy_out                         : out  std_logic;
    gt27_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt27_eyescanreset_in                    : in   std_logic;
    gt27_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt27_eyescandataerror_out               : out  std_logic;
    gt27_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt27_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt27_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt27_rxusrclk_in                        : in   std_logic;
    gt27_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt27_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt27_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt27_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt27_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt27_rxdlyen_in                         : in   std_logic;
    gt27_rxdlysreset_in                     : in   std_logic;
    gt27_rxdlysresetdone_out                : out  std_logic;
    gt27_rxphalign_in                       : in   std_logic;
    gt27_rxphaligndone_out                  : out  std_logic;
    gt27_rxphalignen_in                     : in   std_logic;
    gt27_rxphdlyreset_in                    : in   std_logic;
    gt27_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt27_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt27_rxsyncallin_in                     : in   std_logic;
    gt27_rxsyncdone_out                     : out  std_logic;
    gt27_rxsyncin_in                        : in   std_logic;
    gt27_rxsyncmode_in                      : in   std_logic;
    gt27_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt27_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt27_rxlpmhfhold_in                     : in   std_logic;
    gt27_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt27_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt27_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt27_rxoutclk_out                       : out  std_logic;
    gt27_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt27_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt27_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt27_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt27_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt27_gttxreset_in                       : in   std_logic;
    gt27_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt27_txusrclk_in                        : in   std_logic;
    gt27_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt27_txdlyen_in                         : in   std_logic;
    gt27_txdlysreset_in                     : in   std_logic;
    gt27_txdlysresetdone_out                : out  std_logic;
    gt27_txphalign_in                       : in   std_logic;
    gt27_txphaligndone_out                  : out  std_logic;
    gt27_txphalignen_in                     : in   std_logic;
    gt27_txphdlyreset_in                    : in   std_logic;
    gt27_txphinit_in                        : in   std_logic;
    gt27_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt27_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt27_gthtxn_out                         : out  std_logic;
    gt27_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt27_txoutclk_out                       : out  std_logic;
    gt27_txoutclkfabric_out                 : out  std_logic;
    gt27_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt27_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt27_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT28  (X0Y32)
    --____________________________CHANNEL PORTS________________________________
    GT28_DRP_BUSY_OUT                        : out  std_logic; 
 GT28_RXPMARESETDONE_OUT  : out  std_logic;
 GT28_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt28_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt28_drpclk_in                          : in   std_logic;
    gt28_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt28_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt28_drpen_in                           : in   std_logic;
    gt28_drprdy_out                         : out  std_logic;
    gt28_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt28_eyescanreset_in                    : in   std_logic;
    gt28_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt28_eyescandataerror_out               : out  std_logic;
    gt28_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt28_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt28_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt28_rxusrclk_in                        : in   std_logic;
    gt28_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt28_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt28_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt28_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt28_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt28_rxdlyen_in                         : in   std_logic;
    gt28_rxdlysreset_in                     : in   std_logic;
    gt28_rxdlysresetdone_out                : out  std_logic;
    gt28_rxphalign_in                       : in   std_logic;
    gt28_rxphaligndone_out                  : out  std_logic;
    gt28_rxphalignen_in                     : in   std_logic;
    gt28_rxphdlyreset_in                    : in   std_logic;
    gt28_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt28_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt28_rxsyncallin_in                     : in   std_logic;
    gt28_rxsyncdone_out                     : out  std_logic;
    gt28_rxsyncin_in                        : in   std_logic;
    gt28_rxsyncmode_in                      : in   std_logic;
    gt28_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt28_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt28_rxlpmhfhold_in                     : in   std_logic;
    gt28_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt28_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt28_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt28_rxoutclk_out                       : out  std_logic;
    gt28_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt28_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt28_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt28_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt28_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt28_gttxreset_in                       : in   std_logic;
    gt28_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt28_txusrclk_in                        : in   std_logic;
    gt28_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt28_txdlyen_in                         : in   std_logic;
    gt28_txdlysreset_in                     : in   std_logic;
    gt28_txdlysresetdone_out                : out  std_logic;
    gt28_txphalign_in                       : in   std_logic;
    gt28_txphaligndone_out                  : out  std_logic;
    gt28_txphalignen_in                     : in   std_logic;
    gt28_txphdlyreset_in                    : in   std_logic;
    gt28_txphinit_in                        : in   std_logic;
    gt28_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt28_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt28_gthtxn_out                         : out  std_logic;
    gt28_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt28_txoutclk_out                       : out  std_logic;
    gt28_txoutclkfabric_out                 : out  std_logic;
    gt28_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt28_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt28_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT29  (X0Y33)
    --____________________________CHANNEL PORTS________________________________
    GT29_DRP_BUSY_OUT                        : out  std_logic; 
 GT29_RXPMARESETDONE_OUT  : out  std_logic;
 GT29_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt29_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt29_drpclk_in                          : in   std_logic;
    gt29_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt29_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt29_drpen_in                           : in   std_logic;
    gt29_drprdy_out                         : out  std_logic;
    gt29_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt29_eyescanreset_in                    : in   std_logic;
    gt29_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt29_eyescandataerror_out               : out  std_logic;
    gt29_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt29_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt29_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt29_rxusrclk_in                        : in   std_logic;
    gt29_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt29_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt29_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt29_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt29_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt29_rxdlyen_in                         : in   std_logic;
    gt29_rxdlysreset_in                     : in   std_logic;
    gt29_rxdlysresetdone_out                : out  std_logic;
    gt29_rxphalign_in                       : in   std_logic;
    gt29_rxphaligndone_out                  : out  std_logic;
    gt29_rxphalignen_in                     : in   std_logic;
    gt29_rxphdlyreset_in                    : in   std_logic;
    gt29_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt29_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt29_rxsyncallin_in                     : in   std_logic;
    gt29_rxsyncdone_out                     : out  std_logic;
    gt29_rxsyncin_in                        : in   std_logic;
    gt29_rxsyncmode_in                      : in   std_logic;
    gt29_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt29_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt29_rxlpmhfhold_in                     : in   std_logic;
    gt29_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt29_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt29_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt29_rxoutclk_out                       : out  std_logic;
    gt29_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt29_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt29_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt29_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt29_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt29_gttxreset_in                       : in   std_logic;
    gt29_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt29_txusrclk_in                        : in   std_logic;
    gt29_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt29_txdlyen_in                         : in   std_logic;
    gt29_txdlysreset_in                     : in   std_logic;
    gt29_txdlysresetdone_out                : out  std_logic;
    gt29_txphalign_in                       : in   std_logic;
    gt29_txphaligndone_out                  : out  std_logic;
    gt29_txphalignen_in                     : in   std_logic;
    gt29_txphdlyreset_in                    : in   std_logic;
    gt29_txphinit_in                        : in   std_logic;
    gt29_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt29_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt29_gthtxn_out                         : out  std_logic;
    gt29_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt29_txoutclk_out                       : out  std_logic;
    gt29_txoutclkfabric_out                 : out  std_logic;
    gt29_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt29_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt29_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT30  (X0Y34)
    --____________________________CHANNEL PORTS________________________________
    GT30_DRP_BUSY_OUT                        : out  std_logic; 
 GT30_RXPMARESETDONE_OUT  : out  std_logic;
 GT30_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt30_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt30_drpclk_in                          : in   std_logic;
    gt30_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt30_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt30_drpen_in                           : in   std_logic;
    gt30_drprdy_out                         : out  std_logic;
    gt30_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt30_eyescanreset_in                    : in   std_logic;
    gt30_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt30_eyescandataerror_out               : out  std_logic;
    gt30_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt30_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt30_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt30_rxusrclk_in                        : in   std_logic;
    gt30_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt30_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt30_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt30_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt30_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt30_rxdlyen_in                         : in   std_logic;
    gt30_rxdlysreset_in                     : in   std_logic;
    gt30_rxdlysresetdone_out                : out  std_logic;
    gt30_rxphalign_in                       : in   std_logic;
    gt30_rxphaligndone_out                  : out  std_logic;
    gt30_rxphalignen_in                     : in   std_logic;
    gt30_rxphdlyreset_in                    : in   std_logic;
    gt30_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt30_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt30_rxsyncallin_in                     : in   std_logic;
    gt30_rxsyncdone_out                     : out  std_logic;
    gt30_rxsyncin_in                        : in   std_logic;
    gt30_rxsyncmode_in                      : in   std_logic;
    gt30_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt30_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt30_rxlpmhfhold_in                     : in   std_logic;
    gt30_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt30_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt30_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt30_rxoutclk_out                       : out  std_logic;
    gt30_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt30_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt30_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt30_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt30_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt30_gttxreset_in                       : in   std_logic;
    gt30_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt30_txusrclk_in                        : in   std_logic;
    gt30_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt30_txdlyen_in                         : in   std_logic;
    gt30_txdlysreset_in                     : in   std_logic;
    gt30_txdlysresetdone_out                : out  std_logic;
    gt30_txphalign_in                       : in   std_logic;
    gt30_txphaligndone_out                  : out  std_logic;
    gt30_txphalignen_in                     : in   std_logic;
    gt30_txphdlyreset_in                    : in   std_logic;
    gt30_txphinit_in                        : in   std_logic;
    gt30_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt30_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt30_gthtxn_out                         : out  std_logic;
    gt30_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt30_txoutclk_out                       : out  std_logic;
    gt30_txoutclkfabric_out                 : out  std_logic;
    gt30_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt30_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt30_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT31  (X0Y35)
    --____________________________CHANNEL PORTS________________________________
    GT31_DRP_BUSY_OUT                        : out  std_logic; 
 GT31_RXPMARESETDONE_OUT  : out  std_logic;
 GT31_TXPMARESETDONE_OUT  : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt31_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt31_drpclk_in                          : in   std_logic;
    gt31_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt31_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt31_drpen_in                           : in   std_logic;
    gt31_drprdy_out                         : out  std_logic;
    gt31_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt31_eyescanreset_in                    : in   std_logic;
    gt31_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt31_eyescandataerror_out               : out  std_logic;
    gt31_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt31_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt31_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt31_rxusrclk_in                        : in   std_logic;
    gt31_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt31_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt31_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt31_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt31_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt31_rxdlyen_in                         : in   std_logic;
    gt31_rxdlysreset_in                     : in   std_logic;
    gt31_rxdlysresetdone_out                : out  std_logic;
    gt31_rxphalign_in                       : in   std_logic;
    gt31_rxphaligndone_out                  : out  std_logic;
    gt31_rxphalignen_in                     : in   std_logic;
    gt31_rxphdlyreset_in                    : in   std_logic;
    gt31_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt31_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    gt31_rxsyncallin_in                     : in   std_logic;
    gt31_rxsyncdone_out                     : out  std_logic;
    gt31_rxsyncin_in                        : in   std_logic;
    gt31_rxsyncmode_in                      : in   std_logic;
    gt31_rxsyncout_out                      : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt31_rxbyteisaligned_out                : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt31_rxlpmhfhold_in                     : in   std_logic;
    gt31_rxlpmlfhold_in                     : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt31_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt31_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt31_rxoutclk_out                       : out  std_logic;
    gt31_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt31_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt31_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt31_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt31_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt31_gttxreset_in                       : in   std_logic;
    gt31_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt31_txusrclk_in                        : in   std_logic;
    gt31_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt31_txdlyen_in                         : in   std_logic;
    gt31_txdlysreset_in                     : in   std_logic;
    gt31_txdlysresetdone_out                : out  std_logic;
    gt31_txphalign_in                       : in   std_logic;
    gt31_txphaligndone_out                  : out  std_logic;
    gt31_txphalignen_in                     : in   std_logic;
    gt31_txphdlyreset_in                    : in   std_logic;
    gt31_txphinit_in                        : in   std_logic;
    gt31_txphinitdone_out                   : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt31_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt31_gthtxn_out                         : out  std_logic;
    gt31_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt31_txoutclk_out                       : out  std_logic;
    gt31_txoutclkfabric_out                 : out  std_logic;
    gt31_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt31_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt31_txcharisk_in                       : in   std_logic_vector(7 downto 0);


    --____________________________COMMON PORTS________________________________
     GT0_QPLLOUTCLK_IN : in std_logic;
     GT0_QPLLRESET_IN  : in std_logic;
     GT0_QPLLOUTREFCLK_IN  : in std_logic;
    --____________________________COMMON PORTS________________________________
     GT1_QPLLOUTCLK_IN : in std_logic;
     GT1_QPLLRESET_IN  : in std_logic;
     GT1_QPLLOUTREFCLK_IN  : in std_logic;
    --____________________________COMMON PORTS________________________________
     GT2_QPLLOUTCLK_IN : in std_logic;
     GT2_QPLLRESET_IN  : in std_logic;
     GT2_QPLLOUTREFCLK_IN  : in std_logic;
    --____________________________COMMON PORTS________________________________
     GT3_QPLLOUTCLK_IN : in std_logic;
     GT3_QPLLRESET_IN  : in std_logic;
     GT3_QPLLOUTREFCLK_IN  : in std_logic;
    --____________________________COMMON PORTS________________________________
     GT4_QPLLOUTCLK_IN : in std_logic;
     GT4_QPLLRESET_IN  : in std_logic;
     GT4_QPLLOUTREFCLK_IN  : in std_logic;
    --____________________________COMMON PORTS________________________________
     GT5_QPLLOUTCLK_IN : in std_logic;
     GT5_QPLLRESET_IN  : in std_logic;
     GT5_QPLLOUTREFCLK_IN  : in std_logic;
    --____________________________COMMON PORTS________________________________
     GT6_QPLLOUTCLK_IN : in std_logic;
     GT6_QPLLRESET_IN  : in std_logic;
     GT6_QPLLOUTREFCLK_IN  : in std_logic;
    --____________________________COMMON PORTS________________________________
     GT7_QPLLOUTCLK_IN : in std_logic;
     GT7_QPLLRESET_IN  : in std_logic;
     GT7_QPLLOUTREFCLK_IN  : in std_logic

);


end gtwizard_0_multi_gt;
    
architecture RTL of gtwizard_0_multi_gt is
    attribute DowngradeIPIdentifiedWarnings: string;
    attribute DowngradeIPIdentifiedWarnings of RTL : architecture is "yes";

    attribute CORE_GENERATION_INFO : string;
    attribute CORE_GENERATION_INFO of RTL : architecture is "gtwizard_0_multi_gt,gtwizard_v3_6_9,{protocol_file=Start_from_scratch}";


--***********************************Parameter Declarations********************

    constant DLY : time := 1 ns;

--***************************** Signal Declarations *****************************

    -- ground and tied_to_vcc_i signals
signal  tied_to_ground_i                :   std_logic;
signal  tied_to_ground_vec_i            :   std_logic_vector(63 downto 0);
signal  tied_to_vcc_i                   :   std_logic;
signal   gt0_qplloutclk_i         :   std_logic;
signal   gt0_qplloutrefclk_i      :   std_logic;
signal   gt1_qplloutclk_i         :   std_logic;
signal   gt1_qplloutrefclk_i      :   std_logic;
signal   gt2_qplloutclk_i         :   std_logic;
signal   gt2_qplloutrefclk_i      :   std_logic;
signal   gt3_qplloutclk_i         :   std_logic;
signal   gt3_qplloutrefclk_i      :   std_logic;
signal   gt4_qplloutclk_i         :   std_logic;
signal   gt4_qplloutrefclk_i      :   std_logic;
signal   gt5_qplloutclk_i         :   std_logic;
signal   gt5_qplloutrefclk_i      :   std_logic;
signal   gt6_qplloutclk_i         :   std_logic;
signal   gt6_qplloutrefclk_i      :   std_logic;
signal   gt7_qplloutclk_i         :   std_logic;
signal   gt7_qplloutrefclk_i      :   std_logic;

signal  gt0_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt0_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt1_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt1_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt2_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt2_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt3_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt3_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt4_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt4_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt5_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt5_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt6_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt6_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt7_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt7_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt8_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt8_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt9_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt9_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt10_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt10_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt11_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt11_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt12_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt12_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt13_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt13_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt14_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt14_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt15_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt15_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt16_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt16_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt17_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt17_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt18_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt18_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt19_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt19_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt20_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt20_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt21_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt21_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt22_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt22_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt23_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt23_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt24_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt24_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt25_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt25_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt26_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt26_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt27_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt27_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt28_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt28_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt29_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt29_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt30_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt30_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt31_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt31_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
signal   gt0_qpllclk_i            :   std_logic;
signal   gt0_qpllrefclk_i         :   std_logic;
    signal    gt0_rst_i                       : std_logic;
signal   gt1_qpllclk_i            :   std_logic;
signal   gt1_qpllrefclk_i         :   std_logic;
    signal    gt1_rst_i                       : std_logic;
signal   gt2_qpllclk_i            :   std_logic;
signal   gt2_qpllrefclk_i         :   std_logic;
    signal    gt2_rst_i                       : std_logic;
signal   gt3_qpllclk_i            :   std_logic;
signal   gt3_qpllrefclk_i         :   std_logic;
    signal    gt3_rst_i                       : std_logic;
signal   gt4_qpllclk_i            :   std_logic;
signal   gt4_qpllrefclk_i         :   std_logic;
    signal    gt4_rst_i                       : std_logic;
signal   gt5_qpllclk_i            :   std_logic;
signal   gt5_qpllrefclk_i         :   std_logic;
    signal    gt5_rst_i                       : std_logic;
signal   gt6_qpllclk_i            :   std_logic;
signal   gt6_qpllrefclk_i         :   std_logic;
    signal    gt6_rst_i                       : std_logic;
signal   gt7_qpllclk_i            :   std_logic;
signal   gt7_qpllrefclk_i         :   std_logic;
    signal    gt7_rst_i                       : std_logic;
signal   gt8_qpllclk_i            :   std_logic;
signal   gt8_qpllrefclk_i         :   std_logic;
    signal    gt8_rst_i                       : std_logic;
signal   gt9_qpllclk_i            :   std_logic;
signal   gt9_qpllrefclk_i         :   std_logic;
    signal    gt9_rst_i                       : std_logic;
signal   gt10_qpllclk_i            :   std_logic;
signal   gt10_qpllrefclk_i         :   std_logic;
    signal    gt10_rst_i                      : std_logic;
signal   gt11_qpllclk_i            :   std_logic;
signal   gt11_qpllrefclk_i         :   std_logic;
    signal    gt11_rst_i                      : std_logic;
signal   gt12_qpllclk_i            :   std_logic;
signal   gt12_qpllrefclk_i         :   std_logic;
    signal    gt12_rst_i                      : std_logic;
signal   gt13_qpllclk_i            :   std_logic;
signal   gt13_qpllrefclk_i         :   std_logic;
    signal    gt13_rst_i                      : std_logic;
signal   gt14_qpllclk_i            :   std_logic;
signal   gt14_qpllrefclk_i         :   std_logic;
    signal    gt14_rst_i                      : std_logic;
signal   gt15_qpllclk_i            :   std_logic;
signal   gt15_qpllrefclk_i         :   std_logic;
    signal    gt15_rst_i                      : std_logic;
signal   gt16_qpllclk_i            :   std_logic;
signal   gt16_qpllrefclk_i         :   std_logic;
    signal    gt16_rst_i                      : std_logic;
signal   gt17_qpllclk_i            :   std_logic;
signal   gt17_qpllrefclk_i         :   std_logic;
    signal    gt17_rst_i                      : std_logic;
signal   gt18_qpllclk_i            :   std_logic;
signal   gt18_qpllrefclk_i         :   std_logic;
    signal    gt18_rst_i                      : std_logic;
signal   gt19_qpllclk_i            :   std_logic;
signal   gt19_qpllrefclk_i         :   std_logic;
    signal    gt19_rst_i                      : std_logic;
signal   gt20_qpllclk_i            :   std_logic;
signal   gt20_qpllrefclk_i         :   std_logic;
    signal    gt20_rst_i                      : std_logic;
signal   gt21_qpllclk_i            :   std_logic;
signal   gt21_qpllrefclk_i         :   std_logic;
    signal    gt21_rst_i                      : std_logic;
signal   gt22_qpllclk_i            :   std_logic;
signal   gt22_qpllrefclk_i         :   std_logic;
    signal    gt22_rst_i                      : std_logic;
signal   gt23_qpllclk_i            :   std_logic;
signal   gt23_qpllrefclk_i         :   std_logic;
    signal    gt23_rst_i                      : std_logic;
signal   gt24_qpllclk_i            :   std_logic;
signal   gt24_qpllrefclk_i         :   std_logic;
    signal    gt24_rst_i                      : std_logic;
signal   gt25_qpllclk_i            :   std_logic;
signal   gt25_qpllrefclk_i         :   std_logic;
    signal    gt25_rst_i                      : std_logic;
signal   gt26_qpllclk_i            :   std_logic;
signal   gt26_qpllrefclk_i         :   std_logic;
    signal    gt26_rst_i                      : std_logic;
signal   gt27_qpllclk_i            :   std_logic;
signal   gt27_qpllrefclk_i         :   std_logic;
    signal    gt27_rst_i                      : std_logic;
signal   gt28_qpllclk_i            :   std_logic;
signal   gt28_qpllrefclk_i         :   std_logic;
    signal    gt28_rst_i                      : std_logic;
signal   gt29_qpllclk_i            :   std_logic;
signal   gt29_qpllrefclk_i         :   std_logic;
    signal    gt29_rst_i                      : std_logic;
signal   gt30_qpllclk_i            :   std_logic;
signal   gt30_qpllrefclk_i         :   std_logic;
    signal    gt30_rst_i                      : std_logic;
signal   gt31_qpllclk_i            :   std_logic;
signal   gt31_qpllrefclk_i         :   std_logic;
    signal    gt31_rst_i                      : std_logic;
    signal   gt0_cpllreset_i            :   std_logic;
    signal   gt0_cpllpd_i         :   std_logic;
    signal   gt1_cpllreset_i            :   std_logic;
    signal   gt1_cpllpd_i         :   std_logic;
    signal   gt2_cpllreset_i            :   std_logic;
    signal   gt2_cpllpd_i         :   std_logic;
    signal   gt3_cpllreset_i            :   std_logic;
    signal   gt3_cpllpd_i         :   std_logic;
    signal   gt4_cpllreset_i            :   std_logic;
    signal   gt4_cpllpd_i         :   std_logic;
    signal   gt5_cpllreset_i            :   std_logic;
    signal   gt5_cpllpd_i         :   std_logic;
    signal   gt6_cpllreset_i            :   std_logic;
    signal   gt6_cpllpd_i         :   std_logic;
    signal   gt7_cpllreset_i            :   std_logic;
    signal   gt7_cpllpd_i         :   std_logic;
    signal   gt8_cpllreset_i            :   std_logic;
    signal   gt8_cpllpd_i         :   std_logic;
    signal   gt9_cpllreset_i            :   std_logic;
    signal   gt9_cpllpd_i         :   std_logic;
    signal   gt10_cpllreset_i            :   std_logic;
    signal   gt10_cpllpd_i         :   std_logic;
    signal   gt11_cpllreset_i            :   std_logic;
    signal   gt11_cpllpd_i         :   std_logic;
    signal   gt12_cpllreset_i            :   std_logic;
    signal   gt12_cpllpd_i         :   std_logic;
    signal   gt13_cpllreset_i            :   std_logic;
    signal   gt13_cpllpd_i         :   std_logic;
    signal   gt14_cpllreset_i            :   std_logic;
    signal   gt14_cpllpd_i         :   std_logic;
    signal   gt15_cpllreset_i            :   std_logic;
    signal   gt15_cpllpd_i         :   std_logic;
    signal   gt16_cpllreset_i            :   std_logic;
    signal   gt16_cpllpd_i         :   std_logic;
    signal   gt17_cpllreset_i            :   std_logic;
    signal   gt17_cpllpd_i         :   std_logic;
    signal   gt18_cpllreset_i            :   std_logic;
    signal   gt18_cpllpd_i         :   std_logic;
    signal   gt19_cpllreset_i            :   std_logic;
    signal   gt19_cpllpd_i         :   std_logic;
    signal   gt20_cpllreset_i            :   std_logic;
    signal   gt20_cpllpd_i         :   std_logic;
    signal   gt21_cpllreset_i            :   std_logic;
    signal   gt21_cpllpd_i         :   std_logic;
    signal   gt22_cpllreset_i            :   std_logic;
    signal   gt22_cpllpd_i         :   std_logic;
    signal   gt23_cpllreset_i            :   std_logic;
    signal   gt23_cpllpd_i         :   std_logic;
    signal   gt24_cpllreset_i            :   std_logic;
    signal   gt24_cpllpd_i         :   std_logic;
    signal   gt25_cpllreset_i            :   std_logic;
    signal   gt25_cpllpd_i         :   std_logic;
    signal   gt26_cpllreset_i            :   std_logic;
    signal   gt26_cpllpd_i         :   std_logic;
    signal   gt27_cpllreset_i            :   std_logic;
    signal   gt27_cpllpd_i         :   std_logic;
    signal   gt28_cpllreset_i            :   std_logic;
    signal   gt28_cpllpd_i         :   std_logic;
    signal   gt29_cpllreset_i            :   std_logic;
    signal   gt29_cpllpd_i         :   std_logic;
    signal   gt30_cpllreset_i            :   std_logic;
    signal   gt30_cpllpd_i         :   std_logic;
    signal   gt31_cpllreset_i            :   std_logic;
    signal   gt31_cpllpd_i         :   std_logic;


--*************************** Component Declarations **************************
component gtwizard_0_GT
generic
(
    -- Simulation attributes
    GT_SIM_GTRESET_SPEEDUP    : string := "FALSE";
    EXAMPLE_SIMULATION        : integer  := 0;   
    TXSYNC_OVRD_IN            : bit    := '0';
    SIM_CPLLREFCLK_SEL        : bit_vector (2 downto 0) :=   "001";
    TXSYNC_MULTILANE_IN       : bit    := '0'     
);
port 
(   
    RST_IN                                  : in   std_logic;
    DRP_BUSY_OUT                            : out  std_logic;
 RXPMARESETDONE  : out  std_logic;
 TXPMARESETDONE  : out  std_logic;
     cpllrefclksel_in : in std_logic_vector (2 downto 0);
    ---------------------------- Channel - DRP Ports  --------------------------
    drpaddr_in                              : in   std_logic_vector(8 downto 0);
    drpclk_in                               : in   std_logic;
    drpdi_in                                : in   std_logic_vector(15 downto 0);
    drpdo_out                               : out  std_logic_vector(15 downto 0);
    drpen_in                                : in   std_logic;
    drprdy_out                              : out  std_logic;
    drpwe_in                                : in   std_logic;
    ------------------------------- Clocking Ports -----------------------------
    qpllclk_in                              : in   std_logic;
    qpllrefclk_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    eyescanreset_in                         : in   std_logic;
    rxuserrdy_in                            : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    eyescandataerror_out                    : out  std_logic;
    eyescantrigger_in                       : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    rxslide_in                              : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    dmonitorout_out                         : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    rxusrclk_in                             : in   std_logic;
    rxusrclk2_in                            : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    rxdata_out                              : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    rxdisperr_out                           : out  std_logic_vector(7 downto 0);
    rxnotintable_out                        : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gthrxn_in                               : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    rxdlyen_in                              : in   std_logic;
    rxdlysreset_in                          : in   std_logic;
    rxdlysresetdone_out                     : out  std_logic;
    rxphalign_in                            : in   std_logic;
    rxphaligndone_out                       : out  std_logic;
    rxphalignen_in                          : in   std_logic;
    rxphdlyreset_in                         : in   std_logic;
    rxphmonitor_out                         : out  std_logic_vector(4 downto 0);
    rxphslipmonitor_out                     : out  std_logic_vector(4 downto 0);
    rxsyncallin_in                          : in   std_logic;
    rxsyncdone_out                          : out  std_logic;
    rxsyncin_in                             : in   std_logic;
    rxsyncmode_in                           : in   std_logic;
    rxsyncout_out                           : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    rxbyteisaligned_out                     : out  std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    rxlpmhfhold_in                          : in   std_logic;
    rxlpmlfhold_in                          : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    rxmonitorout_out                        : out  std_logic_vector(6 downto 0);
    rxmonitorsel_in                         : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    rxoutclk_out                            : out  std_logic;
    rxoutclkfabric_out                      : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gtrxreset_in                            : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    rxcharisk_out                           : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gthrxp_in                               : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    rxresetdone_out                         : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gttxreset_in                            : in   std_logic;
    txuserrdy_in                            : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    txusrclk_in                             : in   std_logic;
    txusrclk2_in                            : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    txdlyen_in                              : in   std_logic;
    txdlysreset_in                          : in   std_logic;
    txdlysresetdone_out                     : out  std_logic;
    txphalign_in                            : in   std_logic;
    txphaligndone_out                       : out  std_logic;
    txphalignen_in                          : in   std_logic;
    txphdlyreset_in                         : in   std_logic;
    txphinit_in                             : in   std_logic;
    txphinitdone_out                        : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    txdata_in                               : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gthtxn_out                              : out  std_logic;
    gthtxp_out                              : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    txoutclk_out                            : out  std_logic;
    txoutclkfabric_out                      : out  std_logic;
    txoutclkpcs_out                         : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    txresetdone_out                         : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    txcharisk_in                            : in   std_logic_vector(7 downto 0)


);
end component;



--********************************* Main Body of Code**************************

begin                       

    tied_to_ground_i                    <= '0';
    tied_to_ground_vec_i(63 downto 0)   <= (others => '0');
    tied_to_vcc_i                       <= '1';
    gt0_qpllclk_i    <= GT0_QPLLOUTCLK_IN;  
    gt0_qpllrefclk_i <= GT0_QPLLOUTREFCLK_IN; 
    gt1_qpllclk_i    <= GT0_QPLLOUTCLK_IN;  
    gt1_qpllrefclk_i <= GT0_QPLLOUTREFCLK_IN; 
    gt2_qpllclk_i    <= GT0_QPLLOUTCLK_IN;  
    gt2_qpllrefclk_i <= GT0_QPLLOUTREFCLK_IN; 
    gt3_qpllclk_i    <= GT0_QPLLOUTCLK_IN;  
    gt3_qpllrefclk_i <= GT0_QPLLOUTREFCLK_IN; 
    gt4_qpllclk_i    <= GT1_QPLLOUTCLK_IN;  
    gt4_qpllrefclk_i <= GT1_QPLLOUTREFCLK_IN; 
    gt5_qpllclk_i    <= GT1_QPLLOUTCLK_IN;  
    gt5_qpllrefclk_i <= GT1_QPLLOUTREFCLK_IN; 
    gt6_qpllclk_i    <= GT1_QPLLOUTCLK_IN;  
    gt6_qpllrefclk_i <= GT1_QPLLOUTREFCLK_IN; 
    gt7_qpllclk_i    <= GT1_QPLLOUTCLK_IN;  
    gt7_qpllrefclk_i <= GT1_QPLLOUTREFCLK_IN; 
    gt8_qpllclk_i    <= GT2_QPLLOUTCLK_IN;  
    gt8_qpllrefclk_i <= GT2_QPLLOUTREFCLK_IN; 
    gt9_qpllclk_i    <= GT2_QPLLOUTCLK_IN;  
    gt9_qpllrefclk_i <= GT2_QPLLOUTREFCLK_IN; 
    gt10_qpllclk_i    <= GT2_QPLLOUTCLK_IN;  
    gt10_qpllrefclk_i <= GT2_QPLLOUTREFCLK_IN; 
    gt11_qpllclk_i    <= GT2_QPLLOUTCLK_IN;  
    gt11_qpllrefclk_i <= GT2_QPLLOUTREFCLK_IN; 
    gt12_qpllclk_i    <= GT3_QPLLOUTCLK_IN;  
    gt12_qpllrefclk_i <= GT3_QPLLOUTREFCLK_IN; 
    gt13_qpllclk_i    <= GT3_QPLLOUTCLK_IN;  
    gt13_qpllrefclk_i <= GT3_QPLLOUTREFCLK_IN; 
    gt14_qpllclk_i    <= GT3_QPLLOUTCLK_IN;  
    gt14_qpllrefclk_i <= GT3_QPLLOUTREFCLK_IN; 
    gt15_qpllclk_i    <= GT3_QPLLOUTCLK_IN;  
    gt15_qpllrefclk_i <= GT3_QPLLOUTREFCLK_IN; 
    gt16_qpllclk_i    <= GT4_QPLLOUTCLK_IN;  
    gt16_qpllrefclk_i <= GT4_QPLLOUTREFCLK_IN; 
    gt17_qpllclk_i    <= GT4_QPLLOUTCLK_IN;  
    gt17_qpllrefclk_i <= GT4_QPLLOUTREFCLK_IN; 
    gt18_qpllclk_i    <= GT4_QPLLOUTCLK_IN;  
    gt18_qpllrefclk_i <= GT4_QPLLOUTREFCLK_IN; 
    gt19_qpllclk_i    <= GT4_QPLLOUTCLK_IN;  
    gt19_qpllrefclk_i <= GT4_QPLLOUTREFCLK_IN; 
    gt20_qpllclk_i    <= GT5_QPLLOUTCLK_IN;  
    gt20_qpllrefclk_i <= GT5_QPLLOUTREFCLK_IN; 
    gt21_qpllclk_i    <= GT5_QPLLOUTCLK_IN;  
    gt21_qpllrefclk_i <= GT5_QPLLOUTREFCLK_IN; 
    gt22_qpllclk_i    <= GT5_QPLLOUTCLK_IN;  
    gt22_qpllrefclk_i <= GT5_QPLLOUTREFCLK_IN; 
    gt23_qpllclk_i    <= GT5_QPLLOUTCLK_IN;  
    gt23_qpllrefclk_i <= GT5_QPLLOUTREFCLK_IN; 
    gt24_qpllclk_i    <= GT6_QPLLOUTCLK_IN;  
    gt24_qpllrefclk_i <= GT6_QPLLOUTREFCLK_IN; 
    gt25_qpllclk_i    <= GT6_QPLLOUTCLK_IN;  
    gt25_qpllrefclk_i <= GT6_QPLLOUTREFCLK_IN; 
    gt26_qpllclk_i    <= GT6_QPLLOUTCLK_IN;  
    gt26_qpllrefclk_i <= GT6_QPLLOUTREFCLK_IN; 
    gt27_qpllclk_i    <= GT6_QPLLOUTCLK_IN;  
    gt27_qpllrefclk_i <= GT6_QPLLOUTREFCLK_IN; 
    gt28_qpllclk_i    <= GT7_QPLLOUTCLK_IN;  
    gt28_qpllrefclk_i <= GT7_QPLLOUTREFCLK_IN; 
    gt29_qpllclk_i    <= GT7_QPLLOUTCLK_IN;  
    gt29_qpllrefclk_i <= GT7_QPLLOUTREFCLK_IN; 
    gt30_qpllclk_i    <= GT7_QPLLOUTCLK_IN;  
    gt30_qpllrefclk_i <= GT7_QPLLOUTREFCLK_IN; 
    gt31_qpllclk_i    <= GT7_QPLLOUTCLK_IN;  
    gt31_qpllrefclk_i <= GT7_QPLLOUTREFCLK_IN; 

      gt0_rst_i        <= GT0_QPLLRESET_IN;
   
      gt1_rst_i        <= GT0_QPLLRESET_IN;
   
      gt2_rst_i        <= GT0_QPLLRESET_IN;
   
      gt3_rst_i        <= GT0_QPLLRESET_IN;
   
      gt4_rst_i        <= GT1_QPLLRESET_IN;
   
      gt5_rst_i        <= GT1_QPLLRESET_IN;
   
      gt6_rst_i        <= GT1_QPLLRESET_IN;
   
      gt7_rst_i        <= GT1_QPLLRESET_IN;
   
      gt8_rst_i        <= GT2_QPLLRESET_IN;
   
      gt9_rst_i        <= GT2_QPLLRESET_IN;
   
      gt10_rst_i        <= GT2_QPLLRESET_IN;
   
      gt11_rst_i        <= GT2_QPLLRESET_IN;
   
      gt12_rst_i        <= GT3_QPLLRESET_IN;
   
      gt13_rst_i        <= GT3_QPLLRESET_IN;
   
      gt14_rst_i        <= GT3_QPLLRESET_IN;
   
      gt15_rst_i        <= GT3_QPLLRESET_IN;
   
      gt16_rst_i        <= GT4_QPLLRESET_IN;
   
      gt17_rst_i        <= GT4_QPLLRESET_IN;
   
      gt18_rst_i        <= GT4_QPLLRESET_IN;
   
      gt19_rst_i        <= GT4_QPLLRESET_IN;
   
      gt20_rst_i        <= GT5_QPLLRESET_IN;
   
      gt21_rst_i        <= GT5_QPLLRESET_IN;
   
      gt22_rst_i        <= GT5_QPLLRESET_IN;
   
      gt23_rst_i        <= GT5_QPLLRESET_IN;
   
      gt24_rst_i        <= GT6_QPLLRESET_IN;
   
      gt25_rst_i        <= GT6_QPLLRESET_IN;
   
      gt26_rst_i        <= GT6_QPLLRESET_IN;
   
      gt27_rst_i        <= GT6_QPLLRESET_IN;
   
      gt28_rst_i        <= GT7_QPLLRESET_IN;
   
      gt29_rst_i        <= GT7_QPLLRESET_IN;
   
      gt30_rst_i        <= GT7_QPLLRESET_IN;
   
      gt31_rst_i        <= GT7_QPLLRESET_IN;
   
     

    --------------------------- GT Instances  -------------------------------   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT0  (X0Y4)
gt0_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_OVRD_IN         => ('1'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt0_rst_i,
        DRP_BUSY_OUT                    =>      GT0_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT0_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT0_TXPMARESETDONE_OUT,
        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt0_drpaddr_in,
        drpclk_in                       =>      gt0_drpclk_in,
        drpdi_in                        =>      gt0_drpdi_in,
        drpdo_out                       =>      gt0_drpdo_out,
        drpen_in                        =>      gt0_drpen_in,
        drprdy_out                      =>      gt0_drprdy_out,
        drpwe_in                        =>      gt0_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt0_qpllclk_i,
        qpllrefclk_in                   =>      gt0_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt0_eyescanreset_in,
        rxuserrdy_in                    =>      gt0_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt0_eyescandataerror_out,
        eyescantrigger_in               =>      gt0_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt0_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt0_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt0_rxusrclk_in,
        rxusrclk2_in                    =>      gt0_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt0_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt0_rxdisperr_out,
        rxnotintable_out                =>      gt0_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt0_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt0_rxdlyen_in,
        rxdlysreset_in                  =>      gt0_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt0_rxdlysresetdone_out,
        rxphalign_in                    =>      gt0_rxphalign_in,
        rxphaligndone_out               =>      gt0_rxphaligndone_out,
        rxphalignen_in                  =>      gt0_rxphalignen_in,
        rxphdlyreset_in                 =>      gt0_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt0_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt0_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt0_rxsyncallin_in,
        rxsyncdone_out                  =>      gt0_rxsyncdone_out,
        rxsyncin_in                     =>      gt0_rxsyncin_in,
        rxsyncmode_in                   =>      gt0_rxsyncmode_in,
        rxsyncout_out                   =>      gt0_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt0_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt0_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt0_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt0_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt0_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt0_rxoutclk_out,
        rxoutclkfabric_out              =>      gt0_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt0_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt0_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt0_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt0_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt0_gttxreset_in,
        txuserrdy_in                    =>      gt0_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt0_txusrclk_in,
        txusrclk2_in                    =>      gt0_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt0_txdlyen_in,
        txdlysreset_in                  =>      gt0_txdlysreset_in,
        txdlysresetdone_out             =>      gt0_txdlysresetdone_out,
        txphalign_in                    =>      gt0_txphalign_in,
        txphaligndone_out               =>      gt0_txphaligndone_out,
        txphalignen_in                  =>      gt0_txphalignen_in,
        txphdlyreset_in                 =>      gt0_txphdlyreset_in,
        txphinit_in                     =>      gt0_txphinit_in,
        txphinitdone_out                =>      gt0_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt0_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt0_gthtxn_out,
        gthtxp_out                      =>      gt0_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt0_txoutclk_out,
        txoutclkfabric_out              =>      gt0_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt0_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt0_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt0_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT1  (X0Y5)
gt1_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt1_rst_i,
        DRP_BUSY_OUT                    =>      GT1_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT1_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT1_TXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt1_drpaddr_in,
        drpclk_in                       =>      gt1_drpclk_in,
        drpdi_in                        =>      gt1_drpdi_in,
        drpdo_out                       =>      gt1_drpdo_out,
        drpen_in                        =>      gt1_drpen_in,
        drprdy_out                      =>      gt1_drprdy_out,
        drpwe_in                        =>      gt1_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt1_qpllclk_i,
        qpllrefclk_in                   =>      gt1_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt1_eyescanreset_in,
        rxuserrdy_in                    =>      gt1_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt1_eyescandataerror_out,
        eyescantrigger_in               =>      gt1_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt1_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt1_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt1_rxusrclk_in,
        rxusrclk2_in                    =>      gt1_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt1_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt1_rxdisperr_out,
        rxnotintable_out                =>      gt1_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt1_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt1_rxdlyen_in,
        rxdlysreset_in                  =>      gt1_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt1_rxdlysresetdone_out,
        rxphalign_in                    =>      gt1_rxphalign_in,
        rxphaligndone_out               =>      gt1_rxphaligndone_out,
        rxphalignen_in                  =>      gt1_rxphalignen_in,
        rxphdlyreset_in                 =>      gt1_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt1_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt1_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt1_rxsyncallin_in,
        rxsyncdone_out                  =>      gt1_rxsyncdone_out,
        rxsyncin_in                     =>      gt1_rxsyncin_in,
        rxsyncmode_in                   =>      gt1_rxsyncmode_in,
        rxsyncout_out                   =>      gt1_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt1_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt1_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt1_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt1_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt1_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt1_rxoutclk_out,
        rxoutclkfabric_out              =>      gt1_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt1_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt1_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt1_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt1_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt1_gttxreset_in,
        txuserrdy_in                    =>      gt1_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt1_txusrclk_in,
        txusrclk2_in                    =>      gt1_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt1_txdlyen_in,
        txdlysreset_in                  =>      gt1_txdlysreset_in,
        txdlysresetdone_out             =>      gt1_txdlysresetdone_out,
        txphalign_in                    =>      gt1_txphalign_in,
        txphaligndone_out               =>      gt1_txphaligndone_out,
        txphalignen_in                  =>      gt1_txphalignen_in,
        txphdlyreset_in                 =>      gt1_txphdlyreset_in,
        txphinit_in                     =>      gt1_txphinit_in,
        txphinitdone_out                =>      gt1_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt1_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt1_gthtxn_out,
        gthtxp_out                      =>      gt1_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt1_txoutclk_out,
        txoutclkfabric_out              =>      gt1_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt1_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt1_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt1_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT2  (X0Y6)
gt2_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt2_rst_i,
        DRP_BUSY_OUT                    =>      GT2_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT2_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT2_TXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt2_drpaddr_in,
        drpclk_in                       =>      gt2_drpclk_in,
        drpdi_in                        =>      gt2_drpdi_in,
        drpdo_out                       =>      gt2_drpdo_out,
        drpen_in                        =>      gt2_drpen_in,
        drprdy_out                      =>      gt2_drprdy_out,
        drpwe_in                        =>      gt2_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt2_qpllclk_i,
        qpllrefclk_in                   =>      gt2_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt2_eyescanreset_in,
        rxuserrdy_in                    =>      gt2_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt2_eyescandataerror_out,
        eyescantrigger_in               =>      gt2_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt2_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt2_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt2_rxusrclk_in,
        rxusrclk2_in                    =>      gt2_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt2_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt2_rxdisperr_out,
        rxnotintable_out                =>      gt2_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt2_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt2_rxdlyen_in,
        rxdlysreset_in                  =>      gt2_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt2_rxdlysresetdone_out,
        rxphalign_in                    =>      gt2_rxphalign_in,
        rxphaligndone_out               =>      gt2_rxphaligndone_out,
        rxphalignen_in                  =>      gt2_rxphalignen_in,
        rxphdlyreset_in                 =>      gt2_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt2_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt2_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt2_rxsyncallin_in,
        rxsyncdone_out                  =>      gt2_rxsyncdone_out,
        rxsyncin_in                     =>      gt2_rxsyncin_in,
        rxsyncmode_in                   =>      gt2_rxsyncmode_in,
        rxsyncout_out                   =>      gt2_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt2_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt2_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt2_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt2_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt2_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt2_rxoutclk_out,
        rxoutclkfabric_out              =>      gt2_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt2_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt2_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt2_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt2_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt2_gttxreset_in,
        txuserrdy_in                    =>      gt2_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt2_txusrclk_in,
        txusrclk2_in                    =>      gt2_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt2_txdlyen_in,
        txdlysreset_in                  =>      gt2_txdlysreset_in,
        txdlysresetdone_out             =>      gt2_txdlysresetdone_out,
        txphalign_in                    =>      gt2_txphalign_in,
        txphaligndone_out               =>      gt2_txphaligndone_out,
        txphalignen_in                  =>      gt2_txphalignen_in,
        txphdlyreset_in                 =>      gt2_txphdlyreset_in,
        txphinit_in                     =>      gt2_txphinit_in,
        txphinitdone_out                =>      gt2_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt2_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt2_gthtxn_out,
        gthtxp_out                      =>      gt2_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt2_txoutclk_out,
        txoutclkfabric_out              =>      gt2_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt2_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt2_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt2_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT3  (X0Y7)
gt3_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt3_rst_i,
        DRP_BUSY_OUT                    =>      GT3_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT3_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT3_TXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt3_drpaddr_in,
        drpclk_in                       =>      gt3_drpclk_in,
        drpdi_in                        =>      gt3_drpdi_in,
        drpdo_out                       =>      gt3_drpdo_out,
        drpen_in                        =>      gt3_drpen_in,
        drprdy_out                      =>      gt3_drprdy_out,
        drpwe_in                        =>      gt3_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt3_qpllclk_i,
        qpllrefclk_in                   =>      gt3_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt3_eyescanreset_in,
        rxuserrdy_in                    =>      gt3_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt3_eyescandataerror_out,
        eyescantrigger_in               =>      gt3_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt3_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt3_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt3_rxusrclk_in,
        rxusrclk2_in                    =>      gt3_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt3_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt3_rxdisperr_out,
        rxnotintable_out                =>      gt3_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt3_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt3_rxdlyen_in,
        rxdlysreset_in                  =>      gt3_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt3_rxdlysresetdone_out,
        rxphalign_in                    =>      gt3_rxphalign_in,
        rxphaligndone_out               =>      gt3_rxphaligndone_out,
        rxphalignen_in                  =>      gt3_rxphalignen_in,
        rxphdlyreset_in                 =>      gt3_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt3_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt3_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt3_rxsyncallin_in,
        rxsyncdone_out                  =>      gt3_rxsyncdone_out,
        rxsyncin_in                     =>      gt3_rxsyncin_in,
        rxsyncmode_in                   =>      gt3_rxsyncmode_in,
        rxsyncout_out                   =>      gt3_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt3_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt3_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt3_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt3_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt3_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt3_rxoutclk_out,
        rxoutclkfabric_out              =>      gt3_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt3_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt3_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt3_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt3_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt3_gttxreset_in,
        txuserrdy_in                    =>      gt3_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt3_txusrclk_in,
        txusrclk2_in                    =>      gt3_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt3_txdlyen_in,
        txdlysreset_in                  =>      gt3_txdlysreset_in,
        txdlysresetdone_out             =>      gt3_txdlysresetdone_out,
        txphalign_in                    =>      gt3_txphalign_in,
        txphaligndone_out               =>      gt3_txphaligndone_out,
        txphalignen_in                  =>      gt3_txphalignen_in,
        txphdlyreset_in                 =>      gt3_txphdlyreset_in,
        txphinit_in                     =>      gt3_txphinit_in,
        txphinitdone_out                =>      gt3_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt3_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt3_gthtxn_out,
        gthtxp_out                      =>      gt3_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt3_txoutclk_out,
        txoutclkfabric_out              =>      gt3_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt3_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt3_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt3_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT4  (X0Y8)
gt4_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt4_rst_i,
        DRP_BUSY_OUT                    =>      GT4_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT4_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT4_TXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt4_drpaddr_in,
        drpclk_in                       =>      gt4_drpclk_in,
        drpdi_in                        =>      gt4_drpdi_in,
        drpdo_out                       =>      gt4_drpdo_out,
        drpen_in                        =>      gt4_drpen_in,
        drprdy_out                      =>      gt4_drprdy_out,
        drpwe_in                        =>      gt4_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt4_qpllclk_i,
        qpllrefclk_in                   =>      gt4_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt4_eyescanreset_in,
        rxuserrdy_in                    =>      gt4_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt4_eyescandataerror_out,
        eyescantrigger_in               =>      gt4_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt4_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt4_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt4_rxusrclk_in,
        rxusrclk2_in                    =>      gt4_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt4_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt4_rxdisperr_out,
        rxnotintable_out                =>      gt4_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt4_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt4_rxdlyen_in,
        rxdlysreset_in                  =>      gt4_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt4_rxdlysresetdone_out,
        rxphalign_in                    =>      gt4_rxphalign_in,
        rxphaligndone_out               =>      gt4_rxphaligndone_out,
        rxphalignen_in                  =>      gt4_rxphalignen_in,
        rxphdlyreset_in                 =>      gt4_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt4_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt4_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt4_rxsyncallin_in,
        rxsyncdone_out                  =>      gt4_rxsyncdone_out,
        rxsyncin_in                     =>      gt4_rxsyncin_in,
        rxsyncmode_in                   =>      gt4_rxsyncmode_in,
        rxsyncout_out                   =>      gt4_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt4_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt4_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt4_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt4_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt4_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt4_rxoutclk_out,
        rxoutclkfabric_out              =>      gt4_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt4_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt4_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt4_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt4_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt4_gttxreset_in,
        txuserrdy_in                    =>      gt4_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt4_txusrclk_in,
        txusrclk2_in                    =>      gt4_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt4_txdlyen_in,
        txdlysreset_in                  =>      gt4_txdlysreset_in,
        txdlysresetdone_out             =>      gt4_txdlysresetdone_out,
        txphalign_in                    =>      gt4_txphalign_in,
        txphaligndone_out               =>      gt4_txphaligndone_out,
        txphalignen_in                  =>      gt4_txphalignen_in,
        txphdlyreset_in                 =>      gt4_txphdlyreset_in,
        txphinit_in                     =>      gt4_txphinit_in,
        txphinitdone_out                =>      gt4_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt4_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt4_gthtxn_out,
        gthtxp_out                      =>      gt4_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt4_txoutclk_out,
        txoutclkfabric_out              =>      gt4_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt4_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt4_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt4_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT5  (X0Y9)
gt5_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt5_rst_i,
        DRP_BUSY_OUT                    =>      GT5_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT5_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT5_TXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt5_drpaddr_in,
        drpclk_in                       =>      gt5_drpclk_in,
        drpdi_in                        =>      gt5_drpdi_in,
        drpdo_out                       =>      gt5_drpdo_out,
        drpen_in                        =>      gt5_drpen_in,
        drprdy_out                      =>      gt5_drprdy_out,
        drpwe_in                        =>      gt5_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt5_qpllclk_i,
        qpllrefclk_in                   =>      gt5_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt5_eyescanreset_in,
        rxuserrdy_in                    =>      gt5_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt5_eyescandataerror_out,
        eyescantrigger_in               =>      gt5_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt5_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt5_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt5_rxusrclk_in,
        rxusrclk2_in                    =>      gt5_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt5_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt5_rxdisperr_out,
        rxnotintable_out                =>      gt5_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt5_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt5_rxdlyen_in,
        rxdlysreset_in                  =>      gt5_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt5_rxdlysresetdone_out,
        rxphalign_in                    =>      gt5_rxphalign_in,
        rxphaligndone_out               =>      gt5_rxphaligndone_out,
        rxphalignen_in                  =>      gt5_rxphalignen_in,
        rxphdlyreset_in                 =>      gt5_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt5_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt5_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt5_rxsyncallin_in,
        rxsyncdone_out                  =>      gt5_rxsyncdone_out,
        rxsyncin_in                     =>      gt5_rxsyncin_in,
        rxsyncmode_in                   =>      gt5_rxsyncmode_in,
        rxsyncout_out                   =>      gt5_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt5_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt5_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt5_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt5_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt5_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt5_rxoutclk_out,
        rxoutclkfabric_out              =>      gt5_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt5_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt5_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt5_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt5_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt5_gttxreset_in,
        txuserrdy_in                    =>      gt5_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt5_txusrclk_in,
        txusrclk2_in                    =>      gt5_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt5_txdlyen_in,
        txdlysreset_in                  =>      gt5_txdlysreset_in,
        txdlysresetdone_out             =>      gt5_txdlysresetdone_out,
        txphalign_in                    =>      gt5_txphalign_in,
        txphaligndone_out               =>      gt5_txphaligndone_out,
        txphalignen_in                  =>      gt5_txphalignen_in,
        txphdlyreset_in                 =>      gt5_txphdlyreset_in,
        txphinit_in                     =>      gt5_txphinit_in,
        txphinitdone_out                =>      gt5_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt5_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt5_gthtxn_out,
        gthtxp_out                      =>      gt5_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt5_txoutclk_out,
        txoutclkfabric_out              =>      gt5_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt5_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt5_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt5_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT6  (X0Y10)
gt6_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt6_rst_i,
        DRP_BUSY_OUT                    =>      GT6_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT6_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT6_TXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt6_drpaddr_in,
        drpclk_in                       =>      gt6_drpclk_in,
        drpdi_in                        =>      gt6_drpdi_in,
        drpdo_out                       =>      gt6_drpdo_out,
        drpen_in                        =>      gt6_drpen_in,
        drprdy_out                      =>      gt6_drprdy_out,
        drpwe_in                        =>      gt6_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt6_qpllclk_i,
        qpllrefclk_in                   =>      gt6_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt6_eyescanreset_in,
        rxuserrdy_in                    =>      gt6_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt6_eyescandataerror_out,
        eyescantrigger_in               =>      gt6_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt6_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt6_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt6_rxusrclk_in,
        rxusrclk2_in                    =>      gt6_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt6_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt6_rxdisperr_out,
        rxnotintable_out                =>      gt6_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt6_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt6_rxdlyen_in,
        rxdlysreset_in                  =>      gt6_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt6_rxdlysresetdone_out,
        rxphalign_in                    =>      gt6_rxphalign_in,
        rxphaligndone_out               =>      gt6_rxphaligndone_out,
        rxphalignen_in                  =>      gt6_rxphalignen_in,
        rxphdlyreset_in                 =>      gt6_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt6_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt6_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt6_rxsyncallin_in,
        rxsyncdone_out                  =>      gt6_rxsyncdone_out,
        rxsyncin_in                     =>      gt6_rxsyncin_in,
        rxsyncmode_in                   =>      gt6_rxsyncmode_in,
        rxsyncout_out                   =>      gt6_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt6_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt6_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt6_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt6_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt6_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt6_rxoutclk_out,
        rxoutclkfabric_out              =>      gt6_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt6_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt6_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt6_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt6_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt6_gttxreset_in,
        txuserrdy_in                    =>      gt6_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt6_txusrclk_in,
        txusrclk2_in                    =>      gt6_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt6_txdlyen_in,
        txdlysreset_in                  =>      gt6_txdlysreset_in,
        txdlysresetdone_out             =>      gt6_txdlysresetdone_out,
        txphalign_in                    =>      gt6_txphalign_in,
        txphaligndone_out               =>      gt6_txphaligndone_out,
        txphalignen_in                  =>      gt6_txphalignen_in,
        txphdlyreset_in                 =>      gt6_txphdlyreset_in,
        txphinit_in                     =>      gt6_txphinit_in,
        txphinitdone_out                =>      gt6_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt6_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt6_gthtxn_out,
        gthtxp_out                      =>      gt6_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt6_txoutclk_out,
        txoutclkfabric_out              =>      gt6_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt6_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt6_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt6_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT7  (X0Y11)
gt7_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt7_rst_i,
        DRP_BUSY_OUT                    =>      GT7_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT7_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT7_TXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt7_drpaddr_in,
        drpclk_in                       =>      gt7_drpclk_in,
        drpdi_in                        =>      gt7_drpdi_in,
        drpdo_out                       =>      gt7_drpdo_out,
        drpen_in                        =>      gt7_drpen_in,
        drprdy_out                      =>      gt7_drprdy_out,
        drpwe_in                        =>      gt7_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt7_qpllclk_i,
        qpllrefclk_in                   =>      gt7_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt7_eyescanreset_in,
        rxuserrdy_in                    =>      gt7_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt7_eyescandataerror_out,
        eyescantrigger_in               =>      gt7_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt7_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt7_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt7_rxusrclk_in,
        rxusrclk2_in                    =>      gt7_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt7_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt7_rxdisperr_out,
        rxnotintable_out                =>      gt7_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt7_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt7_rxdlyen_in,
        rxdlysreset_in                  =>      gt7_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt7_rxdlysresetdone_out,
        rxphalign_in                    =>      gt7_rxphalign_in,
        rxphaligndone_out               =>      gt7_rxphaligndone_out,
        rxphalignen_in                  =>      gt7_rxphalignen_in,
        rxphdlyreset_in                 =>      gt7_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt7_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt7_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt7_rxsyncallin_in,
        rxsyncdone_out                  =>      gt7_rxsyncdone_out,
        rxsyncin_in                     =>      gt7_rxsyncin_in,
        rxsyncmode_in                   =>      gt7_rxsyncmode_in,
        rxsyncout_out                   =>      gt7_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt7_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt7_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt7_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt7_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt7_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt7_rxoutclk_out,
        rxoutclkfabric_out              =>      gt7_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt7_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt7_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt7_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt7_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt7_gttxreset_in,
        txuserrdy_in                    =>      gt7_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt7_txusrclk_in,
        txusrclk2_in                    =>      gt7_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt7_txdlyen_in,
        txdlysreset_in                  =>      gt7_txdlysreset_in,
        txdlysresetdone_out             =>      gt7_txdlysresetdone_out,
        txphalign_in                    =>      gt7_txphalign_in,
        txphaligndone_out               =>      gt7_txphaligndone_out,
        txphalignen_in                  =>      gt7_txphalignen_in,
        txphdlyreset_in                 =>      gt7_txphdlyreset_in,
        txphinit_in                     =>      gt7_txphinit_in,
        txphinitdone_out                =>      gt7_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt7_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt7_gthtxn_out,
        gthtxp_out                      =>      gt7_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt7_txoutclk_out,
        txoutclkfabric_out              =>      gt7_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt7_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt7_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt7_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT8  (X0Y12)
gt8_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt8_rst_i,
        DRP_BUSY_OUT                    =>      GT8_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT8_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT8_TXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt8_drpaddr_in,
        drpclk_in                       =>      gt8_drpclk_in,
        drpdi_in                        =>      gt8_drpdi_in,
        drpdo_out                       =>      gt8_drpdo_out,
        drpen_in                        =>      gt8_drpen_in,
        drprdy_out                      =>      gt8_drprdy_out,
        drpwe_in                        =>      gt8_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt8_qpllclk_i,
        qpllrefclk_in                   =>      gt8_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt8_eyescanreset_in,
        rxuserrdy_in                    =>      gt8_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt8_eyescandataerror_out,
        eyescantrigger_in               =>      gt8_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt8_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt8_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt8_rxusrclk_in,
        rxusrclk2_in                    =>      gt8_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt8_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt8_rxdisperr_out,
        rxnotintable_out                =>      gt8_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt8_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt8_rxdlyen_in,
        rxdlysreset_in                  =>      gt8_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt8_rxdlysresetdone_out,
        rxphalign_in                    =>      gt8_rxphalign_in,
        rxphaligndone_out               =>      gt8_rxphaligndone_out,
        rxphalignen_in                  =>      gt8_rxphalignen_in,
        rxphdlyreset_in                 =>      gt8_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt8_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt8_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt8_rxsyncallin_in,
        rxsyncdone_out                  =>      gt8_rxsyncdone_out,
        rxsyncin_in                     =>      gt8_rxsyncin_in,
        rxsyncmode_in                   =>      gt8_rxsyncmode_in,
        rxsyncout_out                   =>      gt8_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt8_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt8_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt8_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt8_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt8_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt8_rxoutclk_out,
        rxoutclkfabric_out              =>      gt8_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt8_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt8_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt8_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt8_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt8_gttxreset_in,
        txuserrdy_in                    =>      gt8_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt8_txusrclk_in,
        txusrclk2_in                    =>      gt8_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt8_txdlyen_in,
        txdlysreset_in                  =>      gt8_txdlysreset_in,
        txdlysresetdone_out             =>      gt8_txdlysresetdone_out,
        txphalign_in                    =>      gt8_txphalign_in,
        txphaligndone_out               =>      gt8_txphaligndone_out,
        txphalignen_in                  =>      gt8_txphalignen_in,
        txphdlyreset_in                 =>      gt8_txphdlyreset_in,
        txphinit_in                     =>      gt8_txphinit_in,
        txphinitdone_out                =>      gt8_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt8_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt8_gthtxn_out,
        gthtxp_out                      =>      gt8_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt8_txoutclk_out,
        txoutclkfabric_out              =>      gt8_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt8_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt8_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt8_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT9  (X0Y13)
gt9_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt9_rst_i,
        DRP_BUSY_OUT                    =>      GT9_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT9_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT9_TXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt9_drpaddr_in,
        drpclk_in                       =>      gt9_drpclk_in,
        drpdi_in                        =>      gt9_drpdi_in,
        drpdo_out                       =>      gt9_drpdo_out,
        drpen_in                        =>      gt9_drpen_in,
        drprdy_out                      =>      gt9_drprdy_out,
        drpwe_in                        =>      gt9_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt9_qpllclk_i,
        qpllrefclk_in                   =>      gt9_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt9_eyescanreset_in,
        rxuserrdy_in                    =>      gt9_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt9_eyescandataerror_out,
        eyescantrigger_in               =>      gt9_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt9_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt9_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt9_rxusrclk_in,
        rxusrclk2_in                    =>      gt9_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt9_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt9_rxdisperr_out,
        rxnotintable_out                =>      gt9_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt9_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt9_rxdlyen_in,
        rxdlysreset_in                  =>      gt9_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt9_rxdlysresetdone_out,
        rxphalign_in                    =>      gt9_rxphalign_in,
        rxphaligndone_out               =>      gt9_rxphaligndone_out,
        rxphalignen_in                  =>      gt9_rxphalignen_in,
        rxphdlyreset_in                 =>      gt9_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt9_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt9_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt9_rxsyncallin_in,
        rxsyncdone_out                  =>      gt9_rxsyncdone_out,
        rxsyncin_in                     =>      gt9_rxsyncin_in,
        rxsyncmode_in                   =>      gt9_rxsyncmode_in,
        rxsyncout_out                   =>      gt9_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt9_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt9_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt9_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt9_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt9_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt9_rxoutclk_out,
        rxoutclkfabric_out              =>      gt9_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt9_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt9_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt9_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt9_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt9_gttxreset_in,
        txuserrdy_in                    =>      gt9_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt9_txusrclk_in,
        txusrclk2_in                    =>      gt9_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt9_txdlyen_in,
        txdlysreset_in                  =>      gt9_txdlysreset_in,
        txdlysresetdone_out             =>      gt9_txdlysresetdone_out,
        txphalign_in                    =>      gt9_txphalign_in,
        txphaligndone_out               =>      gt9_txphaligndone_out,
        txphalignen_in                  =>      gt9_txphalignen_in,
        txphdlyreset_in                 =>      gt9_txphdlyreset_in,
        txphinit_in                     =>      gt9_txphinit_in,
        txphinitdone_out                =>      gt9_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt9_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt9_gthtxn_out,
        gthtxp_out                      =>      gt9_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt9_txoutclk_out,
        txoutclkfabric_out              =>      gt9_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt9_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt9_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt9_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT10  (X0Y14)
gt10_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt10_rst_i,
        DRP_BUSY_OUT                    =>      GT10_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT10_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT10_TXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt10_drpaddr_in,
        drpclk_in                       =>      gt10_drpclk_in,
        drpdi_in                        =>      gt10_drpdi_in,
        drpdo_out                       =>      gt10_drpdo_out,
        drpen_in                        =>      gt10_drpen_in,
        drprdy_out                      =>      gt10_drprdy_out,
        drpwe_in                        =>      gt10_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt10_qpllclk_i,
        qpllrefclk_in                   =>      gt10_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt10_eyescanreset_in,
        rxuserrdy_in                    =>      gt10_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt10_eyescandataerror_out,
        eyescantrigger_in               =>      gt10_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt10_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt10_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt10_rxusrclk_in,
        rxusrclk2_in                    =>      gt10_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt10_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt10_rxdisperr_out,
        rxnotintable_out                =>      gt10_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt10_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt10_rxdlyen_in,
        rxdlysreset_in                  =>      gt10_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt10_rxdlysresetdone_out,
        rxphalign_in                    =>      gt10_rxphalign_in,
        rxphaligndone_out               =>      gt10_rxphaligndone_out,
        rxphalignen_in                  =>      gt10_rxphalignen_in,
        rxphdlyreset_in                 =>      gt10_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt10_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt10_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt10_rxsyncallin_in,
        rxsyncdone_out                  =>      gt10_rxsyncdone_out,
        rxsyncin_in                     =>      gt10_rxsyncin_in,
        rxsyncmode_in                   =>      gt10_rxsyncmode_in,
        rxsyncout_out                   =>      gt10_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt10_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt10_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt10_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt10_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt10_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt10_rxoutclk_out,
        rxoutclkfabric_out              =>      gt10_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt10_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt10_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt10_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt10_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt10_gttxreset_in,
        txuserrdy_in                    =>      gt10_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt10_txusrclk_in,
        txusrclk2_in                    =>      gt10_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt10_txdlyen_in,
        txdlysreset_in                  =>      gt10_txdlysreset_in,
        txdlysresetdone_out             =>      gt10_txdlysresetdone_out,
        txphalign_in                    =>      gt10_txphalign_in,
        txphaligndone_out               =>      gt10_txphaligndone_out,
        txphalignen_in                  =>      gt10_txphalignen_in,
        txphdlyreset_in                 =>      gt10_txphdlyreset_in,
        txphinit_in                     =>      gt10_txphinit_in,
        txphinitdone_out                =>      gt10_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt10_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt10_gthtxn_out,
        gthtxp_out                      =>      gt10_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt10_txoutclk_out,
        txoutclkfabric_out              =>      gt10_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt10_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt10_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt10_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT11  (X0Y15)
gt11_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt11_rst_i,
        DRP_BUSY_OUT                    =>      GT11_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT11_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT11_TXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt11_drpaddr_in,
        drpclk_in                       =>      gt11_drpclk_in,
        drpdi_in                        =>      gt11_drpdi_in,
        drpdo_out                       =>      gt11_drpdo_out,
        drpen_in                        =>      gt11_drpen_in,
        drprdy_out                      =>      gt11_drprdy_out,
        drpwe_in                        =>      gt11_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt11_qpllclk_i,
        qpllrefclk_in                   =>      gt11_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt11_eyescanreset_in,
        rxuserrdy_in                    =>      gt11_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt11_eyescandataerror_out,
        eyescantrigger_in               =>      gt11_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt11_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt11_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt11_rxusrclk_in,
        rxusrclk2_in                    =>      gt11_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt11_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt11_rxdisperr_out,
        rxnotintable_out                =>      gt11_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt11_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt11_rxdlyen_in,
        rxdlysreset_in                  =>      gt11_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt11_rxdlysresetdone_out,
        rxphalign_in                    =>      gt11_rxphalign_in,
        rxphaligndone_out               =>      gt11_rxphaligndone_out,
        rxphalignen_in                  =>      gt11_rxphalignen_in,
        rxphdlyreset_in                 =>      gt11_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt11_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt11_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt11_rxsyncallin_in,
        rxsyncdone_out                  =>      gt11_rxsyncdone_out,
        rxsyncin_in                     =>      gt11_rxsyncin_in,
        rxsyncmode_in                   =>      gt11_rxsyncmode_in,
        rxsyncout_out                   =>      gt11_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt11_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt11_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt11_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt11_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt11_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt11_rxoutclk_out,
        rxoutclkfabric_out              =>      gt11_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt11_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt11_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt11_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt11_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt11_gttxreset_in,
        txuserrdy_in                    =>      gt11_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt11_txusrclk_in,
        txusrclk2_in                    =>      gt11_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt11_txdlyen_in,
        txdlysreset_in                  =>      gt11_txdlysreset_in,
        txdlysresetdone_out             =>      gt11_txdlysresetdone_out,
        txphalign_in                    =>      gt11_txphalign_in,
        txphaligndone_out               =>      gt11_txphaligndone_out,
        txphalignen_in                  =>      gt11_txphalignen_in,
        txphdlyreset_in                 =>      gt11_txphdlyreset_in,
        txphinit_in                     =>      gt11_txphinit_in,
        txphinitdone_out                =>      gt11_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt11_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt11_gthtxn_out,
        gthtxp_out                      =>      gt11_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt11_txoutclk_out,
        txoutclkfabric_out              =>      gt11_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt11_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt11_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt11_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT12  (X0Y16)
gt12_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_OVRD_IN         => ('1'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt12_rst_i,
        DRP_BUSY_OUT                    =>      GT12_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT12_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT12_TXPMARESETDONE_OUT,
        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt12_drpaddr_in,
        drpclk_in                       =>      gt12_drpclk_in,
        drpdi_in                        =>      gt12_drpdi_in,
        drpdo_out                       =>      gt12_drpdo_out,
        drpen_in                        =>      gt12_drpen_in,
        drprdy_out                      =>      gt12_drprdy_out,
        drpwe_in                        =>      gt12_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt12_qpllclk_i,
        qpllrefclk_in                   =>      gt12_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt12_eyescanreset_in,
        rxuserrdy_in                    =>      gt12_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt12_eyescandataerror_out,
        eyescantrigger_in               =>      gt12_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt12_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt12_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt12_rxusrclk_in,
        rxusrclk2_in                    =>      gt12_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt12_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt12_rxdisperr_out,
        rxnotintable_out                =>      gt12_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt12_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt12_rxdlyen_in,
        rxdlysreset_in                  =>      gt12_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt12_rxdlysresetdone_out,
        rxphalign_in                    =>      gt12_rxphalign_in,
        rxphaligndone_out               =>      gt12_rxphaligndone_out,
        rxphalignen_in                  =>      gt12_rxphalignen_in,
        rxphdlyreset_in                 =>      gt12_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt12_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt12_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt12_rxsyncallin_in,
        rxsyncdone_out                  =>      gt12_rxsyncdone_out,
        rxsyncin_in                     =>      gt12_rxsyncin_in,
        rxsyncmode_in                   =>      gt12_rxsyncmode_in,
        rxsyncout_out                   =>      gt12_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt12_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt12_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt12_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt12_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt12_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt12_rxoutclk_out,
        rxoutclkfabric_out              =>      gt12_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt12_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt12_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt12_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt12_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt12_gttxreset_in,
        txuserrdy_in                    =>      gt12_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt12_txusrclk_in,
        txusrclk2_in                    =>      gt12_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt12_txdlyen_in,
        txdlysreset_in                  =>      gt12_txdlysreset_in,
        txdlysresetdone_out             =>      gt12_txdlysresetdone_out,
        txphalign_in                    =>      gt12_txphalign_in,
        txphaligndone_out               =>      gt12_txphaligndone_out,
        txphalignen_in                  =>      gt12_txphalignen_in,
        txphdlyreset_in                 =>      gt12_txphdlyreset_in,
        txphinit_in                     =>      gt12_txphinit_in,
        txphinitdone_out                =>      gt12_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt12_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt12_gthtxn_out,
        gthtxp_out                      =>      gt12_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt12_txoutclk_out,
        txoutclkfabric_out              =>      gt12_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt12_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt12_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt12_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT13  (X0Y17)
gt13_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt13_rst_i,
        DRP_BUSY_OUT                    =>      GT13_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT13_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT13_TXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt13_drpaddr_in,
        drpclk_in                       =>      gt13_drpclk_in,
        drpdi_in                        =>      gt13_drpdi_in,
        drpdo_out                       =>      gt13_drpdo_out,
        drpen_in                        =>      gt13_drpen_in,
        drprdy_out                      =>      gt13_drprdy_out,
        drpwe_in                        =>      gt13_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt13_qpllclk_i,
        qpllrefclk_in                   =>      gt13_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt13_eyescanreset_in,
        rxuserrdy_in                    =>      gt13_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt13_eyescandataerror_out,
        eyescantrigger_in               =>      gt13_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt13_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt13_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt13_rxusrclk_in,
        rxusrclk2_in                    =>      gt13_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt13_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt13_rxdisperr_out,
        rxnotintable_out                =>      gt13_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt13_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt13_rxdlyen_in,
        rxdlysreset_in                  =>      gt13_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt13_rxdlysresetdone_out,
        rxphalign_in                    =>      gt13_rxphalign_in,
        rxphaligndone_out               =>      gt13_rxphaligndone_out,
        rxphalignen_in                  =>      gt13_rxphalignen_in,
        rxphdlyreset_in                 =>      gt13_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt13_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt13_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt13_rxsyncallin_in,
        rxsyncdone_out                  =>      gt13_rxsyncdone_out,
        rxsyncin_in                     =>      gt13_rxsyncin_in,
        rxsyncmode_in                   =>      gt13_rxsyncmode_in,
        rxsyncout_out                   =>      gt13_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt13_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt13_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt13_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt13_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt13_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt13_rxoutclk_out,
        rxoutclkfabric_out              =>      gt13_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt13_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt13_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt13_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt13_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt13_gttxreset_in,
        txuserrdy_in                    =>      gt13_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt13_txusrclk_in,
        txusrclk2_in                    =>      gt13_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt13_txdlyen_in,
        txdlysreset_in                  =>      gt13_txdlysreset_in,
        txdlysresetdone_out             =>      gt13_txdlysresetdone_out,
        txphalign_in                    =>      gt13_txphalign_in,
        txphaligndone_out               =>      gt13_txphaligndone_out,
        txphalignen_in                  =>      gt13_txphalignen_in,
        txphdlyreset_in                 =>      gt13_txphdlyreset_in,
        txphinit_in                     =>      gt13_txphinit_in,
        txphinitdone_out                =>      gt13_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt13_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt13_gthtxn_out,
        gthtxp_out                      =>      gt13_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt13_txoutclk_out,
        txoutclkfabric_out              =>      gt13_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt13_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt13_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt13_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT14  (X0Y18)
gt14_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt14_rst_i,
        DRP_BUSY_OUT                    =>      GT14_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT14_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT14_TXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt14_drpaddr_in,
        drpclk_in                       =>      gt14_drpclk_in,
        drpdi_in                        =>      gt14_drpdi_in,
        drpdo_out                       =>      gt14_drpdo_out,
        drpen_in                        =>      gt14_drpen_in,
        drprdy_out                      =>      gt14_drprdy_out,
        drpwe_in                        =>      gt14_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt14_qpllclk_i,
        qpllrefclk_in                   =>      gt14_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt14_eyescanreset_in,
        rxuserrdy_in                    =>      gt14_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt14_eyescandataerror_out,
        eyescantrigger_in               =>      gt14_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt14_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt14_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt14_rxusrclk_in,
        rxusrclk2_in                    =>      gt14_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt14_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt14_rxdisperr_out,
        rxnotintable_out                =>      gt14_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt14_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt14_rxdlyen_in,
        rxdlysreset_in                  =>      gt14_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt14_rxdlysresetdone_out,
        rxphalign_in                    =>      gt14_rxphalign_in,
        rxphaligndone_out               =>      gt14_rxphaligndone_out,
        rxphalignen_in                  =>      gt14_rxphalignen_in,
        rxphdlyreset_in                 =>      gt14_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt14_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt14_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt14_rxsyncallin_in,
        rxsyncdone_out                  =>      gt14_rxsyncdone_out,
        rxsyncin_in                     =>      gt14_rxsyncin_in,
        rxsyncmode_in                   =>      gt14_rxsyncmode_in,
        rxsyncout_out                   =>      gt14_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt14_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt14_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt14_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt14_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt14_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt14_rxoutclk_out,
        rxoutclkfabric_out              =>      gt14_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt14_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt14_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt14_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt14_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt14_gttxreset_in,
        txuserrdy_in                    =>      gt14_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt14_txusrclk_in,
        txusrclk2_in                    =>      gt14_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt14_txdlyen_in,
        txdlysreset_in                  =>      gt14_txdlysreset_in,
        txdlysresetdone_out             =>      gt14_txdlysresetdone_out,
        txphalign_in                    =>      gt14_txphalign_in,
        txphaligndone_out               =>      gt14_txphaligndone_out,
        txphalignen_in                  =>      gt14_txphalignen_in,
        txphdlyreset_in                 =>      gt14_txphdlyreset_in,
        txphinit_in                     =>      gt14_txphinit_in,
        txphinitdone_out                =>      gt14_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt14_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt14_gthtxn_out,
        gthtxp_out                      =>      gt14_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt14_txoutclk_out,
        txoutclkfabric_out              =>      gt14_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt14_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt14_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt14_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT15  (X0Y19)
gt15_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt15_rst_i,
        DRP_BUSY_OUT                    =>      GT15_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT15_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT15_TXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt15_drpaddr_in,
        drpclk_in                       =>      gt15_drpclk_in,
        drpdi_in                        =>      gt15_drpdi_in,
        drpdo_out                       =>      gt15_drpdo_out,
        drpen_in                        =>      gt15_drpen_in,
        drprdy_out                      =>      gt15_drprdy_out,
        drpwe_in                        =>      gt15_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt15_qpllclk_i,
        qpllrefclk_in                   =>      gt15_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt15_eyescanreset_in,
        rxuserrdy_in                    =>      gt15_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt15_eyescandataerror_out,
        eyescantrigger_in               =>      gt15_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt15_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt15_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt15_rxusrclk_in,
        rxusrclk2_in                    =>      gt15_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt15_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt15_rxdisperr_out,
        rxnotintable_out                =>      gt15_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt15_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt15_rxdlyen_in,
        rxdlysreset_in                  =>      gt15_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt15_rxdlysresetdone_out,
        rxphalign_in                    =>      gt15_rxphalign_in,
        rxphaligndone_out               =>      gt15_rxphaligndone_out,
        rxphalignen_in                  =>      gt15_rxphalignen_in,
        rxphdlyreset_in                 =>      gt15_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt15_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt15_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt15_rxsyncallin_in,
        rxsyncdone_out                  =>      gt15_rxsyncdone_out,
        rxsyncin_in                     =>      gt15_rxsyncin_in,
        rxsyncmode_in                   =>      gt15_rxsyncmode_in,
        rxsyncout_out                   =>      gt15_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt15_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt15_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt15_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt15_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt15_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt15_rxoutclk_out,
        rxoutclkfabric_out              =>      gt15_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt15_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt15_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt15_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt15_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt15_gttxreset_in,
        txuserrdy_in                    =>      gt15_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt15_txusrclk_in,
        txusrclk2_in                    =>      gt15_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt15_txdlyen_in,
        txdlysreset_in                  =>      gt15_txdlysreset_in,
        txdlysresetdone_out             =>      gt15_txdlysresetdone_out,
        txphalign_in                    =>      gt15_txphalign_in,
        txphaligndone_out               =>      gt15_txphaligndone_out,
        txphalignen_in                  =>      gt15_txphalignen_in,
        txphdlyreset_in                 =>      gt15_txphdlyreset_in,
        txphinit_in                     =>      gt15_txphinit_in,
        txphinitdone_out                =>      gt15_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt15_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt15_gthtxn_out,
        gthtxp_out                      =>      gt15_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt15_txoutclk_out,
        txoutclkfabric_out              =>      gt15_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt15_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt15_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt15_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT16  (X0Y20)
gt16_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt16_rst_i,
        DRP_BUSY_OUT                    =>      GT16_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT16_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT16_TXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt16_drpaddr_in,
        drpclk_in                       =>      gt16_drpclk_in,
        drpdi_in                        =>      gt16_drpdi_in,
        drpdo_out                       =>      gt16_drpdo_out,
        drpen_in                        =>      gt16_drpen_in,
        drprdy_out                      =>      gt16_drprdy_out,
        drpwe_in                        =>      gt16_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt16_qpllclk_i,
        qpllrefclk_in                   =>      gt16_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt16_eyescanreset_in,
        rxuserrdy_in                    =>      gt16_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt16_eyescandataerror_out,
        eyescantrigger_in               =>      gt16_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt16_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt16_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt16_rxusrclk_in,
        rxusrclk2_in                    =>      gt16_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt16_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt16_rxdisperr_out,
        rxnotintable_out                =>      gt16_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt16_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt16_rxdlyen_in,
        rxdlysreset_in                  =>      gt16_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt16_rxdlysresetdone_out,
        rxphalign_in                    =>      gt16_rxphalign_in,
        rxphaligndone_out               =>      gt16_rxphaligndone_out,
        rxphalignen_in                  =>      gt16_rxphalignen_in,
        rxphdlyreset_in                 =>      gt16_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt16_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt16_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt16_rxsyncallin_in,
        rxsyncdone_out                  =>      gt16_rxsyncdone_out,
        rxsyncin_in                     =>      gt16_rxsyncin_in,
        rxsyncmode_in                   =>      gt16_rxsyncmode_in,
        rxsyncout_out                   =>      gt16_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt16_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt16_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt16_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt16_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt16_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt16_rxoutclk_out,
        rxoutclkfabric_out              =>      gt16_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt16_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt16_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt16_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt16_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt16_gttxreset_in,
        txuserrdy_in                    =>      gt16_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt16_txusrclk_in,
        txusrclk2_in                    =>      gt16_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt16_txdlyen_in,
        txdlysreset_in                  =>      gt16_txdlysreset_in,
        txdlysresetdone_out             =>      gt16_txdlysresetdone_out,
        txphalign_in                    =>      gt16_txphalign_in,
        txphaligndone_out               =>      gt16_txphaligndone_out,
        txphalignen_in                  =>      gt16_txphalignen_in,
        txphdlyreset_in                 =>      gt16_txphdlyreset_in,
        txphinit_in                     =>      gt16_txphinit_in,
        txphinitdone_out                =>      gt16_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt16_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt16_gthtxn_out,
        gthtxp_out                      =>      gt16_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt16_txoutclk_out,
        txoutclkfabric_out              =>      gt16_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt16_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt16_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt16_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT17  (X0Y21)
gt17_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt17_rst_i,
        DRP_BUSY_OUT                    =>      GT17_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT17_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT17_TXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt17_drpaddr_in,
        drpclk_in                       =>      gt17_drpclk_in,
        drpdi_in                        =>      gt17_drpdi_in,
        drpdo_out                       =>      gt17_drpdo_out,
        drpen_in                        =>      gt17_drpen_in,
        drprdy_out                      =>      gt17_drprdy_out,
        drpwe_in                        =>      gt17_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt17_qpllclk_i,
        qpllrefclk_in                   =>      gt17_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt17_eyescanreset_in,
        rxuserrdy_in                    =>      gt17_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt17_eyescandataerror_out,
        eyescantrigger_in               =>      gt17_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt17_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt17_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt17_rxusrclk_in,
        rxusrclk2_in                    =>      gt17_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt17_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt17_rxdisperr_out,
        rxnotintable_out                =>      gt17_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt17_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt17_rxdlyen_in,
        rxdlysreset_in                  =>      gt17_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt17_rxdlysresetdone_out,
        rxphalign_in                    =>      gt17_rxphalign_in,
        rxphaligndone_out               =>      gt17_rxphaligndone_out,
        rxphalignen_in                  =>      gt17_rxphalignen_in,
        rxphdlyreset_in                 =>      gt17_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt17_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt17_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt17_rxsyncallin_in,
        rxsyncdone_out                  =>      gt17_rxsyncdone_out,
        rxsyncin_in                     =>      gt17_rxsyncin_in,
        rxsyncmode_in                   =>      gt17_rxsyncmode_in,
        rxsyncout_out                   =>      gt17_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt17_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt17_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt17_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt17_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt17_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt17_rxoutclk_out,
        rxoutclkfabric_out              =>      gt17_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt17_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt17_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt17_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt17_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt17_gttxreset_in,
        txuserrdy_in                    =>      gt17_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt17_txusrclk_in,
        txusrclk2_in                    =>      gt17_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt17_txdlyen_in,
        txdlysreset_in                  =>      gt17_txdlysreset_in,
        txdlysresetdone_out             =>      gt17_txdlysresetdone_out,
        txphalign_in                    =>      gt17_txphalign_in,
        txphaligndone_out               =>      gt17_txphaligndone_out,
        txphalignen_in                  =>      gt17_txphalignen_in,
        txphdlyreset_in                 =>      gt17_txphdlyreset_in,
        txphinit_in                     =>      gt17_txphinit_in,
        txphinitdone_out                =>      gt17_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt17_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt17_gthtxn_out,
        gthtxp_out                      =>      gt17_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt17_txoutclk_out,
        txoutclkfabric_out              =>      gt17_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt17_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt17_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt17_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT18  (X0Y22)
gt18_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt18_rst_i,
        DRP_BUSY_OUT                    =>      GT18_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT18_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT18_TXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt18_drpaddr_in,
        drpclk_in                       =>      gt18_drpclk_in,
        drpdi_in                        =>      gt18_drpdi_in,
        drpdo_out                       =>      gt18_drpdo_out,
        drpen_in                        =>      gt18_drpen_in,
        drprdy_out                      =>      gt18_drprdy_out,
        drpwe_in                        =>      gt18_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt18_qpllclk_i,
        qpllrefclk_in                   =>      gt18_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt18_eyescanreset_in,
        rxuserrdy_in                    =>      gt18_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt18_eyescandataerror_out,
        eyescantrigger_in               =>      gt18_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt18_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt18_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt18_rxusrclk_in,
        rxusrclk2_in                    =>      gt18_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt18_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt18_rxdisperr_out,
        rxnotintable_out                =>      gt18_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt18_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt18_rxdlyen_in,
        rxdlysreset_in                  =>      gt18_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt18_rxdlysresetdone_out,
        rxphalign_in                    =>      gt18_rxphalign_in,
        rxphaligndone_out               =>      gt18_rxphaligndone_out,
        rxphalignen_in                  =>      gt18_rxphalignen_in,
        rxphdlyreset_in                 =>      gt18_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt18_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt18_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt18_rxsyncallin_in,
        rxsyncdone_out                  =>      gt18_rxsyncdone_out,
        rxsyncin_in                     =>      gt18_rxsyncin_in,
        rxsyncmode_in                   =>      gt18_rxsyncmode_in,
        rxsyncout_out                   =>      gt18_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt18_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt18_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt18_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt18_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt18_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt18_rxoutclk_out,
        rxoutclkfabric_out              =>      gt18_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt18_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt18_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt18_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt18_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt18_gttxreset_in,
        txuserrdy_in                    =>      gt18_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt18_txusrclk_in,
        txusrclk2_in                    =>      gt18_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt18_txdlyen_in,
        txdlysreset_in                  =>      gt18_txdlysreset_in,
        txdlysresetdone_out             =>      gt18_txdlysresetdone_out,
        txphalign_in                    =>      gt18_txphalign_in,
        txphaligndone_out               =>      gt18_txphaligndone_out,
        txphalignen_in                  =>      gt18_txphalignen_in,
        txphdlyreset_in                 =>      gt18_txphdlyreset_in,
        txphinit_in                     =>      gt18_txphinit_in,
        txphinitdone_out                =>      gt18_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt18_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt18_gthtxn_out,
        gthtxp_out                      =>      gt18_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt18_txoutclk_out,
        txoutclkfabric_out              =>      gt18_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt18_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt18_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt18_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT19  (X0Y23)
gt19_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt19_rst_i,
        DRP_BUSY_OUT                    =>      GT19_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT19_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT19_TXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt19_drpaddr_in,
        drpclk_in                       =>      gt19_drpclk_in,
        drpdi_in                        =>      gt19_drpdi_in,
        drpdo_out                       =>      gt19_drpdo_out,
        drpen_in                        =>      gt19_drpen_in,
        drprdy_out                      =>      gt19_drprdy_out,
        drpwe_in                        =>      gt19_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt19_qpllclk_i,
        qpllrefclk_in                   =>      gt19_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt19_eyescanreset_in,
        rxuserrdy_in                    =>      gt19_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt19_eyescandataerror_out,
        eyescantrigger_in               =>      gt19_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt19_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt19_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt19_rxusrclk_in,
        rxusrclk2_in                    =>      gt19_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt19_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt19_rxdisperr_out,
        rxnotintable_out                =>      gt19_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt19_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt19_rxdlyen_in,
        rxdlysreset_in                  =>      gt19_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt19_rxdlysresetdone_out,
        rxphalign_in                    =>      gt19_rxphalign_in,
        rxphaligndone_out               =>      gt19_rxphaligndone_out,
        rxphalignen_in                  =>      gt19_rxphalignen_in,
        rxphdlyreset_in                 =>      gt19_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt19_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt19_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt19_rxsyncallin_in,
        rxsyncdone_out                  =>      gt19_rxsyncdone_out,
        rxsyncin_in                     =>      gt19_rxsyncin_in,
        rxsyncmode_in                   =>      gt19_rxsyncmode_in,
        rxsyncout_out                   =>      gt19_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt19_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt19_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt19_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt19_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt19_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt19_rxoutclk_out,
        rxoutclkfabric_out              =>      gt19_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt19_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt19_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt19_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt19_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt19_gttxreset_in,
        txuserrdy_in                    =>      gt19_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt19_txusrclk_in,
        txusrclk2_in                    =>      gt19_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt19_txdlyen_in,
        txdlysreset_in                  =>      gt19_txdlysreset_in,
        txdlysresetdone_out             =>      gt19_txdlysresetdone_out,
        txphalign_in                    =>      gt19_txphalign_in,
        txphaligndone_out               =>      gt19_txphaligndone_out,
        txphalignen_in                  =>      gt19_txphalignen_in,
        txphdlyreset_in                 =>      gt19_txphdlyreset_in,
        txphinit_in                     =>      gt19_txphinit_in,
        txphinitdone_out                =>      gt19_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt19_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt19_gthtxn_out,
        gthtxp_out                      =>      gt19_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt19_txoutclk_out,
        txoutclkfabric_out              =>      gt19_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt19_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt19_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt19_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT20  (X0Y24)
gt20_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt20_rst_i,
        DRP_BUSY_OUT                    =>      GT20_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT20_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT20_TXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt20_drpaddr_in,
        drpclk_in                       =>      gt20_drpclk_in,
        drpdi_in                        =>      gt20_drpdi_in,
        drpdo_out                       =>      gt20_drpdo_out,
        drpen_in                        =>      gt20_drpen_in,
        drprdy_out                      =>      gt20_drprdy_out,
        drpwe_in                        =>      gt20_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt20_qpllclk_i,
        qpllrefclk_in                   =>      gt20_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt20_eyescanreset_in,
        rxuserrdy_in                    =>      gt20_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt20_eyescandataerror_out,
        eyescantrigger_in               =>      gt20_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt20_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt20_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt20_rxusrclk_in,
        rxusrclk2_in                    =>      gt20_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt20_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt20_rxdisperr_out,
        rxnotintable_out                =>      gt20_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt20_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt20_rxdlyen_in,
        rxdlysreset_in                  =>      gt20_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt20_rxdlysresetdone_out,
        rxphalign_in                    =>      gt20_rxphalign_in,
        rxphaligndone_out               =>      gt20_rxphaligndone_out,
        rxphalignen_in                  =>      gt20_rxphalignen_in,
        rxphdlyreset_in                 =>      gt20_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt20_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt20_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt20_rxsyncallin_in,
        rxsyncdone_out                  =>      gt20_rxsyncdone_out,
        rxsyncin_in                     =>      gt20_rxsyncin_in,
        rxsyncmode_in                   =>      gt20_rxsyncmode_in,
        rxsyncout_out                   =>      gt20_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt20_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt20_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt20_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt20_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt20_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt20_rxoutclk_out,
        rxoutclkfabric_out              =>      gt20_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt20_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt20_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt20_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt20_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt20_gttxreset_in,
        txuserrdy_in                    =>      gt20_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt20_txusrclk_in,
        txusrclk2_in                    =>      gt20_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt20_txdlyen_in,
        txdlysreset_in                  =>      gt20_txdlysreset_in,
        txdlysresetdone_out             =>      gt20_txdlysresetdone_out,
        txphalign_in                    =>      gt20_txphalign_in,
        txphaligndone_out               =>      gt20_txphaligndone_out,
        txphalignen_in                  =>      gt20_txphalignen_in,
        txphdlyreset_in                 =>      gt20_txphdlyreset_in,
        txphinit_in                     =>      gt20_txphinit_in,
        txphinitdone_out                =>      gt20_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt20_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt20_gthtxn_out,
        gthtxp_out                      =>      gt20_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt20_txoutclk_out,
        txoutclkfabric_out              =>      gt20_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt20_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt20_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt20_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT21  (X0Y25)
gt21_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt21_rst_i,
        DRP_BUSY_OUT                    =>      GT21_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT21_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT21_TXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt21_drpaddr_in,
        drpclk_in                       =>      gt21_drpclk_in,
        drpdi_in                        =>      gt21_drpdi_in,
        drpdo_out                       =>      gt21_drpdo_out,
        drpen_in                        =>      gt21_drpen_in,
        drprdy_out                      =>      gt21_drprdy_out,
        drpwe_in                        =>      gt21_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt21_qpllclk_i,
        qpllrefclk_in                   =>      gt21_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt21_eyescanreset_in,
        rxuserrdy_in                    =>      gt21_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt21_eyescandataerror_out,
        eyescantrigger_in               =>      gt21_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt21_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt21_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt21_rxusrclk_in,
        rxusrclk2_in                    =>      gt21_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt21_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt21_rxdisperr_out,
        rxnotintable_out                =>      gt21_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt21_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt21_rxdlyen_in,
        rxdlysreset_in                  =>      gt21_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt21_rxdlysresetdone_out,
        rxphalign_in                    =>      gt21_rxphalign_in,
        rxphaligndone_out               =>      gt21_rxphaligndone_out,
        rxphalignen_in                  =>      gt21_rxphalignen_in,
        rxphdlyreset_in                 =>      gt21_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt21_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt21_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt21_rxsyncallin_in,
        rxsyncdone_out                  =>      gt21_rxsyncdone_out,
        rxsyncin_in                     =>      gt21_rxsyncin_in,
        rxsyncmode_in                   =>      gt21_rxsyncmode_in,
        rxsyncout_out                   =>      gt21_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt21_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt21_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt21_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt21_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt21_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt21_rxoutclk_out,
        rxoutclkfabric_out              =>      gt21_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt21_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt21_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt21_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt21_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt21_gttxreset_in,
        txuserrdy_in                    =>      gt21_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt21_txusrclk_in,
        txusrclk2_in                    =>      gt21_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt21_txdlyen_in,
        txdlysreset_in                  =>      gt21_txdlysreset_in,
        txdlysresetdone_out             =>      gt21_txdlysresetdone_out,
        txphalign_in                    =>      gt21_txphalign_in,
        txphaligndone_out               =>      gt21_txphaligndone_out,
        txphalignen_in                  =>      gt21_txphalignen_in,
        txphdlyreset_in                 =>      gt21_txphdlyreset_in,
        txphinit_in                     =>      gt21_txphinit_in,
        txphinitdone_out                =>      gt21_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt21_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt21_gthtxn_out,
        gthtxp_out                      =>      gt21_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt21_txoutclk_out,
        txoutclkfabric_out              =>      gt21_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt21_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt21_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt21_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT22  (X0Y26)
gt22_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt22_rst_i,
        DRP_BUSY_OUT                    =>      GT22_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT22_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT22_TXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt22_drpaddr_in,
        drpclk_in                       =>      gt22_drpclk_in,
        drpdi_in                        =>      gt22_drpdi_in,
        drpdo_out                       =>      gt22_drpdo_out,
        drpen_in                        =>      gt22_drpen_in,
        drprdy_out                      =>      gt22_drprdy_out,
        drpwe_in                        =>      gt22_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt22_qpllclk_i,
        qpllrefclk_in                   =>      gt22_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt22_eyescanreset_in,
        rxuserrdy_in                    =>      gt22_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt22_eyescandataerror_out,
        eyescantrigger_in               =>      gt22_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt22_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt22_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt22_rxusrclk_in,
        rxusrclk2_in                    =>      gt22_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt22_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt22_rxdisperr_out,
        rxnotintable_out                =>      gt22_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt22_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt22_rxdlyen_in,
        rxdlysreset_in                  =>      gt22_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt22_rxdlysresetdone_out,
        rxphalign_in                    =>      gt22_rxphalign_in,
        rxphaligndone_out               =>      gt22_rxphaligndone_out,
        rxphalignen_in                  =>      gt22_rxphalignen_in,
        rxphdlyreset_in                 =>      gt22_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt22_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt22_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt22_rxsyncallin_in,
        rxsyncdone_out                  =>      gt22_rxsyncdone_out,
        rxsyncin_in                     =>      gt22_rxsyncin_in,
        rxsyncmode_in                   =>      gt22_rxsyncmode_in,
        rxsyncout_out                   =>      gt22_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt22_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt22_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt22_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt22_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt22_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt22_rxoutclk_out,
        rxoutclkfabric_out              =>      gt22_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt22_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt22_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt22_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt22_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt22_gttxreset_in,
        txuserrdy_in                    =>      gt22_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt22_txusrclk_in,
        txusrclk2_in                    =>      gt22_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt22_txdlyen_in,
        txdlysreset_in                  =>      gt22_txdlysreset_in,
        txdlysresetdone_out             =>      gt22_txdlysresetdone_out,
        txphalign_in                    =>      gt22_txphalign_in,
        txphaligndone_out               =>      gt22_txphaligndone_out,
        txphalignen_in                  =>      gt22_txphalignen_in,
        txphdlyreset_in                 =>      gt22_txphdlyreset_in,
        txphinit_in                     =>      gt22_txphinit_in,
        txphinitdone_out                =>      gt22_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt22_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt22_gthtxn_out,
        gthtxp_out                      =>      gt22_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt22_txoutclk_out,
        txoutclkfabric_out              =>      gt22_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt22_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt22_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt22_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT23  (X0Y27)
gt23_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt23_rst_i,
        DRP_BUSY_OUT                    =>      GT23_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT23_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT23_TXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt23_drpaddr_in,
        drpclk_in                       =>      gt23_drpclk_in,
        drpdi_in                        =>      gt23_drpdi_in,
        drpdo_out                       =>      gt23_drpdo_out,
        drpen_in                        =>      gt23_drpen_in,
        drprdy_out                      =>      gt23_drprdy_out,
        drpwe_in                        =>      gt23_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt23_qpllclk_i,
        qpllrefclk_in                   =>      gt23_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt23_eyescanreset_in,
        rxuserrdy_in                    =>      gt23_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt23_eyescandataerror_out,
        eyescantrigger_in               =>      gt23_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt23_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt23_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt23_rxusrclk_in,
        rxusrclk2_in                    =>      gt23_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt23_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt23_rxdisperr_out,
        rxnotintable_out                =>      gt23_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt23_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt23_rxdlyen_in,
        rxdlysreset_in                  =>      gt23_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt23_rxdlysresetdone_out,
        rxphalign_in                    =>      gt23_rxphalign_in,
        rxphaligndone_out               =>      gt23_rxphaligndone_out,
        rxphalignen_in                  =>      gt23_rxphalignen_in,
        rxphdlyreset_in                 =>      gt23_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt23_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt23_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt23_rxsyncallin_in,
        rxsyncdone_out                  =>      gt23_rxsyncdone_out,
        rxsyncin_in                     =>      gt23_rxsyncin_in,
        rxsyncmode_in                   =>      gt23_rxsyncmode_in,
        rxsyncout_out                   =>      gt23_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt23_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt23_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt23_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt23_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt23_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt23_rxoutclk_out,
        rxoutclkfabric_out              =>      gt23_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt23_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt23_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt23_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt23_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt23_gttxreset_in,
        txuserrdy_in                    =>      gt23_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt23_txusrclk_in,
        txusrclk2_in                    =>      gt23_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt23_txdlyen_in,
        txdlysreset_in                  =>      gt23_txdlysreset_in,
        txdlysresetdone_out             =>      gt23_txdlysresetdone_out,
        txphalign_in                    =>      gt23_txphalign_in,
        txphaligndone_out               =>      gt23_txphaligndone_out,
        txphalignen_in                  =>      gt23_txphalignen_in,
        txphdlyreset_in                 =>      gt23_txphdlyreset_in,
        txphinit_in                     =>      gt23_txphinit_in,
        txphinitdone_out                =>      gt23_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt23_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt23_gthtxn_out,
        gthtxp_out                      =>      gt23_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt23_txoutclk_out,
        txoutclkfabric_out              =>      gt23_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt23_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt23_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt23_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT24  (X0Y28)
gt24_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_OVRD_IN         => ('1'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt24_rst_i,
        DRP_BUSY_OUT                    =>      GT24_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT24_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT24_TXPMARESETDONE_OUT,
        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt24_drpaddr_in,
        drpclk_in                       =>      gt24_drpclk_in,
        drpdi_in                        =>      gt24_drpdi_in,
        drpdo_out                       =>      gt24_drpdo_out,
        drpen_in                        =>      gt24_drpen_in,
        drprdy_out                      =>      gt24_drprdy_out,
        drpwe_in                        =>      gt24_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt24_qpllclk_i,
        qpllrefclk_in                   =>      gt24_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt24_eyescanreset_in,
        rxuserrdy_in                    =>      gt24_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt24_eyescandataerror_out,
        eyescantrigger_in               =>      gt24_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt24_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt24_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt24_rxusrclk_in,
        rxusrclk2_in                    =>      gt24_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt24_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt24_rxdisperr_out,
        rxnotintable_out                =>      gt24_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt24_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt24_rxdlyen_in,
        rxdlysreset_in                  =>      gt24_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt24_rxdlysresetdone_out,
        rxphalign_in                    =>      gt24_rxphalign_in,
        rxphaligndone_out               =>      gt24_rxphaligndone_out,
        rxphalignen_in                  =>      gt24_rxphalignen_in,
        rxphdlyreset_in                 =>      gt24_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt24_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt24_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt24_rxsyncallin_in,
        rxsyncdone_out                  =>      gt24_rxsyncdone_out,
        rxsyncin_in                     =>      gt24_rxsyncin_in,
        rxsyncmode_in                   =>      gt24_rxsyncmode_in,
        rxsyncout_out                   =>      gt24_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt24_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt24_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt24_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt24_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt24_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt24_rxoutclk_out,
        rxoutclkfabric_out              =>      gt24_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt24_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt24_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt24_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt24_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt24_gttxreset_in,
        txuserrdy_in                    =>      gt24_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt24_txusrclk_in,
        txusrclk2_in                    =>      gt24_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt24_txdlyen_in,
        txdlysreset_in                  =>      gt24_txdlysreset_in,
        txdlysresetdone_out             =>      gt24_txdlysresetdone_out,
        txphalign_in                    =>      gt24_txphalign_in,
        txphaligndone_out               =>      gt24_txphaligndone_out,
        txphalignen_in                  =>      gt24_txphalignen_in,
        txphdlyreset_in                 =>      gt24_txphdlyreset_in,
        txphinit_in                     =>      gt24_txphinit_in,
        txphinitdone_out                =>      gt24_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt24_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt24_gthtxn_out,
        gthtxp_out                      =>      gt24_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt24_txoutclk_out,
        txoutclkfabric_out              =>      gt24_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt24_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt24_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt24_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT25  (X0Y29)
gt25_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt25_rst_i,
        DRP_BUSY_OUT                    =>      GT25_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT25_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT25_TXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt25_drpaddr_in,
        drpclk_in                       =>      gt25_drpclk_in,
        drpdi_in                        =>      gt25_drpdi_in,
        drpdo_out                       =>      gt25_drpdo_out,
        drpen_in                        =>      gt25_drpen_in,
        drprdy_out                      =>      gt25_drprdy_out,
        drpwe_in                        =>      gt25_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt25_qpllclk_i,
        qpllrefclk_in                   =>      gt25_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt25_eyescanreset_in,
        rxuserrdy_in                    =>      gt25_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt25_eyescandataerror_out,
        eyescantrigger_in               =>      gt25_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt25_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt25_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt25_rxusrclk_in,
        rxusrclk2_in                    =>      gt25_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt25_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt25_rxdisperr_out,
        rxnotintable_out                =>      gt25_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt25_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt25_rxdlyen_in,
        rxdlysreset_in                  =>      gt25_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt25_rxdlysresetdone_out,
        rxphalign_in                    =>      gt25_rxphalign_in,
        rxphaligndone_out               =>      gt25_rxphaligndone_out,
        rxphalignen_in                  =>      gt25_rxphalignen_in,
        rxphdlyreset_in                 =>      gt25_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt25_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt25_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt25_rxsyncallin_in,
        rxsyncdone_out                  =>      gt25_rxsyncdone_out,
        rxsyncin_in                     =>      gt25_rxsyncin_in,
        rxsyncmode_in                   =>      gt25_rxsyncmode_in,
        rxsyncout_out                   =>      gt25_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt25_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt25_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt25_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt25_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt25_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt25_rxoutclk_out,
        rxoutclkfabric_out              =>      gt25_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt25_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt25_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt25_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt25_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt25_gttxreset_in,
        txuserrdy_in                    =>      gt25_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt25_txusrclk_in,
        txusrclk2_in                    =>      gt25_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt25_txdlyen_in,
        txdlysreset_in                  =>      gt25_txdlysreset_in,
        txdlysresetdone_out             =>      gt25_txdlysresetdone_out,
        txphalign_in                    =>      gt25_txphalign_in,
        txphaligndone_out               =>      gt25_txphaligndone_out,
        txphalignen_in                  =>      gt25_txphalignen_in,
        txphdlyreset_in                 =>      gt25_txphdlyreset_in,
        txphinit_in                     =>      gt25_txphinit_in,
        txphinitdone_out                =>      gt25_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt25_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt25_gthtxn_out,
        gthtxp_out                      =>      gt25_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt25_txoutclk_out,
        txoutclkfabric_out              =>      gt25_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt25_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt25_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt25_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT26  (X0Y30)
gt26_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt26_rst_i,
        DRP_BUSY_OUT                    =>      GT26_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT26_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT26_TXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt26_drpaddr_in,
        drpclk_in                       =>      gt26_drpclk_in,
        drpdi_in                        =>      gt26_drpdi_in,
        drpdo_out                       =>      gt26_drpdo_out,
        drpen_in                        =>      gt26_drpen_in,
        drprdy_out                      =>      gt26_drprdy_out,
        drpwe_in                        =>      gt26_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt26_qpllclk_i,
        qpllrefclk_in                   =>      gt26_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt26_eyescanreset_in,
        rxuserrdy_in                    =>      gt26_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt26_eyescandataerror_out,
        eyescantrigger_in               =>      gt26_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt26_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt26_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt26_rxusrclk_in,
        rxusrclk2_in                    =>      gt26_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt26_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt26_rxdisperr_out,
        rxnotintable_out                =>      gt26_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt26_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt26_rxdlyen_in,
        rxdlysreset_in                  =>      gt26_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt26_rxdlysresetdone_out,
        rxphalign_in                    =>      gt26_rxphalign_in,
        rxphaligndone_out               =>      gt26_rxphaligndone_out,
        rxphalignen_in                  =>      gt26_rxphalignen_in,
        rxphdlyreset_in                 =>      gt26_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt26_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt26_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt26_rxsyncallin_in,
        rxsyncdone_out                  =>      gt26_rxsyncdone_out,
        rxsyncin_in                     =>      gt26_rxsyncin_in,
        rxsyncmode_in                   =>      gt26_rxsyncmode_in,
        rxsyncout_out                   =>      gt26_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt26_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt26_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt26_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt26_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt26_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt26_rxoutclk_out,
        rxoutclkfabric_out              =>      gt26_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt26_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt26_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt26_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt26_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt26_gttxreset_in,
        txuserrdy_in                    =>      gt26_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt26_txusrclk_in,
        txusrclk2_in                    =>      gt26_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt26_txdlyen_in,
        txdlysreset_in                  =>      gt26_txdlysreset_in,
        txdlysresetdone_out             =>      gt26_txdlysresetdone_out,
        txphalign_in                    =>      gt26_txphalign_in,
        txphaligndone_out               =>      gt26_txphaligndone_out,
        txphalignen_in                  =>      gt26_txphalignen_in,
        txphdlyreset_in                 =>      gt26_txphdlyreset_in,
        txphinit_in                     =>      gt26_txphinit_in,
        txphinitdone_out                =>      gt26_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt26_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt26_gthtxn_out,
        gthtxp_out                      =>      gt26_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt26_txoutclk_out,
        txoutclkfabric_out              =>      gt26_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt26_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt26_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt26_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT27  (X0Y31)
gt27_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt27_rst_i,
        DRP_BUSY_OUT                    =>      GT27_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT27_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT27_TXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt27_drpaddr_in,
        drpclk_in                       =>      gt27_drpclk_in,
        drpdi_in                        =>      gt27_drpdi_in,
        drpdo_out                       =>      gt27_drpdo_out,
        drpen_in                        =>      gt27_drpen_in,
        drprdy_out                      =>      gt27_drprdy_out,
        drpwe_in                        =>      gt27_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt27_qpllclk_i,
        qpllrefclk_in                   =>      gt27_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt27_eyescanreset_in,
        rxuserrdy_in                    =>      gt27_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt27_eyescandataerror_out,
        eyescantrigger_in               =>      gt27_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt27_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt27_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt27_rxusrclk_in,
        rxusrclk2_in                    =>      gt27_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt27_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt27_rxdisperr_out,
        rxnotintable_out                =>      gt27_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt27_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt27_rxdlyen_in,
        rxdlysreset_in                  =>      gt27_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt27_rxdlysresetdone_out,
        rxphalign_in                    =>      gt27_rxphalign_in,
        rxphaligndone_out               =>      gt27_rxphaligndone_out,
        rxphalignen_in                  =>      gt27_rxphalignen_in,
        rxphdlyreset_in                 =>      gt27_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt27_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt27_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt27_rxsyncallin_in,
        rxsyncdone_out                  =>      gt27_rxsyncdone_out,
        rxsyncin_in                     =>      gt27_rxsyncin_in,
        rxsyncmode_in                   =>      gt27_rxsyncmode_in,
        rxsyncout_out                   =>      gt27_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt27_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt27_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt27_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt27_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt27_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt27_rxoutclk_out,
        rxoutclkfabric_out              =>      gt27_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt27_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt27_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt27_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt27_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt27_gttxreset_in,
        txuserrdy_in                    =>      gt27_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt27_txusrclk_in,
        txusrclk2_in                    =>      gt27_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt27_txdlyen_in,
        txdlysreset_in                  =>      gt27_txdlysreset_in,
        txdlysresetdone_out             =>      gt27_txdlysresetdone_out,
        txphalign_in                    =>      gt27_txphalign_in,
        txphaligndone_out               =>      gt27_txphaligndone_out,
        txphalignen_in                  =>      gt27_txphalignen_in,
        txphdlyreset_in                 =>      gt27_txphdlyreset_in,
        txphinit_in                     =>      gt27_txphinit_in,
        txphinitdone_out                =>      gt27_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt27_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt27_gthtxn_out,
        gthtxp_out                      =>      gt27_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt27_txoutclk_out,
        txoutclkfabric_out              =>      gt27_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt27_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt27_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt27_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT28  (X0Y32)
gt28_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt28_rst_i,
        DRP_BUSY_OUT                    =>      GT28_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT28_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT28_TXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt28_drpaddr_in,
        drpclk_in                       =>      gt28_drpclk_in,
        drpdi_in                        =>      gt28_drpdi_in,
        drpdo_out                       =>      gt28_drpdo_out,
        drpen_in                        =>      gt28_drpen_in,
        drprdy_out                      =>      gt28_drprdy_out,
        drpwe_in                        =>      gt28_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt28_qpllclk_i,
        qpllrefclk_in                   =>      gt28_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt28_eyescanreset_in,
        rxuserrdy_in                    =>      gt28_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt28_eyescandataerror_out,
        eyescantrigger_in               =>      gt28_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt28_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt28_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt28_rxusrclk_in,
        rxusrclk2_in                    =>      gt28_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt28_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt28_rxdisperr_out,
        rxnotintable_out                =>      gt28_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt28_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt28_rxdlyen_in,
        rxdlysreset_in                  =>      gt28_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt28_rxdlysresetdone_out,
        rxphalign_in                    =>      gt28_rxphalign_in,
        rxphaligndone_out               =>      gt28_rxphaligndone_out,
        rxphalignen_in                  =>      gt28_rxphalignen_in,
        rxphdlyreset_in                 =>      gt28_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt28_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt28_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt28_rxsyncallin_in,
        rxsyncdone_out                  =>      gt28_rxsyncdone_out,
        rxsyncin_in                     =>      gt28_rxsyncin_in,
        rxsyncmode_in                   =>      gt28_rxsyncmode_in,
        rxsyncout_out                   =>      gt28_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt28_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt28_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt28_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt28_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt28_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt28_rxoutclk_out,
        rxoutclkfabric_out              =>      gt28_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt28_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt28_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt28_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt28_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt28_gttxreset_in,
        txuserrdy_in                    =>      gt28_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt28_txusrclk_in,
        txusrclk2_in                    =>      gt28_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt28_txdlyen_in,
        txdlysreset_in                  =>      gt28_txdlysreset_in,
        txdlysresetdone_out             =>      gt28_txdlysresetdone_out,
        txphalign_in                    =>      gt28_txphalign_in,
        txphaligndone_out               =>      gt28_txphaligndone_out,
        txphalignen_in                  =>      gt28_txphalignen_in,
        txphdlyreset_in                 =>      gt28_txphdlyreset_in,
        txphinit_in                     =>      gt28_txphinit_in,
        txphinitdone_out                =>      gt28_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt28_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt28_gthtxn_out,
        gthtxp_out                      =>      gt28_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt28_txoutclk_out,
        txoutclkfabric_out              =>      gt28_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt28_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt28_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt28_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT29  (X0Y33)
gt29_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt29_rst_i,
        DRP_BUSY_OUT                    =>      GT29_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT29_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT29_TXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt29_drpaddr_in,
        drpclk_in                       =>      gt29_drpclk_in,
        drpdi_in                        =>      gt29_drpdi_in,
        drpdo_out                       =>      gt29_drpdo_out,
        drpen_in                        =>      gt29_drpen_in,
        drprdy_out                      =>      gt29_drprdy_out,
        drpwe_in                        =>      gt29_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt29_qpllclk_i,
        qpllrefclk_in                   =>      gt29_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt29_eyescanreset_in,
        rxuserrdy_in                    =>      gt29_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt29_eyescandataerror_out,
        eyescantrigger_in               =>      gt29_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt29_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt29_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt29_rxusrclk_in,
        rxusrclk2_in                    =>      gt29_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt29_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt29_rxdisperr_out,
        rxnotintable_out                =>      gt29_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt29_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt29_rxdlyen_in,
        rxdlysreset_in                  =>      gt29_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt29_rxdlysresetdone_out,
        rxphalign_in                    =>      gt29_rxphalign_in,
        rxphaligndone_out               =>      gt29_rxphaligndone_out,
        rxphalignen_in                  =>      gt29_rxphalignen_in,
        rxphdlyreset_in                 =>      gt29_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt29_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt29_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt29_rxsyncallin_in,
        rxsyncdone_out                  =>      gt29_rxsyncdone_out,
        rxsyncin_in                     =>      gt29_rxsyncin_in,
        rxsyncmode_in                   =>      gt29_rxsyncmode_in,
        rxsyncout_out                   =>      gt29_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt29_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt29_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt29_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt29_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt29_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt29_rxoutclk_out,
        rxoutclkfabric_out              =>      gt29_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt29_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt29_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt29_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt29_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt29_gttxreset_in,
        txuserrdy_in                    =>      gt29_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt29_txusrclk_in,
        txusrclk2_in                    =>      gt29_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt29_txdlyen_in,
        txdlysreset_in                  =>      gt29_txdlysreset_in,
        txdlysresetdone_out             =>      gt29_txdlysresetdone_out,
        txphalign_in                    =>      gt29_txphalign_in,
        txphaligndone_out               =>      gt29_txphaligndone_out,
        txphalignen_in                  =>      gt29_txphalignen_in,
        txphdlyreset_in                 =>      gt29_txphdlyreset_in,
        txphinit_in                     =>      gt29_txphinit_in,
        txphinitdone_out                =>      gt29_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt29_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt29_gthtxn_out,
        gthtxp_out                      =>      gt29_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt29_txoutclk_out,
        txoutclkfabric_out              =>      gt29_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt29_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt29_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt29_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT30  (X0Y34)
gt30_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt30_rst_i,
        DRP_BUSY_OUT                    =>      GT30_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT30_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT30_TXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt30_drpaddr_in,
        drpclk_in                       =>      gt30_drpclk_in,
        drpdi_in                        =>      gt30_drpdi_in,
        drpdo_out                       =>      gt30_drpdo_out,
        drpen_in                        =>      gt30_drpen_in,
        drprdy_out                      =>      gt30_drprdy_out,
        drpwe_in                        =>      gt30_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt30_qpllclk_i,
        qpllrefclk_in                   =>      gt30_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt30_eyescanreset_in,
        rxuserrdy_in                    =>      gt30_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt30_eyescandataerror_out,
        eyescantrigger_in               =>      gt30_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt30_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt30_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt30_rxusrclk_in,
        rxusrclk2_in                    =>      gt30_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt30_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt30_rxdisperr_out,
        rxnotintable_out                =>      gt30_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt30_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt30_rxdlyen_in,
        rxdlysreset_in                  =>      gt30_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt30_rxdlysresetdone_out,
        rxphalign_in                    =>      gt30_rxphalign_in,
        rxphaligndone_out               =>      gt30_rxphaligndone_out,
        rxphalignen_in                  =>      gt30_rxphalignen_in,
        rxphdlyreset_in                 =>      gt30_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt30_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt30_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt30_rxsyncallin_in,
        rxsyncdone_out                  =>      gt30_rxsyncdone_out,
        rxsyncin_in                     =>      gt30_rxsyncin_in,
        rxsyncmode_in                   =>      gt30_rxsyncmode_in,
        rxsyncout_out                   =>      gt30_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt30_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt30_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt30_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt30_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt30_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt30_rxoutclk_out,
        rxoutclkfabric_out              =>      gt30_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt30_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt30_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt30_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt30_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt30_gttxreset_in,
        txuserrdy_in                    =>      gt30_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt30_txusrclk_in,
        txusrclk2_in                    =>      gt30_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt30_txdlyen_in,
        txdlysreset_in                  =>      gt30_txdlysreset_in,
        txdlysresetdone_out             =>      gt30_txdlysresetdone_out,
        txphalign_in                    =>      gt30_txphalign_in,
        txphaligndone_out               =>      gt30_txphaligndone_out,
        txphalignen_in                  =>      gt30_txphalignen_in,
        txphdlyreset_in                 =>      gt30_txphdlyreset_in,
        txphinit_in                     =>      gt30_txphinit_in,
        txphinitdone_out                =>      gt30_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt30_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt30_gthtxn_out,
        gthtxp_out                      =>      gt30_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt30_txoutclk_out,
        txoutclkfabric_out              =>      gt30_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt30_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt30_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt30_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT31  (X0Y35)
gt31_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        SIM_CPLLREFCLK_SEL     =>  "001",
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt31_rst_i,
        DRP_BUSY_OUT                    =>      GT31_DRP_BUSY_OUT,
        RXPMARESETDONE                  =>      GT31_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT31_TXPMARESETDONE_OUT,

        cpllrefclksel_in => "001",
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt31_drpaddr_in,
        drpclk_in                       =>      gt31_drpclk_in,
        drpdi_in                        =>      gt31_drpdi_in,
        drpdo_out                       =>      gt31_drpdo_out,
        drpen_in                        =>      gt31_drpen_in,
        drprdy_out                      =>      gt31_drprdy_out,
        drpwe_in                        =>      gt31_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt31_qpllclk_i,
        qpllrefclk_in                   =>      gt31_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt31_eyescanreset_in,
        rxuserrdy_in                    =>      gt31_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt31_eyescandataerror_out,
        eyescantrigger_in               =>      gt31_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        rxslide_in                      =>      gt31_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt31_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt31_rxusrclk_in,
        rxusrclk2_in                    =>      gt31_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt31_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt31_rxdisperr_out,
        rxnotintable_out                =>      gt31_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt31_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt31_rxdlyen_in,
        rxdlysreset_in                  =>      gt31_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt31_rxdlysresetdone_out,
        rxphalign_in                    =>      gt31_rxphalign_in,
        rxphaligndone_out               =>      gt31_rxphaligndone_out,
        rxphalignen_in                  =>      gt31_rxphalignen_in,
        rxphdlyreset_in                 =>      gt31_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt31_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt31_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt31_rxsyncallin_in,
        rxsyncdone_out                  =>      gt31_rxsyncdone_out,
        rxsyncin_in                     =>      gt31_rxsyncin_in,
        rxsyncmode_in                   =>      gt31_rxsyncmode_in,
        rxsyncout_out                   =>      gt31_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt31_rxbyteisaligned_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt31_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt31_rxlpmlfhold_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxmonitorout_out                =>      gt31_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt31_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt31_rxoutclk_out,
        rxoutclkfabric_out              =>      gt31_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt31_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt31_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt31_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt31_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt31_gttxreset_in,
        txuserrdy_in                    =>      gt31_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt31_txusrclk_in,
        txusrclk2_in                    =>      gt31_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt31_txdlyen_in,
        txdlysreset_in                  =>      gt31_txdlysreset_in,
        txdlysresetdone_out             =>      gt31_txdlysresetdone_out,
        txphalign_in                    =>      gt31_txphalign_in,
        txphaligndone_out               =>      gt31_txphaligndone_out,
        txphalignen_in                  =>      gt31_txphalignen_in,
        txphdlyreset_in                 =>      gt31_txphdlyreset_in,
        txphinit_in                     =>      gt31_txphinit_in,
        txphinitdone_out                =>      gt31_txphinitdone_out,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt31_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt31_gthtxn_out,
        gthtxp_out                      =>      gt31_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt31_txoutclk_out,
        txoutclkfabric_out              =>      gt31_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt31_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt31_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt31_txcharisk_in

    );
    

end RTL;
     
