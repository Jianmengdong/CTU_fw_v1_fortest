
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
library UNISIM;
use UNISIM.VComponents.all;

package CTU_pack is

    type t_array8 is array (integer range<>) of std_logic_vector(7 downto 0);
    type t_array16 is array (integer range<>) of std_logic_vector(15 downto 0);
    type t_array48 is array (integer range<>) of std_logic_vector(47 downto 0);
    type t_array64 is array (integer range<>) of std_logic_vector(63 downto 0);
    type t_array672 is array (integer range<>) of std_logic_vector(671 downto 0);
    
    type t_uarray16 is array (integer range<>) of unsigned(15 downto 0);
    constant VFL_NUMBER : integer range 1 to 180 := 110;
    --constant delay_cycle_vector : t_array672(VFL_NUMBER - 1 downto 0) := 
        --(0=> x"888887777777777766666666666666665555555555555555555555554444444444444444444444444444444333333333533333333333333333333222222222222222222221111111111111111111000000000000"
        --1=> x"888877777777777666666666666666655555555555555555555555544444444444444444444444444444443333333335333333333333333333332222222222222222222211111111111111111110000000000008",
        --2=> x"888777777777776666666666666666555555555555555555555555444444444444444444444444444444433333333353333333333333333333322222222222222222222111111111111111111100000000000088",
        --3=> x"887777777777766666666666666665555555555555555555555554444444444444444444444444444444333333333533333333333333333333222222222222222222221111111111111111111000000000000888",
        --4=> x"877777777777666666666666666655555555555555555555555544444444444444444444444444444443333333335333333333333333333332222222222222222222211111111111111111110000000000008888",
        --5=> x"777777777776666666666666666555555555555555555555555444444444444444444444444444444433333333353333333333333333333322222222222222222222111111111111111111100000000000088888",
        --6=> x"777777777766666666666666665555555555555555555555554444444444444444444444444444444333333333533333333333333333333222222222222222222221111111111111111111000000000000888887",
        --7=> x"777777777666666666666666655555555555555555555555544444444444444444444444444444443333333335333333333333333333332222222222222222222211111111111111111110000000000008888877",
        --8=> x"777777776666666666666666555555555555555555555555444444444444444444444444444444433333333353333333333333333333322222222222222222222111111111111111111100000000000088888777",
        --9=> x"777777766666666666666665555555555555555555555554444444444444444444444444444444333333333533333333333333333333222222222222222222221111111111111111111000000000000888887777",
        --10=> x"777777666666666666666655555555555555555555555544444444444444444444444444444443333333335333333333333333333332222222222222222222211111111111111111110000000000008888877777",
        --11=> x"777777666666666666666655555555555555555555555544444444444444444444444444444443333333335333333333333333333332222222222222222222211111111111111111110000000000008888877777",
        --12=> x"777776666666666666666555555555555555555555555444444444444444444444444444444433333333353333333333333333333322222222222222222222111111111111111111100000000000088888777777",
        --13=> x"777766666666666666665555555555555555555555554444444444444444444444444444444333333333533333333333333333333222222222222222222221111111111111111111000000000000888887777777",
        --14=> x"777666666666666666655555555555555555555555544444444444444444444444444444443333333335333333333333333333332222222222222222222211111111111111111110000000000008888877777777",
        --15=> x"776666666666666666555555555555555555555555444444444444444444444444444444433333333353333333333333333333322222222222222222222111111111111111111100000000000088888777777777",
        --16=> x"766666666666666665555555555555555555555554444444444444444444444444444444333333333533333333333333333333222222222222222222221111111111111111111000000000000888887777777777",
        --17=> x"666666666666666655555555555555555555555544444444444444444444444444444443333333335333333333333333333332222222222222222222211111111111111111110000000000008888877777777777",
        --18=> x"666666666666666555555555555555555555555444444444444444444444444444444433333333353333333333333333333322222222222222222222111111111111111111100000000000088888777777777776",
        --19=> x"666666666666665555555555555555555555554444444444444444444444444444444333333333533333333333333333333222222222222222222221111111111111111111000000000000888887777777777766",
        --20=> x"666666666666655555555555555555555555544444444444444444444444444444443333333335333333333333333333332222222222222222222211111111111111111110000000000008888877777777777666",
        --21=> x"666666666666555555555555555555555555444444444444444444444444444444433333333353333333333333333333322222222222222222222111111111111111111100000000000088888777777777776666",
        --22=> x"666666666665555555555555555555555554444444444444444444444444444444333333333533333333333333333333222222222222222222221111111111111111111000000000000888887777777777766666",
        --23=> x"666666666655555555555555555555555544444444444444444444444444444443333333335333333333333333333332222222222222222222211111111111111111110000000000008888877777777777666666",
        --24=> x"666666666555555555555555555555555444444444444444444444444444444433333333353333333333333333333322222222222222222222111111111111111111100000000000088888777777777776666666",
        --25=> x"666666665555555555555555555555554444444444444444444444444444444333333333533333333333333333333222222222222222222221111111111111111111000000000000888887777777777766666666",
        --26=> x"666666655555555555555555555555544444444444444444444444444444443333333335333333333333333333332222222222222222222211111111111111111110000000000008888877777777777666666666",
        --27=> x"666666555555555555555555555555444444444444444444444444444444433333333353333333333333333333322222222222222222222111111111111111111100000000000088888777777777776666666666",
        --28=> x"666665555555555555555555555554444444444444444444444444444444333333333533333333333333333333222222222222222222221111111111111111111000000000000888887777777777766666666666",
        --29=> x"666655555555555555555555555544444444444444444444444444444443333333335333333333333333333332222222222222222222211111111111111111110000000000008888877777777777666666666666",
        --30=> x"666555555555555555555555555444444444444444444444444444444433333333353333333333333333333322222222222222222222111111111111111111100000000000088888777777777776666666666666",
        --31=> x"665555555555555555555555554444444444444444444444444444444333333333533333333333333333333222222222222222222221111111111111111111000000000000888887777777777766666666666666",
        --32=> x"655555555555555555555555544444444444444444444444444444443333333335333333333333333333332222222222222222222211111111111111111110000000000008888877777777777666666666666666",
        --33=> x"555555555555555555555555444444444444444444444444444444433333333353333333333333333333322222222222222222222111111111111111111100000000000088888777777777776666666666666666",
        --34=> x"555555555555555555555554444444444444444444444444444444333333333533333333333333333333222222222222222222221111111111111111111000000000000888887777777777766666666666666665",
        --35=> x"555555555555555555555544444444444444444444444444444443333333335333333333333333333332222222222222222222211111111111111111110000000000008888877777777777666666666666666655",
        --36=> x"555555555555555555555444444444444444444444444444444433333333353333333333333333333322222222222222222222111111111111111111100000000000088888777777777776666666666666666555",
        --37=> x"555555555555555555554444444444444444444444444444444333333333533333333333333333333222222222222222222221111111111111111111000000000000888887777777777766666666666666665555",
        --38=> x"555555555555555555544444444444444444444444444444443333333335333333333333333333332222222222222222222211111111111111111110000000000008888877777777777666666666666666655555",
        --39=> x"555555555555555555444444444444444444444444444444433333333353333333333333333333322222222222222222222111111111111111111100000000000088888777777777776666666666666666555555",
        --40=> x"555555555555555554444444444444444444444444444444333333333533333333333333333333222222222222222222221111111111111111111000000000000888887777777777766666666666666665555555",
        --41=> x"555555555555555544444444444444444444444444444443333333335333333333333333333332222222222222222222211111111111111111110000000000008888877777777777666666666666666655555555",
        --42=> x"555555555555555444444444444444444444444444444433333333353333333333333333333322222222222222222222111111111111111111100000000000088888777777777776666666666666666555555555",
        --43=> x"555555555555554444444444444444444444444444444333333333533333333333333333333222222222222222222221111111111111111111000000000000888887777777777766666666666666665555555555",
        --44=> x"555555555555544444444444444444444444444444443333333335333333333333333333332222222222222222222211111111111111111110000000000008888877777777777666666666666666655555555555",
        --45=> x"555555555555444444444444444444444444444444433333333353333333333333333333322222222222222222222111111111111111111100000000000088888777777777776666666666666666555555555555",
        --46=> x"555555555554444444444444444444444444444444333333333533333333333333333333222222222222222222221111111111111111111000000000000888887777777777766666666666666665555555555555",
        --47=> x"555555555544444444444444444444444444444443333333335333333333333333333332222222222222222222211111111111111111110000000000008888877777777777666666666666666655555555555555",
        --48=> x"555555555444444444444444444444444444444433333333353333333333333333333322222222222222222222111111111111111111100000000000088888777777777776666666666666666555555555555555",
        --49=> x"555555554444444444444444444444444444444333333333533333333333333333333222222222222222222221111111111111111111000000000000888887777777777766666666666666665555555555555555",
        --50=> x"555555544444444444444444444444444444443333333335333333333333333333332222222222222222222211111111111111111110000000000008888877777777777666666666666666655555555555555555",
        --51=> x"555555544444444444444444444444444444443333333335333333333333333333332222222222222222222211111111111111111110000000000008888877777777777666666666666666655555555555555555",
        --52=> x"555555444444444444444444444444444444433333333353333333333333333333322222222222222222222111111111111111111100000000000088888777777777776666666666666666555555555555555555",
        --53=> x"555554444444444444444444444444444444333333333533333333333333333333222222222222222222221111111111111111111000000000000888887777777777766666666666666665555555555555555555",
        --54=> x"555544444444444444444444444444444443333333335333333333333333333332222222222222222222211111111111111111110000000000008888877777777777666666666666666655555555555555555555",
        --55=> x"555444444444444444444444444444444433333333353333333333333333333322222222222222222222111111111111111111100000000000088888777777777776666666666666666555555555555555555555",
        --56=> x"554444444444444444444444444444444333333333533333333333333333333222222222222222222221111111111111111111000000000000888887777777777766666666666666665555555555555555555555",
        --57=> x"544444444444444444444444444444443333333335333333333333333333332222222222222222222211111111111111111110000000000008888877777777777666666666666666655555555555555555555555",
        --58=> x"444444444444444444444444444444433333333353333333333333333333322222222222222222222111111111111111111100000000000088888777777777776666666666666666555555555555555555555555",
        --59=> x"444444444444444444444444444444333333333533333333333333333333222222222222222222221111111111111111111000000000000888887777777777766666666666666665555555555555555555555554",
        --60=> x"444444444444444444444444444443333333335333333333333333333332222222222222222222211111111111111111110000000000008888877777777777666666666666666655555555555555555555555544",
        --61=> x"444444444444444444444444444433333333353333333333333333333322222222222222222222111111111111111111100000000000088888777777777776666666666666666555555555555555555555555444",
        --62=> x"444444444444444444444444444333333333533333333333333333333222222222222222222221111111111111111111000000000000888887777777777766666666666666665555555555555555555555554444",
        --63=> x"444444444444444444444444443333333335333333333333333333332222222222222222222211111111111111111110000000000008888877777777777666666666666666655555555555555555555555544444",
        --64=> x"444444444444444444444444433333333353333333333333333333322222222222222222222111111111111111111100000000000088888777777777776666666666666666555555555555555555555555444444",
        --65=> x"444444444444444444444444333333333533333333333333333333222222222222222222221111111111111111111000000000000888887777777777766666666666666665555555555555555555555554444444",
        --66=> x"444444444444444444444443333333335333333333333333333332222222222222222222211111111111111111110000000000008888877777777777666666666666666655555555555555555555555544444444",
        --67=> x"444444444444444444444433333333353333333333333333333322222222222222222222111111111111111111100000000000088888777777777776666666666666666555555555555555555555555444444444",
        --68=> x"444444444444444444444333333333533333333333333333333222222222222222222221111111111111111111000000000000888887777777777766666666666666665555555555555555555555554444444444",
        --69=> x"444444444444444444443333333335333333333333333333332222222222222222222211111111111111111110000000000008888877777777777666666666666666655555555555555555555555544444444444",
        --70=> x"444444444444444444433333333353333333333333333333322222222222222222222111111111111111111100000000000088888777777777776666666666666666555555555555555555555555444444444444",
        --71=> x"444444444444444444333333333533333333333333333333222222222222222222221111111111111111111000000000000888887777777777766666666666666665555555555555555555555554444444444444",
        --72=> x"444444444444444443333333335333333333333333333332222222222222222222211111111111111111110000000000008888877777777777666666666666666655555555555555555555555544444444444444",
        --73=> x"444444444444444433333333353333333333333333333322222222222222222222111111111111111111100000000000088888777777777776666666666666666555555555555555555555555444444444444444",
        --74=> x"444444444444444333333333533333333333333333333222222222222222222221111111111111111111000000000000888887777777777766666666666666665555555555555555555555554444444444444444",
        --75=> x"444444444444443333333335333333333333333333332222222222222222222211111111111111111110000000000008888877777777777666666666666666655555555555555555555555544444444444444444",
        --76=> x"444444444444433333333353333333333333333333322222222222222222222111111111111111111100000000000088888777777777776666666666666666555555555555555555555555444444444444444444",
        --77=> x"444444444444333333333533333333333333333333222222222222222222221111111111111111111000000000000888887777777777766666666666666665555555555555555555555554444444444444444444",
        --78=> x"444444444443333333335333333333333333333332222222222222222222211111111111111111110000000000008888877777777777666666666666666655555555555555555555555544444444444444444444",
        --79=> x"444444444433333333353333333333333333333322222222222222222222111111111111111111100000000000088888777777777776666666666666666555555555555555555555555444444444444444444444",
        --80=> x"444444444333333333533333333333333333333222222222222222222221111111111111111111000000000000888887777777777766666666666666665555555555555555555555554444444444444444444444",
        --81=> x"444444443333333335333333333333333333332222222222222222222211111111111111111110000000000008888877777777777666666666666666655555555555555555555555544444444444444444444444",
        --82=> x"444444433333333353333333333333333333322222222222222222222111111111111111111100000000000088888777777777776666666666666666555555555555555555555555444444444444444444444444",
        --83=> x"444444333333333533333333333333333333222222222222222222221111111111111111111000000000000888887777777777766666666666666665555555555555555555555554444444444444444444444444",
        --84=> x"444443333333335333333333333333333332222222222222222222211111111111111111110000000000008888877777777777666666666666666655555555555555555555555544444444444444444444444444",
        --85=> x"444433333333353333333333333333333322222222222222222222111111111111111111100000000000088888777777777776666666666666666555555555555555555555555444444444444444444444444444",
        --86=> x"444333333333533333333333333333333222222222222222222221111111111111111111000000000000888887777777777766666666666666665555555555555555555555554444444444444444444444444444",
        --87=> x"443333333335333333333333333333332222222222222222222211111111111111111110000000000008888877777777777666666666666666655555555555555555555555544444444444444444444444444444",
        --88=> x"433333333353333333333333333333322222222222222222222111111111111111111100000000000088888777777777776666666666666666555555555555555555555555444444444444444444444444444444",
        --89=> x"333333333533333333333333333333222222222222222222221111111111111111111000000000000888887777777777766666666666666665555555555555555555555554444444444444444444444444444444",
        --90=> x"333333335333333333333333333332222222222222222222211111111111111111110000000000008888877777777777666666666666666655555555555555555555555544444444444444444444444444444443",
        --91=> x"333333335333333333333333333332222222222222222222211111111111111111110000000000008888877777777777666666666666666655555555555555555555555544444444444444444444444444444443",
        --92=> x"333333353333333333333333333322222222222222222222111111111111111111100000000000088888777777777776666666666666666555555555555555555555555444444444444444444444444444444433",
        --93=> x"333333533333333333333333333222222222222222222221111111111111111111000000000000888887777777777766666666666666665555555555555555555555554444444444444444444444444444444333",
        --94=> x"333335333333333333333333332222222222222222222211111111111111111110000000000008888877777777777666666666666666655555555555555555555555544444444444444444444444444444443333",
        --95=> x"333353333333333333333333322222222222222222222111111111111111111100000000000088888777777777776666666666666666555555555555555555555555444444444444444444444444444444433333",
        --96=> x"333533333333333333333333222222222222222222221111111111111111111000000000000888887777777777766666666666666665555555555555555555555554444444444444444444444444444444333333",
        --97=> x"335333333333333333333332222222222222222222211111111111111111110000000000008888877777777777666666666666666655555555555555555555555544444444444444444444444444444443333333",
        --98=> x"353333333333333333333322222222222222222222111111111111111111100000000000088888777777777776666666666666666555555555555555555555555444444444444444444444444444444433333333",
        --99=> x"533333333333333333333222222222222222222221111111111111111111000000000000888887777777777766666666666666665555555555555555555555554444444444444444444444444444444333333333",
        --100=> x"333333333333333333332222222222222222222211111111111111111110000000000008888877777777777666666666666666655555555555555555555555544444444444444444444444444444443333333335",
        --101=> x"333333333333333333322222222222222222222111111111111111111100000000000088888777777777776666666666666666555555555555555555555555444444444444444444444444444444433333333353",
        --102=> x"333333333333333333222222222222222222221111111111111111111000000000000888887777777777766666666666666665555555555555555555555554444444444444444444444444444444333333333533",
        --103=> x"333333333333333332222222222222222222211111111111111111110000000000008888877777777777666666666666666655555555555555555555555544444444444444444444444444444443333333335333",
        --104=> x"333333333333333322222222222222222222111111111111111111100000000000088888777777777776666666666666666555555555555555555555555444444444444444444444444444444433333333353333",
        --105=> x"333333333333333222222222222222222221111111111111111111000000000000888887777777777766666666666666665555555555555555555555554444444444444444444444444444444333333333533333",
        --106=> x"333333333333332222222222222222222211111111111111111110000000000008888877777777777666666666666666655555555555555555555555544444444444444444444444444444443333333335333333",
        --107=> x"333333333333322222222222222222222111111111111111111100000000000088888777777777776666666666666666555555555555555555555555444444444444444444444444444444433333333353333333",
        --108=> x"333333333333222222222222222222221111111111111111111000000000000888887777777777766666666666666665555555555555555555555554444444444444444444444444444444333333333533333333",
        --109=> x"333333333332222222222222222222211111111111111111110000000000008888877777777777666666666666666655555555555555555555555544444444444444444444444444444443333333335333333333",
        --110=> x"333333333322222222222222222222111111111111111111100000000000088888777777777776666666666666666555555555555555555555555444444444444444444444444444444433333333353333333333",
        --111=> x"333333333222222222222222222221111111111111111111000000000000888887777777777766666666666666665555555555555555555555554444444444444444444444444444444333333333533333333333",
        --112=> x"333333332222222222222222222211111111111111111110000000000008888877777777777666666666666666655555555555555555555555544444444444444444444444444444443333333335333333333333",
        --113=> x"333333322222222222222222222111111111111111111100000000000088888777777777776666666666666666555555555555555555555555444444444444444444444444444444433333333353333333333333",
        --114=> x"333333222222222222222222221111111111111111111000000000000888887777777777766666666666666665555555555555555555555554444444444444444444444444444444333333333533333333333333",
        --115=> x"333332222222222222222222211111111111111111110000000000008888877777777777666666666666666655555555555555555555555544444444444444444444444444444443333333335333333333333333",
        --116=> x"333322222222222222222222111111111111111111100000000000088888777777777776666666666666666555555555555555555555555444444444444444444444444444444433333333353333333333333333",
        --117=> x"333222222222222222222221111111111111111111000000000000888887777777777766666666666666665555555555555555555555554444444444444444444444444444444333333333533333333333333333",
        --118=> x"332222222222222222222211111111111111111110000000000008888877777777777666666666666666655555555555555555555555544444444444444444444444444444443333333335333333333333333333",
        --119=> x"322222222222222222222111111111111111111100000000000088888777777777776666666666666666555555555555555555555555444444444444444444444444444444433333333353333333333333333333",
        --120=> x"222222222222111111111111111111100000000000088888777777777776666666666666666555555555555555555555555444444444444444444444444444444433333333353333333333333333333322222222",
        --121=> x"222222222221111111111111111111000000000000888887777777777766666666666666665555555555555555555555554444444444444444444444444444444333333333533333333333333333333222222222",
        --122=> x"222222222211111111111111111110000000000008888877777777777666666666666666655555555555555555555555544444444444444444444444444444443333333335333333333333333333332222222222",
        --123=> x"222222222111111111111111111100000000000088888777777777776666666666666666555555555555555555555555444444444444444444444444444444433333333353333333333333333333322222222222",
        --124=> x"222222221111111111111111111000000000000888887777777777766666666666666665555555555555555555555554444444444444444444444444444444333333333533333333333333333333222222222222",
        --125=> x"222222211111111111111111110000000000008888877777777777666666666666666655555555555555555555555544444444444444444444444444444443333333335333333333333333333332222222222222",
        --126=> x"222222111111111111111111100000000000088888777777777776666666666666666555555555555555555555555444444444444444444444444444444433333333353333333333333333333322222222222222",
        --127=> x"222221111111111111111111000000000000888887777777777766666666666666665555555555555555555555554444444444444444444444444444444333333333533333333333333333333222222222222222",
        --128=> x"222211111111111111111110000000000008888877777777777666666666666666655555555555555555555555544444444444444444444444444444443333333335333333333333333333332222222222222222",
        --129=> x"222111111111111111111100000000000088888777777777776666666666666666555555555555555555555555444444444444444444444444444444433333333353333333333333333333322222222222222222",
        --130=> x"221111111111111111111000000000000888887777777777766666666666666665555555555555555555555554444444444444444444444444444444333333333533333333333333333333222222222222222222",
        --131=> x"211111111111111111110000000000008888877777777777666666666666666655555555555555555555555544444444444444444444444444444443333333335333333333333333333332222222222222222222",
        --132=> x"111111111111111111100000000000088888777777777776666666666666666555555555555555555555555444444444444444444444444444444433333333353333333333333333333322222222222222222222",
        --133=> x"111111111111111111000000000000888887777777777766666666666666665555555555555555555555554444444444444444444444444444444333333333533333333333333333333222222222222222222221",
        --134=> x"111111111111111110000000000008888877777777777666666666666666655555555555555555555555544444444444444444444444444444443333333335333333333333333333332222222222222222222211",
        --135=> x"111111111111111100000000000088888777777777776666666666666666555555555555555555555555444444444444444444444444444444433333333353333333333333333333322222222222222222222111",
        --136=> x"111111111111111000000000000888887777777777766666666666666665555555555555555555555554444444444444444444444444444444333333333533333333333333333333222222222222222222221111",
        --137=> x"111111111111110000000000008888877777777777666666666666666655555555555555555555555544444444444444444444444444444443333333335333333333333333333332222222222222222222211111",
        --138=> x"111111111111100000000000088888777777777776666666666666666555555555555555555555555444444444444444444444444444444433333333353333333333333333333322222222222222222222111111",
        --139=> x"111111111111000000000000888887777777777766666666666666665555555555555555555555554444444444444444444444444444444333333333533333333333333333333222222222222222222221111111",
        --140=> x"111111111110000000000008888877777777777666666666666666655555555555555555555555544444444444444444444444444444443333333335333333333333333333332222222222222222222211111111",
        --141=> x"111111111100000000000088888777777777776666666666666666555555555555555555555555444444444444444444444444444444433333333353333333333333333333322222222222222222222111111111",
        --142=> x"111111111000000000000888887777777777766666666666666665555555555555555555555554444444444444444444444444444444333333333533333333333333333333222222222222222222221111111111",
        --143=> x"111111110000000000008888877777777777666666666666666655555555555555555555555544444444444444444444444444444443333333335333333333333333333332222222222222222222211111111111",
        --144=> x"111111100000000000088888777777777776666666666666666555555555555555555555555444444444444444444444444444444433333333353333333333333333333322222222222222222222111111111111",
        --145=> x"111111000000000000888887777777777766666666666666665555555555555555555555554444444444444444444444444444444333333333533333333333333333333222222222222222222221111111111111",
        --146=> x"111110000000000008888877777777777666666666666666655555555555555555555555544444444444444444444444444444443333333335333333333333333333332222222222222222222211111111111111",
        --147=> x"111100000000000088888777777777776666666666666666555555555555555555555555444444444444444444444444444444433333333353333333333333333333322222222222222222222111111111111111",
        --148=> x"111000000000000888887777777777766666666666666665555555555555555555555554444444444444444444444444444444333333333533333333333333333333222222222222222222221111111111111111",
        --149=> x"110000000000008888877777777777666666666666666655555555555555555555555544444444444444444444444444444443333333335333333333333333333332222222222222222222211111111111111111",
        --150=> x"100000000000088888777777777776666666666666666555555555555555555555555444444444444444444444444444444433333333353333333333333333333322222222222222222222111111111111111111",
        --151=> x"000000000000888887777777777766666666666666665555555555555555555555554444444444444444444444444444444333333333533333333333333333333222222222222222222221111111111111111111",
        --152=> x"000000000008888877777777777666666666666666655555555555555555555555544444444444444444444444444444443333333335333333333333333333332222222222222222222211111111111111111110",
        --153=> x"000000000088888777777777776666666666666666555555555555555555555555444444444444444444444444444444433333333353333333333333333333322222222222222222222111111111111111111100",
        --154=> x"000000000888887777777777766666666666666665555555555555555555555554444444444444444444444444444444333333333533333333333333333333222222222222222222221111111111111111111000",
        --155=> x"000000008888877777777777666666666666666655555555555555555555555544444444444444444444444444444443333333335333333333333333333332222222222222222222211111111111111111110000",
        --156=> x"000000088888777777777776666666666666666555555555555555555555555444444444444444444444444444444433333333353333333333333333333322222222222222222222111111111111111111100000",
        --157=> x"000000888887777777777766666666666666665555555555555555555555554444444444444444444444444444444333333333533333333333333333333222222222222222222221111111111111111111000000",
        --158=> x"000008888877777777777666666666666666655555555555555555555555544444444444444444444444444444443333333335333333333333333333332222222222222222222211111111111111111110000000",
        --159=> x"000088888777777777776666666666666666555555555555555555555555444444444444444444444444444444433333333353333333333333333333322222222222222222222111111111111111111100000000"
        --);
    subtype t_hamming is std_logic_vector(3 downto 0);
    
    function f_hamming_encoder_4bit(data_in: std_logic_vector(3 downto 0)) return t_hamming;

end CTU_pack;

package body CTU_pack is
function f_hamming_encoder_4bit(data_in: std_logic_vector(3 downto 0)) return t_hamming is
    variable parity : std_logic_vector(3 downto 0);
    begin
        parity(3) := data_in(0) xor data_in(1) xor data_in(2);
        parity(2) := data_in(0) xor data_in(1) xor data_in(3);
        parity(1) := data_in(1) xor data_in(2) xor data_in(3);
        parity(0) := data_in(0) xor data_in(1) xor data_in(2) xor data_in(3) 
                     xor parity(1) xor parity(2) xor parity(3);
        return parity;
    end f_hamming_encoder_4bit;

end CTU_pack;
