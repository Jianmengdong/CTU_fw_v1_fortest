------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 3.6
--  \   \         Application : 7 Series FPGAs Transceivers Wizard 
--  /   /         Filename : gtwizard_0_support.vhd
-- /___/   /\      
-- \   \  /  \ 
--  \___\/\___\
--
--  Description : This module instantiates the modules required for
--                reset and initialisation of the Transceiver
--
-- Module gtwizard_0_support
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;
--***********************************Entity Declaration************************

entity gtwizard_0_support is
generic
(
    EXAMPLE_SIM_GTRESET_SPEEDUP             : string    := "TRUE";     -- simulation setting for GT SecureIP model
    STABLE_CLOCK_PERIOD                     : integer   := 8  

);
port
(
    SOFT_RESET_TX_IN                        : in   std_logic;
    SOFT_RESET_RX_IN                        : in   std_logic;
    DONT_RESET_ON_DATA_ERROR_IN             : in   std_logic;
    Q2_CLK0_GTREFCLK_PAD_N_IN               : in   std_logic;
    Q2_CLK0_GTREFCLK_PAD_P_IN               : in   std_logic;
    Q5_CLK0_GTREFCLK_PAD_N_IN               : in   std_logic;
    Q5_CLK0_GTREFCLK_PAD_P_IN               : in   std_logic;
    Q7_CLK0_GTREFCLK_PAD_N_IN               : in   std_logic;
    Q7_CLK0_GTREFCLK_PAD_P_IN               : in   std_logic;
    
    txusrclk2_in : in std_logic;
    txusrclk_in : in std_logic;

    GT0_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_DATA_VALID_IN                       : in   std_logic;
    GT0_TX_MMCM_LOCK_OUT                    : out  std_logic;
    GT0_RX_MMCM_LOCK_OUT                    : out  std_logic;
    GT1_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT1_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT1_DATA_VALID_IN                       : in   std_logic;
    GT1_TX_MMCM_LOCK_OUT                    : out  std_logic;
    GT1_RX_MMCM_LOCK_OUT                    : out  std_logic;
    GT2_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT2_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT2_DATA_VALID_IN                       : in   std_logic;
    GT2_TX_MMCM_LOCK_OUT                    : out  std_logic;
    GT2_RX_MMCM_LOCK_OUT                    : out  std_logic;
    GT3_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT3_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT3_DATA_VALID_IN                       : in   std_logic;
    GT3_TX_MMCM_LOCK_OUT                    : out  std_logic;
    GT3_RX_MMCM_LOCK_OUT                    : out  std_logic;
    GT4_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT4_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT4_DATA_VALID_IN                       : in   std_logic;
    GT4_TX_MMCM_LOCK_OUT                    : out  std_logic;
    GT4_RX_MMCM_LOCK_OUT                    : out  std_logic;
    GT5_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT5_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT5_DATA_VALID_IN                       : in   std_logic;
    GT5_TX_MMCM_LOCK_OUT                    : out  std_logic;
    GT5_RX_MMCM_LOCK_OUT                    : out  std_logic;
    GT6_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT6_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT6_DATA_VALID_IN                       : in   std_logic;
    GT6_TX_MMCM_LOCK_OUT                    : out  std_logic;
    GT6_RX_MMCM_LOCK_OUT                    : out  std_logic;
    GT7_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT7_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT7_DATA_VALID_IN                       : in   std_logic;
    GT7_TX_MMCM_LOCK_OUT                    : out  std_logic;
    GT7_RX_MMCM_LOCK_OUT                    : out  std_logic;
    GT8_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT8_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT8_DATA_VALID_IN                       : in   std_logic;
    GT8_TX_MMCM_LOCK_OUT                    : out  std_logic;
    GT8_RX_MMCM_LOCK_OUT                    : out  std_logic;
    GT9_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT9_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT9_DATA_VALID_IN                       : in   std_logic;
    GT9_TX_MMCM_LOCK_OUT                    : out  std_logic;
    GT9_RX_MMCM_LOCK_OUT                    : out  std_logic;
    GT10_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT10_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT10_DATA_VALID_IN                      : in   std_logic;
    GT10_TX_MMCM_LOCK_OUT                   : out  std_logic;
    GT10_RX_MMCM_LOCK_OUT                   : out  std_logic;
    GT11_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT11_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT11_DATA_VALID_IN                      : in   std_logic;
    GT11_TX_MMCM_LOCK_OUT                   : out  std_logic;
    GT11_RX_MMCM_LOCK_OUT                   : out  std_logic;
    GT12_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT12_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT12_DATA_VALID_IN                      : in   std_logic;
    GT12_TX_MMCM_LOCK_OUT                   : out  std_logic;
    GT12_RX_MMCM_LOCK_OUT                   : out  std_logic;
    GT13_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT13_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT13_DATA_VALID_IN                      : in   std_logic;
    GT13_TX_MMCM_LOCK_OUT                   : out  std_logic;
    GT13_RX_MMCM_LOCK_OUT                   : out  std_logic;
    GT14_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT14_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT14_DATA_VALID_IN                      : in   std_logic;
    GT14_TX_MMCM_LOCK_OUT                   : out  std_logic;
    GT14_RX_MMCM_LOCK_OUT                   : out  std_logic;
    GT15_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT15_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT15_DATA_VALID_IN                      : in   std_logic;
    GT15_TX_MMCM_LOCK_OUT                   : out  std_logic;
    GT15_RX_MMCM_LOCK_OUT                   : out  std_logic;
    GT16_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT16_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT16_DATA_VALID_IN                      : in   std_logic;
    GT16_TX_MMCM_LOCK_OUT                   : out  std_logic;
    GT16_RX_MMCM_LOCK_OUT                   : out  std_logic;
    GT17_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT17_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT17_DATA_VALID_IN                      : in   std_logic;
    GT17_TX_MMCM_LOCK_OUT                   : out  std_logic;
    GT17_RX_MMCM_LOCK_OUT                   : out  std_logic;
    GT18_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT18_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT18_DATA_VALID_IN                      : in   std_logic;
    GT18_TX_MMCM_LOCK_OUT                   : out  std_logic;
    GT18_RX_MMCM_LOCK_OUT                   : out  std_logic;
    GT19_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT19_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT19_DATA_VALID_IN                      : in   std_logic;
    GT19_TX_MMCM_LOCK_OUT                   : out  std_logic;
    GT19_RX_MMCM_LOCK_OUT                   : out  std_logic;
    GT20_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT20_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT20_DATA_VALID_IN                      : in   std_logic;
    GT20_TX_MMCM_LOCK_OUT                   : out  std_logic;
    GT20_RX_MMCM_LOCK_OUT                   : out  std_logic;
    GT21_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT21_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT21_DATA_VALID_IN                      : in   std_logic;
    GT21_TX_MMCM_LOCK_OUT                   : out  std_logic;
    GT21_RX_MMCM_LOCK_OUT                   : out  std_logic;
    GT22_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT22_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT22_DATA_VALID_IN                      : in   std_logic;
    GT22_TX_MMCM_LOCK_OUT                   : out  std_logic;
    GT22_RX_MMCM_LOCK_OUT                   : out  std_logic;
    GT23_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT23_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT23_DATA_VALID_IN                      : in   std_logic;
    GT23_TX_MMCM_LOCK_OUT                   : out  std_logic;
    GT23_RX_MMCM_LOCK_OUT                   : out  std_logic;
    GT24_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT24_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT24_DATA_VALID_IN                      : in   std_logic;
    GT24_TX_MMCM_LOCK_OUT                   : out  std_logic;
    GT24_RX_MMCM_LOCK_OUT                   : out  std_logic;
    GT25_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT25_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT25_DATA_VALID_IN                      : in   std_logic;
    GT25_TX_MMCM_LOCK_OUT                   : out  std_logic;
    GT25_RX_MMCM_LOCK_OUT                   : out  std_logic;
    GT26_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT26_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT26_DATA_VALID_IN                      : in   std_logic;
    GT26_TX_MMCM_LOCK_OUT                   : out  std_logic;
    GT26_RX_MMCM_LOCK_OUT                   : out  std_logic;
    GT27_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT27_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT27_DATA_VALID_IN                      : in   std_logic;
    GT27_TX_MMCM_LOCK_OUT                   : out  std_logic;
    GT27_RX_MMCM_LOCK_OUT                   : out  std_logic;
    GT28_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT28_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT28_DATA_VALID_IN                      : in   std_logic;
    GT28_TX_MMCM_LOCK_OUT                   : out  std_logic;
    GT28_RX_MMCM_LOCK_OUT                   : out  std_logic;
    GT29_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT29_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT29_DATA_VALID_IN                      : in   std_logic;
    GT29_TX_MMCM_LOCK_OUT                   : out  std_logic;
    GT29_RX_MMCM_LOCK_OUT                   : out  std_logic;
    GT30_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT30_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT30_DATA_VALID_IN                      : in   std_logic;
    GT30_TX_MMCM_LOCK_OUT                   : out  std_logic;
    GT30_RX_MMCM_LOCK_OUT                   : out  std_logic;
    GT31_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT31_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT31_DATA_VALID_IN                      : in   std_logic;
    GT31_TX_MMCM_LOCK_OUT                   : out  std_logic;
    GT31_RX_MMCM_LOCK_OUT                   : out  std_logic;
 
    GT0_TXUSRCLK_OUT                        : out  std_logic;
    GT0_TXUSRCLK2_OUT                       : out  std_logic;
    GT0_RXUSRCLK_OUT                        : out  std_logic;
    GT0_RXUSRCLK2_OUT                       : out  std_logic;
 
    GT1_TXUSRCLK_OUT                        : out  std_logic;
    GT1_TXUSRCLK2_OUT                       : out  std_logic;
    GT1_RXUSRCLK_OUT                        : out  std_logic;
    GT1_RXUSRCLK2_OUT                       : out  std_logic;
 
    GT2_TXUSRCLK_OUT                        : out  std_logic;
    GT2_TXUSRCLK2_OUT                       : out  std_logic;
    GT2_RXUSRCLK_OUT                        : out  std_logic;
    GT2_RXUSRCLK2_OUT                       : out  std_logic;
 
    GT3_TXUSRCLK_OUT                        : out  std_logic;
    GT3_TXUSRCLK2_OUT                       : out  std_logic;
    GT3_RXUSRCLK_OUT                        : out  std_logic;
    GT3_RXUSRCLK2_OUT                       : out  std_logic;
 
    GT4_TXUSRCLK_OUT                        : out  std_logic;
    GT4_TXUSRCLK2_OUT                       : out  std_logic;
    GT4_RXUSRCLK_OUT                        : out  std_logic;
    GT4_RXUSRCLK2_OUT                       : out  std_logic;
 
    GT5_TXUSRCLK_OUT                        : out  std_logic;
    GT5_TXUSRCLK2_OUT                       : out  std_logic;
    GT5_RXUSRCLK_OUT                        : out  std_logic;
    GT5_RXUSRCLK2_OUT                       : out  std_logic;
 
    GT6_TXUSRCLK_OUT                        : out  std_logic;
    GT6_TXUSRCLK2_OUT                       : out  std_logic;
    GT6_RXUSRCLK_OUT                        : out  std_logic;
    GT6_RXUSRCLK2_OUT                       : out  std_logic;
 
    GT7_TXUSRCLK_OUT                        : out  std_logic;
    GT7_TXUSRCLK2_OUT                       : out  std_logic;
    GT7_RXUSRCLK_OUT                        : out  std_logic;
    GT7_RXUSRCLK2_OUT                       : out  std_logic;
 
    GT8_TXUSRCLK_OUT                        : out  std_logic;
    GT8_TXUSRCLK2_OUT                       : out  std_logic;
    GT8_RXUSRCLK_OUT                        : out  std_logic;
    GT8_RXUSRCLK2_OUT                       : out  std_logic;
 
    GT9_TXUSRCLK_OUT                        : out  std_logic;
    GT9_TXUSRCLK2_OUT                       : out  std_logic;
    GT9_RXUSRCLK_OUT                        : out  std_logic;
    GT9_RXUSRCLK2_OUT                       : out  std_logic;
 
    GT10_TXUSRCLK_OUT                       : out  std_logic;
    GT10_TXUSRCLK2_OUT                      : out  std_logic;
    GT10_RXUSRCLK_OUT                       : out  std_logic;
    GT10_RXUSRCLK2_OUT                      : out  std_logic;
 
    GT11_TXUSRCLK_OUT                       : out  std_logic;
    GT11_TXUSRCLK2_OUT                      : out  std_logic;
    GT11_RXUSRCLK_OUT                       : out  std_logic;
    GT11_RXUSRCLK2_OUT                      : out  std_logic;
 
    GT12_TXUSRCLK_OUT                       : out  std_logic;
    GT12_TXUSRCLK2_OUT                      : out  std_logic;
    GT12_RXUSRCLK_OUT                       : out  std_logic;
    GT12_RXUSRCLK2_OUT                      : out  std_logic;
 
    GT13_TXUSRCLK_OUT                       : out  std_logic;
    GT13_TXUSRCLK2_OUT                      : out  std_logic;
    GT13_RXUSRCLK_OUT                       : out  std_logic;
    GT13_RXUSRCLK2_OUT                      : out  std_logic;
 
    GT14_TXUSRCLK_OUT                       : out  std_logic;
    GT14_TXUSRCLK2_OUT                      : out  std_logic;
    GT14_RXUSRCLK_OUT                       : out  std_logic;
    GT14_RXUSRCLK2_OUT                      : out  std_logic;
 
    GT15_TXUSRCLK_OUT                       : out  std_logic;
    GT15_TXUSRCLK2_OUT                      : out  std_logic;
    GT15_RXUSRCLK_OUT                       : out  std_logic;
    GT15_RXUSRCLK2_OUT                      : out  std_logic;
 
    GT16_TXUSRCLK_OUT                       : out  std_logic;
    GT16_TXUSRCLK2_OUT                      : out  std_logic;
    GT16_RXUSRCLK_OUT                       : out  std_logic;
    GT16_RXUSRCLK2_OUT                      : out  std_logic;
 
    GT17_TXUSRCLK_OUT                       : out  std_logic;
    GT17_TXUSRCLK2_OUT                      : out  std_logic;
    GT17_RXUSRCLK_OUT                       : out  std_logic;
    GT17_RXUSRCLK2_OUT                      : out  std_logic;
 
    GT18_TXUSRCLK_OUT                       : out  std_logic;
    GT18_TXUSRCLK2_OUT                      : out  std_logic;
    GT18_RXUSRCLK_OUT                       : out  std_logic;
    GT18_RXUSRCLK2_OUT                      : out  std_logic;
 
    GT19_TXUSRCLK_OUT                       : out  std_logic;
    GT19_TXUSRCLK2_OUT                      : out  std_logic;
    GT19_RXUSRCLK_OUT                       : out  std_logic;
    GT19_RXUSRCLK2_OUT                      : out  std_logic;
 
    GT20_TXUSRCLK_OUT                       : out  std_logic;
    GT20_TXUSRCLK2_OUT                      : out  std_logic;
    GT20_RXUSRCLK_OUT                       : out  std_logic;
    GT20_RXUSRCLK2_OUT                      : out  std_logic;
 
    GT21_TXUSRCLK_OUT                       : out  std_logic;
    GT21_TXUSRCLK2_OUT                      : out  std_logic;
    GT21_RXUSRCLK_OUT                       : out  std_logic;
    GT21_RXUSRCLK2_OUT                      : out  std_logic;
 
    GT22_TXUSRCLK_OUT                       : out  std_logic;
    GT22_TXUSRCLK2_OUT                      : out  std_logic;
    GT22_RXUSRCLK_OUT                       : out  std_logic;
    GT22_RXUSRCLK2_OUT                      : out  std_logic;
 
    GT23_TXUSRCLK_OUT                       : out  std_logic;
    GT23_TXUSRCLK2_OUT                      : out  std_logic;
    GT23_RXUSRCLK_OUT                       : out  std_logic;
    GT23_RXUSRCLK2_OUT                      : out  std_logic;
 
    GT24_TXUSRCLK_OUT                       : out  std_logic;
    GT24_TXUSRCLK2_OUT                      : out  std_logic;
    GT24_RXUSRCLK_OUT                       : out  std_logic;
    GT24_RXUSRCLK2_OUT                      : out  std_logic;
 
    GT25_TXUSRCLK_OUT                       : out  std_logic;
    GT25_TXUSRCLK2_OUT                      : out  std_logic;
    GT25_RXUSRCLK_OUT                       : out  std_logic;
    GT25_RXUSRCLK2_OUT                      : out  std_logic;
 
    GT26_TXUSRCLK_OUT                       : out  std_logic;
    GT26_TXUSRCLK2_OUT                      : out  std_logic;
    GT26_RXUSRCLK_OUT                       : out  std_logic;
    GT26_RXUSRCLK2_OUT                      : out  std_logic;
 
    GT27_TXUSRCLK_OUT                       : out  std_logic;
    GT27_TXUSRCLK2_OUT                      : out  std_logic;
    GT27_RXUSRCLK_OUT                       : out  std_logic;
    GT27_RXUSRCLK2_OUT                      : out  std_logic;
 
    GT28_TXUSRCLK_OUT                       : out  std_logic;
    GT28_TXUSRCLK2_OUT                      : out  std_logic;
    GT28_RXUSRCLK_OUT                       : out  std_logic;
    GT28_RXUSRCLK2_OUT                      : out  std_logic;
 
    GT29_TXUSRCLK_OUT                       : out  std_logic;
    GT29_TXUSRCLK2_OUT                      : out  std_logic;
    GT29_RXUSRCLK_OUT                       : out  std_logic;
    GT29_RXUSRCLK2_OUT                      : out  std_logic;
 
    GT30_TXUSRCLK_OUT                       : out  std_logic;
    GT30_TXUSRCLK2_OUT                      : out  std_logic;
    GT30_RXUSRCLK_OUT                       : out  std_logic;
    GT30_RXUSRCLK2_OUT                      : out  std_logic;
 
    GT31_TXUSRCLK_OUT                       : out  std_logic;
    GT31_TXUSRCLK2_OUT                      : out  std_logic;
    GT31_RXUSRCLK_OUT                       : out  std_logic;
    GT31_RXUSRCLK2_OUT                      : out  std_logic;

    --_________________________________________________________________________
    --GT0  (X1Y4)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt0_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt0_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt0_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt0_drpen_in                            : in   std_logic;
    gt0_drprdy_out                          : out  std_logic;
    gt0_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt0_eyescanreset_in                     : in   std_logic;
    gt0_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt0_eyescandataerror_out                : out  std_logic;
    gt0_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt0_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt0_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt0_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt0_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt0_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt0_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt0_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt0_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt0_rxbyteisaligned_out                 : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt0_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt0_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt0_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt0_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt0_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt0_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt0_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt0_gttxreset_in                        : in   std_logic;
    gt0_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt0_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt0_gthtxn_out                          : out  std_logic;
    gt0_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt0_txoutclkfabric_out                  : out  std_logic;
    gt0_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt0_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt0_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT1  (X1Y5)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt1_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt1_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt1_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt1_drpen_in                            : in   std_logic;
    gt1_drprdy_out                          : out  std_logic;
    gt1_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt1_eyescanreset_in                     : in   std_logic;
    gt1_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt1_eyescandataerror_out                : out  std_logic;
    gt1_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt1_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt1_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt1_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt1_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt1_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt1_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt1_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt1_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt1_rxbyteisaligned_out                 : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt1_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt1_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt1_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt1_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt1_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt1_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt1_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt1_gttxreset_in                        : in   std_logic;
    gt1_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt1_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt1_gthtxn_out                          : out  std_logic;
    gt1_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt1_txoutclkfabric_out                  : out  std_logic;
    gt1_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt1_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt1_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT2  (X1Y6)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt2_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt2_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt2_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt2_drpen_in                            : in   std_logic;
    gt2_drprdy_out                          : out  std_logic;
    gt2_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt2_eyescanreset_in                     : in   std_logic;
    gt2_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt2_eyescandataerror_out                : out  std_logic;
    gt2_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt2_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt2_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt2_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt2_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt2_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt2_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt2_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt2_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt2_rxbyteisaligned_out                 : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt2_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt2_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt2_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt2_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt2_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt2_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt2_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt2_gttxreset_in                        : in   std_logic;
    gt2_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt2_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt2_gthtxn_out                          : out  std_logic;
    gt2_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt2_txoutclkfabric_out                  : out  std_logic;
    gt2_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt2_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt2_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT3  (X1Y7)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt3_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt3_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt3_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt3_drpen_in                            : in   std_logic;
    gt3_drprdy_out                          : out  std_logic;
    gt3_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt3_eyescanreset_in                     : in   std_logic;
    gt3_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt3_eyescandataerror_out                : out  std_logic;
    gt3_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt3_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt3_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt3_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt3_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt3_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt3_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt3_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt3_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt3_rxbyteisaligned_out                 : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt3_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt3_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt3_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt3_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt3_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt3_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt3_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt3_gttxreset_in                        : in   std_logic;
    gt3_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt3_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt3_gthtxn_out                          : out  std_logic;
    gt3_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt3_txoutclkfabric_out                  : out  std_logic;
    gt3_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt3_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt3_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT4  (X1Y8)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt4_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt4_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt4_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt4_drpen_in                            : in   std_logic;
    gt4_drprdy_out                          : out  std_logic;
    gt4_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt4_eyescanreset_in                     : in   std_logic;
    gt4_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt4_eyescandataerror_out                : out  std_logic;
    gt4_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt4_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt4_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt4_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt4_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt4_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt4_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt4_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt4_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt4_rxbyteisaligned_out                 : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt4_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt4_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt4_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt4_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt4_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt4_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt4_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt4_gttxreset_in                        : in   std_logic;
    gt4_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt4_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt4_gthtxn_out                          : out  std_logic;
    gt4_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt4_txoutclkfabric_out                  : out  std_logic;
    gt4_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt4_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt4_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT5  (X1Y9)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt5_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt5_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt5_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt5_drpen_in                            : in   std_logic;
    gt5_drprdy_out                          : out  std_logic;
    gt5_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt5_eyescanreset_in                     : in   std_logic;
    gt5_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt5_eyescandataerror_out                : out  std_logic;
    gt5_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt5_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt5_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt5_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt5_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt5_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt5_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt5_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt5_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt5_rxbyteisaligned_out                 : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt5_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt5_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt5_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt5_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt5_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt5_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt5_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt5_gttxreset_in                        : in   std_logic;
    gt5_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt5_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt5_gthtxn_out                          : out  std_logic;
    gt5_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt5_txoutclkfabric_out                  : out  std_logic;
    gt5_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt5_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt5_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT6  (X1Y10)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt6_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt6_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt6_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt6_drpen_in                            : in   std_logic;
    gt6_drprdy_out                          : out  std_logic;
    gt6_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt6_eyescanreset_in                     : in   std_logic;
    gt6_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt6_eyescandataerror_out                : out  std_logic;
    gt6_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt6_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt6_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt6_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt6_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt6_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt6_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt6_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt6_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt6_rxbyteisaligned_out                 : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt6_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt6_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt6_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt6_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt6_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt6_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt6_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt6_gttxreset_in                        : in   std_logic;
    gt6_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt6_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt6_gthtxn_out                          : out  std_logic;
    gt6_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt6_txoutclkfabric_out                  : out  std_logic;
    gt6_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt6_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt6_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT7  (X1Y11)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt7_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt7_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt7_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt7_drpen_in                            : in   std_logic;
    gt7_drprdy_out                          : out  std_logic;
    gt7_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt7_eyescanreset_in                     : in   std_logic;
    gt7_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt7_eyescandataerror_out                : out  std_logic;
    gt7_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt7_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt7_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt7_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt7_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt7_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt7_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt7_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt7_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt7_rxbyteisaligned_out                 : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt7_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt7_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt7_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt7_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt7_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt7_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt7_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt7_gttxreset_in                        : in   std_logic;
    gt7_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt7_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt7_gthtxn_out                          : out  std_logic;
    gt7_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt7_txoutclkfabric_out                  : out  std_logic;
    gt7_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt7_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt7_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT8  (X1Y12)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt8_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt8_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt8_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt8_drpen_in                            : in   std_logic;
    gt8_drprdy_out                          : out  std_logic;
    gt8_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt8_eyescanreset_in                     : in   std_logic;
    gt8_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt8_eyescandataerror_out                : out  std_logic;
    gt8_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt8_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt8_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt8_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt8_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt8_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt8_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt8_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt8_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt8_rxbyteisaligned_out                 : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt8_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt8_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt8_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt8_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt8_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt8_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt8_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt8_gttxreset_in                        : in   std_logic;
    gt8_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt8_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt8_gthtxn_out                          : out  std_logic;
    gt8_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt8_txoutclkfabric_out                  : out  std_logic;
    gt8_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt8_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt8_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT9  (X1Y13)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt9_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt9_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt9_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt9_drpen_in                            : in   std_logic;
    gt9_drprdy_out                          : out  std_logic;
    gt9_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt9_eyescanreset_in                     : in   std_logic;
    gt9_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt9_eyescandataerror_out                : out  std_logic;
    gt9_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt9_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt9_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt9_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt9_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt9_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt9_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt9_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt9_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt9_rxbyteisaligned_out                 : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt9_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt9_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt9_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt9_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt9_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt9_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt9_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt9_gttxreset_in                        : in   std_logic;
    gt9_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt9_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt9_gthtxn_out                          : out  std_logic;
    gt9_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt9_txoutclkfabric_out                  : out  std_logic;
    gt9_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt9_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt9_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT10  (X1Y14)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt10_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt10_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt10_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt10_drpen_in                           : in   std_logic;
    gt10_drprdy_out                         : out  std_logic;
    gt10_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt10_eyescanreset_in                    : in   std_logic;
    gt10_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt10_eyescandataerror_out               : out  std_logic;
    gt10_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt10_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt10_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt10_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt10_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt10_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt10_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt10_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt10_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt10_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt10_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt10_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt10_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt10_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt10_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt10_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt10_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt10_gttxreset_in                       : in   std_logic;
    gt10_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt10_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt10_gthtxn_out                         : out  std_logic;
    gt10_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt10_txoutclkfabric_out                 : out  std_logic;
    gt10_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt10_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt10_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT11  (X1Y15)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt11_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt11_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt11_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt11_drpen_in                           : in   std_logic;
    gt11_drprdy_out                         : out  std_logic;
    gt11_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt11_eyescanreset_in                    : in   std_logic;
    gt11_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt11_eyescandataerror_out               : out  std_logic;
    gt11_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt11_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt11_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt11_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt11_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt11_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt11_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt11_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt11_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt11_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt11_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt11_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt11_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt11_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt11_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt11_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt11_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt11_gttxreset_in                       : in   std_logic;
    gt11_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt11_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt11_gthtxn_out                         : out  std_logic;
    gt11_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt11_txoutclkfabric_out                 : out  std_logic;
    gt11_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt11_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt11_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT12  (X1Y16)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt12_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt12_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt12_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt12_drpen_in                           : in   std_logic;
    gt12_drprdy_out                         : out  std_logic;
    gt12_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt12_eyescanreset_in                    : in   std_logic;
    gt12_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt12_eyescandataerror_out               : out  std_logic;
    gt12_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt12_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt12_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt12_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt12_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt12_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt12_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt12_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt12_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt12_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt12_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt12_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt12_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt12_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt12_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt12_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt12_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt12_gttxreset_in                       : in   std_logic;
    gt12_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt12_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt12_gthtxn_out                         : out  std_logic;
    gt12_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt12_txoutclkfabric_out                 : out  std_logic;
    gt12_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt12_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt12_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT13  (X1Y17)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt13_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt13_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt13_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt13_drpen_in                           : in   std_logic;
    gt13_drprdy_out                         : out  std_logic;
    gt13_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt13_eyescanreset_in                    : in   std_logic;
    gt13_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt13_eyescandataerror_out               : out  std_logic;
    gt13_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt13_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt13_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt13_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt13_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt13_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt13_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt13_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt13_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt13_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt13_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt13_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt13_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt13_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt13_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt13_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt13_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt13_gttxreset_in                       : in   std_logic;
    gt13_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt13_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt13_gthtxn_out                         : out  std_logic;
    gt13_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt13_txoutclkfabric_out                 : out  std_logic;
    gt13_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt13_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt13_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT14  (X1Y18)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt14_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt14_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt14_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt14_drpen_in                           : in   std_logic;
    gt14_drprdy_out                         : out  std_logic;
    gt14_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt14_eyescanreset_in                    : in   std_logic;
    gt14_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt14_eyescandataerror_out               : out  std_logic;
    gt14_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt14_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt14_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt14_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt14_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt14_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt14_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt14_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt14_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt14_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt14_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt14_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt14_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt14_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt14_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt14_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt14_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt14_gttxreset_in                       : in   std_logic;
    gt14_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt14_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt14_gthtxn_out                         : out  std_logic;
    gt14_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt14_txoutclkfabric_out                 : out  std_logic;
    gt14_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt14_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt14_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT15  (X1Y19)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt15_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt15_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt15_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt15_drpen_in                           : in   std_logic;
    gt15_drprdy_out                         : out  std_logic;
    gt15_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt15_eyescanreset_in                    : in   std_logic;
    gt15_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt15_eyescandataerror_out               : out  std_logic;
    gt15_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt15_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt15_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt15_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt15_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt15_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt15_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt15_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt15_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt15_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt15_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt15_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt15_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt15_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt15_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt15_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt15_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt15_gttxreset_in                       : in   std_logic;
    gt15_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt15_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt15_gthtxn_out                         : out  std_logic;
    gt15_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt15_txoutclkfabric_out                 : out  std_logic;
    gt15_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt15_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt15_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT16  (X1Y20)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt16_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt16_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt16_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt16_drpen_in                           : in   std_logic;
    gt16_drprdy_out                         : out  std_logic;
    gt16_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt16_eyescanreset_in                    : in   std_logic;
    gt16_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt16_eyescandataerror_out               : out  std_logic;
    gt16_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt16_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt16_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt16_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt16_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt16_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt16_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt16_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt16_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt16_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt16_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt16_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt16_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt16_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt16_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt16_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt16_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt16_gttxreset_in                       : in   std_logic;
    gt16_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt16_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt16_gthtxn_out                         : out  std_logic;
    gt16_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt16_txoutclkfabric_out                 : out  std_logic;
    gt16_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt16_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt16_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT17  (X1Y21)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt17_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt17_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt17_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt17_drpen_in                           : in   std_logic;
    gt17_drprdy_out                         : out  std_logic;
    gt17_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt17_eyescanreset_in                    : in   std_logic;
    gt17_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt17_eyescandataerror_out               : out  std_logic;
    gt17_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt17_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt17_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt17_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt17_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt17_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt17_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt17_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt17_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt17_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt17_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt17_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt17_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt17_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt17_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt17_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt17_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt17_gttxreset_in                       : in   std_logic;
    gt17_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt17_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt17_gthtxn_out                         : out  std_logic;
    gt17_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt17_txoutclkfabric_out                 : out  std_logic;
    gt17_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt17_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt17_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT18  (X1Y22)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt18_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt18_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt18_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt18_drpen_in                           : in   std_logic;
    gt18_drprdy_out                         : out  std_logic;
    gt18_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt18_eyescanreset_in                    : in   std_logic;
    gt18_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt18_eyescandataerror_out               : out  std_logic;
    gt18_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt18_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt18_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt18_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt18_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt18_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt18_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt18_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt18_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt18_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt18_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt18_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt18_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt18_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt18_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt18_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt18_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt18_gttxreset_in                       : in   std_logic;
    gt18_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt18_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt18_gthtxn_out                         : out  std_logic;
    gt18_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt18_txoutclkfabric_out                 : out  std_logic;
    gt18_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt18_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt18_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT19  (X1Y23)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt19_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt19_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt19_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt19_drpen_in                           : in   std_logic;
    gt19_drprdy_out                         : out  std_logic;
    gt19_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt19_eyescanreset_in                    : in   std_logic;
    gt19_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt19_eyescandataerror_out               : out  std_logic;
    gt19_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt19_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt19_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt19_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt19_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt19_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt19_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt19_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt19_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt19_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt19_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt19_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt19_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt19_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt19_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt19_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt19_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt19_gttxreset_in                       : in   std_logic;
    gt19_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt19_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt19_gthtxn_out                         : out  std_logic;
    gt19_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt19_txoutclkfabric_out                 : out  std_logic;
    gt19_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt19_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt19_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT20  (X1Y24)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt20_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt20_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt20_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt20_drpen_in                           : in   std_logic;
    gt20_drprdy_out                         : out  std_logic;
    gt20_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt20_eyescanreset_in                    : in   std_logic;
    gt20_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt20_eyescandataerror_out               : out  std_logic;
    gt20_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt20_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt20_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt20_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt20_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt20_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt20_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt20_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt20_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt20_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt20_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt20_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt20_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt20_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt20_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt20_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt20_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt20_gttxreset_in                       : in   std_logic;
    gt20_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt20_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt20_gthtxn_out                         : out  std_logic;
    gt20_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt20_txoutclkfabric_out                 : out  std_logic;
    gt20_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt20_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt20_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT21  (X1Y25)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt21_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt21_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt21_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt21_drpen_in                           : in   std_logic;
    gt21_drprdy_out                         : out  std_logic;
    gt21_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt21_eyescanreset_in                    : in   std_logic;
    gt21_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt21_eyescandataerror_out               : out  std_logic;
    gt21_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt21_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt21_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt21_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt21_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt21_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt21_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt21_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt21_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt21_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt21_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt21_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt21_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt21_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt21_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt21_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt21_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt21_gttxreset_in                       : in   std_logic;
    gt21_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt21_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt21_gthtxn_out                         : out  std_logic;
    gt21_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt21_txoutclkfabric_out                 : out  std_logic;
    gt21_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt21_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt21_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT22  (X1Y26)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt22_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt22_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt22_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt22_drpen_in                           : in   std_logic;
    gt22_drprdy_out                         : out  std_logic;
    gt22_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt22_eyescanreset_in                    : in   std_logic;
    gt22_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt22_eyescandataerror_out               : out  std_logic;
    gt22_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt22_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt22_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt22_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt22_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt22_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt22_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt22_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt22_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt22_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt22_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt22_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt22_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt22_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt22_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt22_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt22_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt22_gttxreset_in                       : in   std_logic;
    gt22_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt22_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt22_gthtxn_out                         : out  std_logic;
    gt22_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt22_txoutclkfabric_out                 : out  std_logic;
    gt22_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt22_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt22_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT23  (X1Y27)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt23_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt23_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt23_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt23_drpen_in                           : in   std_logic;
    gt23_drprdy_out                         : out  std_logic;
    gt23_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt23_eyescanreset_in                    : in   std_logic;
    gt23_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt23_eyescandataerror_out               : out  std_logic;
    gt23_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt23_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt23_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt23_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt23_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt23_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt23_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt23_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt23_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt23_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt23_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt23_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt23_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt23_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt23_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt23_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt23_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt23_gttxreset_in                       : in   std_logic;
    gt23_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt23_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt23_gthtxn_out                         : out  std_logic;
    gt23_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt23_txoutclkfabric_out                 : out  std_logic;
    gt23_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt23_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt23_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT24  (X1Y28)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt24_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt24_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt24_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt24_drpen_in                           : in   std_logic;
    gt24_drprdy_out                         : out  std_logic;
    gt24_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt24_eyescanreset_in                    : in   std_logic;
    gt24_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt24_eyescandataerror_out               : out  std_logic;
    gt24_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt24_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt24_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt24_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt24_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt24_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt24_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt24_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt24_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt24_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt24_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt24_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt24_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt24_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt24_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt24_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt24_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt24_gttxreset_in                       : in   std_logic;
    gt24_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt24_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt24_gthtxn_out                         : out  std_logic;
    gt24_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt24_txoutclkfabric_out                 : out  std_logic;
    gt24_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt24_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt24_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT25  (X1Y29)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt25_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt25_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt25_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt25_drpen_in                           : in   std_logic;
    gt25_drprdy_out                         : out  std_logic;
    gt25_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt25_eyescanreset_in                    : in   std_logic;
    gt25_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt25_eyescandataerror_out               : out  std_logic;
    gt25_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt25_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt25_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt25_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt25_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt25_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt25_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt25_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt25_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt25_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt25_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt25_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt25_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt25_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt25_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt25_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt25_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt25_gttxreset_in                       : in   std_logic;
    gt25_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt25_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt25_gthtxn_out                         : out  std_logic;
    gt25_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt25_txoutclkfabric_out                 : out  std_logic;
    gt25_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt25_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt25_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT26  (X1Y30)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt26_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt26_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt26_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt26_drpen_in                           : in   std_logic;
    gt26_drprdy_out                         : out  std_logic;
    gt26_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt26_eyescanreset_in                    : in   std_logic;
    gt26_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt26_eyescandataerror_out               : out  std_logic;
    gt26_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt26_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt26_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt26_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt26_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt26_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt26_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt26_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt26_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt26_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt26_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt26_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt26_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt26_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt26_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt26_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt26_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt26_gttxreset_in                       : in   std_logic;
    gt26_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt26_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt26_gthtxn_out                         : out  std_logic;
    gt26_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt26_txoutclkfabric_out                 : out  std_logic;
    gt26_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt26_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt26_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT27  (X1Y31)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt27_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt27_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt27_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt27_drpen_in                           : in   std_logic;
    gt27_drprdy_out                         : out  std_logic;
    gt27_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt27_eyescanreset_in                    : in   std_logic;
    gt27_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt27_eyescandataerror_out               : out  std_logic;
    gt27_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt27_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt27_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt27_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt27_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt27_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt27_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt27_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt27_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt27_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt27_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt27_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt27_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt27_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt27_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt27_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt27_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt27_gttxreset_in                       : in   std_logic;
    gt27_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt27_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt27_gthtxn_out                         : out  std_logic;
    gt27_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt27_txoutclkfabric_out                 : out  std_logic;
    gt27_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt27_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt27_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT28  (X1Y32)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt28_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt28_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt28_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt28_drpen_in                           : in   std_logic;
    gt28_drprdy_out                         : out  std_logic;
    gt28_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt28_eyescanreset_in                    : in   std_logic;
    gt28_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt28_eyescandataerror_out               : out  std_logic;
    gt28_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt28_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt28_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt28_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt28_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt28_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt28_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt28_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt28_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt28_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt28_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt28_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt28_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt28_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt28_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt28_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt28_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt28_gttxreset_in                       : in   std_logic;
    gt28_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt28_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt28_gthtxn_out                         : out  std_logic;
    gt28_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt28_txoutclkfabric_out                 : out  std_logic;
    gt28_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt28_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt28_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT29  (X1Y33)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt29_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt29_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt29_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt29_drpen_in                           : in   std_logic;
    gt29_drprdy_out                         : out  std_logic;
    gt29_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt29_eyescanreset_in                    : in   std_logic;
    gt29_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt29_eyescandataerror_out               : out  std_logic;
    gt29_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt29_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt29_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt29_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt29_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt29_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt29_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt29_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt29_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt29_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt29_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt29_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt29_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt29_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt29_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt29_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt29_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt29_gttxreset_in                       : in   std_logic;
    gt29_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt29_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt29_gthtxn_out                         : out  std_logic;
    gt29_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt29_txoutclkfabric_out                 : out  std_logic;
    gt29_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt29_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt29_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT30  (X1Y34)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt30_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt30_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt30_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt30_drpen_in                           : in   std_logic;
    gt30_drprdy_out                         : out  std_logic;
    gt30_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt30_eyescanreset_in                    : in   std_logic;
    gt30_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt30_eyescandataerror_out               : out  std_logic;
    gt30_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt30_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt30_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt30_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt30_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt30_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt30_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt30_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt30_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt30_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt30_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt30_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt30_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt30_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt30_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt30_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt30_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt30_gttxreset_in                       : in   std_logic;
    gt30_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt30_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt30_gthtxn_out                         : out  std_logic;
    gt30_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt30_txoutclkfabric_out                 : out  std_logic;
    gt30_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt30_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt30_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT31  (X1Y35)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt31_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt31_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt31_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt31_drpen_in                           : in   std_logic;
    gt31_drprdy_out                         : out  std_logic;
    gt31_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt31_eyescanreset_in                    : in   std_logic;
    gt31_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt31_eyescandataerror_out               : out  std_logic;
    gt31_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt31_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt31_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt31_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt31_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt31_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt31_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt31_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt31_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt31_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt31_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt31_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt31_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt31_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt31_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt31_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt31_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt31_gttxreset_in                       : in   std_logic;
    gt31_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt31_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt31_gthtxn_out                         : out  std_logic;
    gt31_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt31_txoutclkfabric_out                 : out  std_logic;
    gt31_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt31_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt31_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --____________________________COMMON PORTS________________________________
    GT0_QPLLLOCK_OUT : out std_logic;
    GT0_QPLLREFCLKLOST_OUT  : out std_logic;
    GT0_QPLLRESET_OUT  : out std_logic;
     GT0_QPLLOUTCLK_OUT  : out std_logic;
     GT0_QPLLOUTREFCLK_OUT : out std_logic;
    --____________________________COMMON PORTS________________________________
    GT1_QPLLLOCK_OUT : out std_logic;
    GT1_QPLLREFCLKLOST_OUT  : out std_logic;
    GT1_QPLLRESET_OUT  : out std_logic;
     GT1_QPLLOUTCLK_OUT  : out std_logic;
     GT1_QPLLOUTREFCLK_OUT : out std_logic;
    --____________________________COMMON PORTS________________________________
    GT2_QPLLLOCK_OUT : out std_logic;
    GT2_QPLLREFCLKLOST_OUT  : out std_logic;
    GT2_QPLLRESET_OUT  : out std_logic;
     GT2_QPLLOUTCLK_OUT  : out std_logic;
     GT2_QPLLOUTREFCLK_OUT : out std_logic;
    --____________________________COMMON PORTS________________________________
    GT3_QPLLLOCK_OUT : out std_logic;
    GT3_QPLLREFCLKLOST_OUT  : out std_logic;
    GT3_QPLLRESET_OUT  : out std_logic;
     GT3_QPLLOUTCLK_OUT  : out std_logic;
     GT3_QPLLOUTREFCLK_OUT : out std_logic;
    --____________________________COMMON PORTS________________________________
    GT4_QPLLLOCK_OUT : out std_logic;
    GT4_QPLLREFCLKLOST_OUT  : out std_logic;
    GT4_QPLLRESET_OUT  : out std_logic;
     GT4_QPLLOUTCLK_OUT  : out std_logic;
     GT4_QPLLOUTREFCLK_OUT : out std_logic;
    --____________________________COMMON PORTS________________________________
    GT5_QPLLLOCK_OUT : out std_logic;
    GT5_QPLLREFCLKLOST_OUT  : out std_logic;
    GT5_QPLLRESET_OUT  : out std_logic;
     GT5_QPLLOUTCLK_OUT  : out std_logic;
     GT5_QPLLOUTREFCLK_OUT : out std_logic;
    --____________________________COMMON PORTS________________________________
    GT6_QPLLLOCK_OUT : out std_logic;
    GT6_QPLLREFCLKLOST_OUT  : out std_logic;
    GT6_QPLLRESET_OUT  : out std_logic;
     GT6_QPLLOUTCLK_OUT  : out std_logic;
     GT6_QPLLOUTREFCLK_OUT : out std_logic;
    --____________________________COMMON PORTS________________________________
    GT7_QPLLLOCK_OUT : out std_logic;
    GT7_QPLLREFCLKLOST_OUT  : out std_logic;
    GT7_QPLLRESET_OUT  : out std_logic;
     GT7_QPLLOUTCLK_OUT  : out std_logic;
     GT7_QPLLOUTREFCLK_OUT : out std_logic;
       sysclk_in        : in std_logic

);

end gtwizard_0_support;
    
architecture RTL of gtwizard_0_support is
attribute DowngradeIPIdentifiedWarnings: string;
attribute DowngradeIPIdentifiedWarnings of RTL : architecture is "yes";

--**************************Component Declarations*****************************

component gtwizard_0_init
 
port
(
    SYSCLK_IN                               : in   std_logic;
    SOFT_RESET_TX_IN                        : in   std_logic;
    SOFT_RESET_RX_IN                        : in   std_logic;
    DONT_RESET_ON_DATA_ERROR_IN             : in   std_logic;
    GT0_DRP_BUSY_OUT                        : out  std_logic;
    GT0_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_DATA_VALID_IN                       : in   std_logic;
    GT0_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT0_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT0_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT0_RX_MMCM_RESET_OUT                   : out  std_logic;
    GT1_DRP_BUSY_OUT                        : out  std_logic;
    GT1_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT1_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT1_DATA_VALID_IN                       : in   std_logic;
    GT1_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT1_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT1_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT1_RX_MMCM_RESET_OUT                   : out  std_logic;
    GT2_DRP_BUSY_OUT                        : out  std_logic;
    GT2_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT2_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT2_DATA_VALID_IN                       : in   std_logic;
    GT2_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT2_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT2_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT2_RX_MMCM_RESET_OUT                   : out  std_logic;
    GT3_DRP_BUSY_OUT                        : out  std_logic;
    GT3_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT3_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT3_DATA_VALID_IN                       : in   std_logic;
    GT3_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT3_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT3_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT3_RX_MMCM_RESET_OUT                   : out  std_logic;
    GT4_DRP_BUSY_OUT                        : out  std_logic;
    GT4_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT4_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT4_DATA_VALID_IN                       : in   std_logic;
    GT4_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT4_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT4_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT4_RX_MMCM_RESET_OUT                   : out  std_logic;
    GT5_DRP_BUSY_OUT                        : out  std_logic;
    GT5_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT5_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT5_DATA_VALID_IN                       : in   std_logic;
    GT5_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT5_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT5_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT5_RX_MMCM_RESET_OUT                   : out  std_logic;
    GT6_DRP_BUSY_OUT                        : out  std_logic;
    GT6_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT6_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT6_DATA_VALID_IN                       : in   std_logic;
    GT6_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT6_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT6_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT6_RX_MMCM_RESET_OUT                   : out  std_logic;
    GT7_DRP_BUSY_OUT                        : out  std_logic;
    GT7_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT7_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT7_DATA_VALID_IN                       : in   std_logic;
    GT7_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT7_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT7_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT7_RX_MMCM_RESET_OUT                   : out  std_logic;
    GT8_DRP_BUSY_OUT                        : out  std_logic;
    GT8_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT8_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT8_DATA_VALID_IN                       : in   std_logic;
    GT8_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT8_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT8_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT8_RX_MMCM_RESET_OUT                   : out  std_logic;
    GT9_DRP_BUSY_OUT                        : out  std_logic;
    GT9_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT9_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT9_DATA_VALID_IN                       : in   std_logic;
    GT9_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT9_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT9_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT9_RX_MMCM_RESET_OUT                   : out  std_logic;
    GT10_DRP_BUSY_OUT                       : out  std_logic;
    GT10_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT10_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT10_DATA_VALID_IN                      : in   std_logic;
    GT10_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT10_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT10_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT10_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT11_DRP_BUSY_OUT                       : out  std_logic;
    GT11_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT11_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT11_DATA_VALID_IN                      : in   std_logic;
    GT11_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT11_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT11_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT11_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT12_DRP_BUSY_OUT                       : out  std_logic;
    GT12_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT12_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT12_DATA_VALID_IN                      : in   std_logic;
    GT12_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT12_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT12_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT12_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT13_DRP_BUSY_OUT                       : out  std_logic;
    GT13_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT13_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT13_DATA_VALID_IN                      : in   std_logic;
    GT13_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT13_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT13_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT13_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT14_DRP_BUSY_OUT                       : out  std_logic;
    GT14_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT14_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT14_DATA_VALID_IN                      : in   std_logic;
    GT14_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT14_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT14_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT14_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT15_DRP_BUSY_OUT                       : out  std_logic;
    GT15_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT15_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT15_DATA_VALID_IN                      : in   std_logic;
    GT15_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT15_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT15_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT15_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT16_DRP_BUSY_OUT                       : out  std_logic;
    GT16_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT16_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT16_DATA_VALID_IN                      : in   std_logic;
    GT16_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT16_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT16_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT16_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT17_DRP_BUSY_OUT                       : out  std_logic;
    GT17_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT17_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT17_DATA_VALID_IN                      : in   std_logic;
    GT17_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT17_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT17_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT17_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT18_DRP_BUSY_OUT                       : out  std_logic;
    GT18_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT18_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT18_DATA_VALID_IN                      : in   std_logic;
    GT18_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT18_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT18_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT18_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT19_DRP_BUSY_OUT                       : out  std_logic;
    GT19_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT19_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT19_DATA_VALID_IN                      : in   std_logic;
    GT19_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT19_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT19_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT19_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT20_DRP_BUSY_OUT                       : out  std_logic;
    GT20_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT20_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT20_DATA_VALID_IN                      : in   std_logic;
    GT20_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT20_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT20_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT20_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT21_DRP_BUSY_OUT                       : out  std_logic;
    GT21_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT21_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT21_DATA_VALID_IN                      : in   std_logic;
    GT21_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT21_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT21_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT21_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT22_DRP_BUSY_OUT                       : out  std_logic;
    GT22_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT22_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT22_DATA_VALID_IN                      : in   std_logic;
    GT22_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT22_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT22_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT22_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT23_DRP_BUSY_OUT                       : out  std_logic;
    GT23_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT23_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT23_DATA_VALID_IN                      : in   std_logic;
    GT23_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT23_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT23_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT23_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT24_DRP_BUSY_OUT                       : out  std_logic;
    GT24_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT24_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT24_DATA_VALID_IN                      : in   std_logic;
    GT24_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT24_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT24_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT24_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT25_DRP_BUSY_OUT                       : out  std_logic;
    GT25_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT25_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT25_DATA_VALID_IN                      : in   std_logic;
    GT25_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT25_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT25_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT25_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT26_DRP_BUSY_OUT                       : out  std_logic;
    GT26_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT26_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT26_DATA_VALID_IN                      : in   std_logic;
    GT26_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT26_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT26_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT26_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT27_DRP_BUSY_OUT                       : out  std_logic;
    GT27_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT27_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT27_DATA_VALID_IN                      : in   std_logic;
    GT27_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT27_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT27_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT27_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT28_DRP_BUSY_OUT                       : out  std_logic;
    GT28_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT28_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT28_DATA_VALID_IN                      : in   std_logic;
    GT28_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT28_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT28_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT28_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT29_DRP_BUSY_OUT                       : out  std_logic;
    GT29_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT29_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT29_DATA_VALID_IN                      : in   std_logic;
    GT29_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT29_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT29_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT29_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT30_DRP_BUSY_OUT                       : out  std_logic;
    GT30_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT30_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT30_DATA_VALID_IN                      : in   std_logic;
    GT30_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT30_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT30_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT30_RX_MMCM_RESET_OUT                  : out  std_logic;
    GT31_DRP_BUSY_OUT                       : out  std_logic;
    GT31_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT31_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT31_DATA_VALID_IN                      : in   std_logic;
    GT31_TX_MMCM_LOCK_IN                    : in   std_logic;
    GT31_TX_MMCM_RESET_OUT                  : out  std_logic;
    GT31_RX_MMCM_LOCK_IN                    : in   std_logic;
    GT31_RX_MMCM_RESET_OUT                  : out  std_logic;

    --_________________________________________________________________________
    --GT0  (X1Y4)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt0_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt0_drpclk_in                           : in   std_logic;
    gt0_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt0_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt0_drpen_in                            : in   std_logic;
    gt0_drprdy_out                          : out  std_logic;
    gt0_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt0_eyescanreset_in                     : in   std_logic;
    gt0_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt0_eyescandataerror_out                : out  std_logic;
    gt0_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt0_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt0_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt0_rxusrclk_in                         : in   std_logic;
    gt0_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt0_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt0_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt0_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt0_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt0_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt0_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt0_rxbyteisaligned_out                 : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt0_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt0_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt0_rxoutclk_out                        : out  std_logic;
    gt0_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt0_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt0_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt0_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt0_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt0_gttxreset_in                        : in   std_logic;
    gt0_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt0_txusrclk_in                         : in   std_logic;
    gt0_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt0_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt0_gthtxn_out                          : out  std_logic;
    gt0_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt0_txoutclk_out                        : out  std_logic;
    gt0_txoutclkfabric_out                  : out  std_logic;
    gt0_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt0_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt0_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT1  (X1Y5)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt1_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt1_drpclk_in                           : in   std_logic;
    gt1_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt1_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt1_drpen_in                            : in   std_logic;
    gt1_drprdy_out                          : out  std_logic;
    gt1_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt1_eyescanreset_in                     : in   std_logic;
    gt1_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt1_eyescandataerror_out                : out  std_logic;
    gt1_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt1_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt1_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt1_rxusrclk_in                         : in   std_logic;
    gt1_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt1_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt1_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt1_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt1_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt1_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt1_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt1_rxbyteisaligned_out                 : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt1_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt1_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt1_rxoutclk_out                        : out  std_logic;
    gt1_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt1_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt1_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt1_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt1_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt1_gttxreset_in                        : in   std_logic;
    gt1_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt1_txusrclk_in                         : in   std_logic;
    gt1_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt1_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt1_gthtxn_out                          : out  std_logic;
    gt1_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt1_txoutclk_out                        : out  std_logic;
    gt1_txoutclkfabric_out                  : out  std_logic;
    gt1_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt1_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt1_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT2  (X1Y6)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt2_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt2_drpclk_in                           : in   std_logic;
    gt2_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt2_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt2_drpen_in                            : in   std_logic;
    gt2_drprdy_out                          : out  std_logic;
    gt2_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt2_eyescanreset_in                     : in   std_logic;
    gt2_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt2_eyescandataerror_out                : out  std_logic;
    gt2_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt2_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt2_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt2_rxusrclk_in                         : in   std_logic;
    gt2_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt2_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt2_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt2_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt2_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt2_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt2_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt2_rxbyteisaligned_out                 : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt2_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt2_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt2_rxoutclk_out                        : out  std_logic;
    gt2_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt2_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt2_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt2_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt2_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt2_gttxreset_in                        : in   std_logic;
    gt2_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt2_txusrclk_in                         : in   std_logic;
    gt2_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt2_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt2_gthtxn_out                          : out  std_logic;
    gt2_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt2_txoutclk_out                        : out  std_logic;
    gt2_txoutclkfabric_out                  : out  std_logic;
    gt2_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt2_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt2_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT3  (X1Y7)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt3_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt3_drpclk_in                           : in   std_logic;
    gt3_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt3_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt3_drpen_in                            : in   std_logic;
    gt3_drprdy_out                          : out  std_logic;
    gt3_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt3_eyescanreset_in                     : in   std_logic;
    gt3_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt3_eyescandataerror_out                : out  std_logic;
    gt3_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt3_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt3_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt3_rxusrclk_in                         : in   std_logic;
    gt3_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt3_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt3_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt3_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt3_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt3_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt3_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt3_rxbyteisaligned_out                 : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt3_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt3_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt3_rxoutclk_out                        : out  std_logic;
    gt3_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt3_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt3_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt3_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt3_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt3_gttxreset_in                        : in   std_logic;
    gt3_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt3_txusrclk_in                         : in   std_logic;
    gt3_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt3_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt3_gthtxn_out                          : out  std_logic;
    gt3_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt3_txoutclk_out                        : out  std_logic;
    gt3_txoutclkfabric_out                  : out  std_logic;
    gt3_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt3_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt3_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT4  (X1Y8)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt4_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt4_drpclk_in                           : in   std_logic;
    gt4_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt4_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt4_drpen_in                            : in   std_logic;
    gt4_drprdy_out                          : out  std_logic;
    gt4_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt4_eyescanreset_in                     : in   std_logic;
    gt4_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt4_eyescandataerror_out                : out  std_logic;
    gt4_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt4_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt4_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt4_rxusrclk_in                         : in   std_logic;
    gt4_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt4_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt4_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt4_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt4_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt4_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt4_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt4_rxbyteisaligned_out                 : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt4_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt4_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt4_rxoutclk_out                        : out  std_logic;
    gt4_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt4_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt4_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt4_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt4_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt4_gttxreset_in                        : in   std_logic;
    gt4_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt4_txusrclk_in                         : in   std_logic;
    gt4_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt4_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt4_gthtxn_out                          : out  std_logic;
    gt4_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt4_txoutclk_out                        : out  std_logic;
    gt4_txoutclkfabric_out                  : out  std_logic;
    gt4_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt4_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt4_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT5  (X1Y9)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt5_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt5_drpclk_in                           : in   std_logic;
    gt5_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt5_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt5_drpen_in                            : in   std_logic;
    gt5_drprdy_out                          : out  std_logic;
    gt5_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt5_eyescanreset_in                     : in   std_logic;
    gt5_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt5_eyescandataerror_out                : out  std_logic;
    gt5_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt5_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt5_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt5_rxusrclk_in                         : in   std_logic;
    gt5_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt5_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt5_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt5_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt5_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt5_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt5_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt5_rxbyteisaligned_out                 : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt5_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt5_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt5_rxoutclk_out                        : out  std_logic;
    gt5_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt5_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt5_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt5_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt5_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt5_gttxreset_in                        : in   std_logic;
    gt5_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt5_txusrclk_in                         : in   std_logic;
    gt5_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt5_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt5_gthtxn_out                          : out  std_logic;
    gt5_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt5_txoutclk_out                        : out  std_logic;
    gt5_txoutclkfabric_out                  : out  std_logic;
    gt5_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt5_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt5_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT6  (X1Y10)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt6_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt6_drpclk_in                           : in   std_logic;
    gt6_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt6_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt6_drpen_in                            : in   std_logic;
    gt6_drprdy_out                          : out  std_logic;
    gt6_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt6_eyescanreset_in                     : in   std_logic;
    gt6_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt6_eyescandataerror_out                : out  std_logic;
    gt6_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt6_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt6_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt6_rxusrclk_in                         : in   std_logic;
    gt6_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt6_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt6_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt6_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt6_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt6_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt6_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt6_rxbyteisaligned_out                 : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt6_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt6_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt6_rxoutclk_out                        : out  std_logic;
    gt6_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt6_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt6_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt6_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt6_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt6_gttxreset_in                        : in   std_logic;
    gt6_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt6_txusrclk_in                         : in   std_logic;
    gt6_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt6_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt6_gthtxn_out                          : out  std_logic;
    gt6_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt6_txoutclk_out                        : out  std_logic;
    gt6_txoutclkfabric_out                  : out  std_logic;
    gt6_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt6_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt6_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT7  (X1Y11)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt7_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt7_drpclk_in                           : in   std_logic;
    gt7_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt7_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt7_drpen_in                            : in   std_logic;
    gt7_drprdy_out                          : out  std_logic;
    gt7_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt7_eyescanreset_in                     : in   std_logic;
    gt7_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt7_eyescandataerror_out                : out  std_logic;
    gt7_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt7_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt7_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt7_rxusrclk_in                         : in   std_logic;
    gt7_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt7_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt7_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt7_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt7_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt7_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt7_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt7_rxbyteisaligned_out                 : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt7_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt7_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt7_rxoutclk_out                        : out  std_logic;
    gt7_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt7_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt7_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt7_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt7_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt7_gttxreset_in                        : in   std_logic;
    gt7_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt7_txusrclk_in                         : in   std_logic;
    gt7_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt7_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt7_gthtxn_out                          : out  std_logic;
    gt7_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt7_txoutclk_out                        : out  std_logic;
    gt7_txoutclkfabric_out                  : out  std_logic;
    gt7_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt7_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt7_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT8  (X1Y12)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt8_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt8_drpclk_in                           : in   std_logic;
    gt8_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt8_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt8_drpen_in                            : in   std_logic;
    gt8_drprdy_out                          : out  std_logic;
    gt8_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt8_eyescanreset_in                     : in   std_logic;
    gt8_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt8_eyescandataerror_out                : out  std_logic;
    gt8_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt8_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt8_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt8_rxusrclk_in                         : in   std_logic;
    gt8_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt8_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt8_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt8_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt8_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt8_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt8_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt8_rxbyteisaligned_out                 : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt8_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt8_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt8_rxoutclk_out                        : out  std_logic;
    gt8_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt8_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt8_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt8_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt8_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt8_gttxreset_in                        : in   std_logic;
    gt8_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt8_txusrclk_in                         : in   std_logic;
    gt8_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt8_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt8_gthtxn_out                          : out  std_logic;
    gt8_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt8_txoutclk_out                        : out  std_logic;
    gt8_txoutclkfabric_out                  : out  std_logic;
    gt8_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt8_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt8_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT9  (X1Y13)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt9_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt9_drpclk_in                           : in   std_logic;
    gt9_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt9_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt9_drpen_in                            : in   std_logic;
    gt9_drprdy_out                          : out  std_logic;
    gt9_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt9_eyescanreset_in                     : in   std_logic;
    gt9_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt9_eyescandataerror_out                : out  std_logic;
    gt9_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt9_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt9_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt9_rxusrclk_in                         : in   std_logic;
    gt9_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt9_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt9_rxdisperr_out                       : out  std_logic_vector(7 downto 0);
    gt9_rxnotintable_out                    : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt9_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt9_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt9_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt9_rxbyteisaligned_out                 : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt9_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt9_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt9_rxoutclk_out                        : out  std_logic;
    gt9_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt9_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt9_rxcharisk_out                       : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt9_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt9_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt9_gttxreset_in                        : in   std_logic;
    gt9_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt9_txusrclk_in                         : in   std_logic;
    gt9_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt9_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt9_gthtxn_out                          : out  std_logic;
    gt9_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt9_txoutclk_out                        : out  std_logic;
    gt9_txoutclkfabric_out                  : out  std_logic;
    gt9_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt9_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt9_txcharisk_in                        : in   std_logic_vector(7 downto 0);

    --GT10  (X1Y14)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt10_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt10_drpclk_in                          : in   std_logic;
    gt10_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt10_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt10_drpen_in                           : in   std_logic;
    gt10_drprdy_out                         : out  std_logic;
    gt10_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt10_eyescanreset_in                    : in   std_logic;
    gt10_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt10_eyescandataerror_out               : out  std_logic;
    gt10_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt10_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt10_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt10_rxusrclk_in                        : in   std_logic;
    gt10_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt10_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt10_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt10_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt10_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt10_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt10_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt10_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt10_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt10_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt10_rxoutclk_out                       : out  std_logic;
    gt10_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt10_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt10_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt10_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt10_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt10_gttxreset_in                       : in   std_logic;
    gt10_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt10_txusrclk_in                        : in   std_logic;
    gt10_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt10_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt10_gthtxn_out                         : out  std_logic;
    gt10_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt10_txoutclk_out                       : out  std_logic;
    gt10_txoutclkfabric_out                 : out  std_logic;
    gt10_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt10_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt10_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT11  (X1Y15)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt11_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt11_drpclk_in                          : in   std_logic;
    gt11_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt11_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt11_drpen_in                           : in   std_logic;
    gt11_drprdy_out                         : out  std_logic;
    gt11_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt11_eyescanreset_in                    : in   std_logic;
    gt11_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt11_eyescandataerror_out               : out  std_logic;
    gt11_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt11_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt11_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt11_rxusrclk_in                        : in   std_logic;
    gt11_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt11_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt11_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt11_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt11_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt11_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt11_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt11_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt11_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt11_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt11_rxoutclk_out                       : out  std_logic;
    gt11_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt11_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt11_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt11_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt11_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt11_gttxreset_in                       : in   std_logic;
    gt11_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt11_txusrclk_in                        : in   std_logic;
    gt11_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt11_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt11_gthtxn_out                         : out  std_logic;
    gt11_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt11_txoutclk_out                       : out  std_logic;
    gt11_txoutclkfabric_out                 : out  std_logic;
    gt11_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt11_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt11_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT12  (X1Y16)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt12_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt12_drpclk_in                          : in   std_logic;
    gt12_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt12_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt12_drpen_in                           : in   std_logic;
    gt12_drprdy_out                         : out  std_logic;
    gt12_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt12_eyescanreset_in                    : in   std_logic;
    gt12_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt12_eyescandataerror_out               : out  std_logic;
    gt12_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt12_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt12_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt12_rxusrclk_in                        : in   std_logic;
    gt12_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt12_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt12_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt12_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt12_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt12_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt12_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt12_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt12_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt12_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt12_rxoutclk_out                       : out  std_logic;
    gt12_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt12_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt12_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt12_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt12_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt12_gttxreset_in                       : in   std_logic;
    gt12_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt12_txusrclk_in                        : in   std_logic;
    gt12_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt12_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt12_gthtxn_out                         : out  std_logic;
    gt12_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt12_txoutclk_out                       : out  std_logic;
    gt12_txoutclkfabric_out                 : out  std_logic;
    gt12_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt12_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt12_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT13  (X1Y17)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt13_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt13_drpclk_in                          : in   std_logic;
    gt13_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt13_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt13_drpen_in                           : in   std_logic;
    gt13_drprdy_out                         : out  std_logic;
    gt13_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt13_eyescanreset_in                    : in   std_logic;
    gt13_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt13_eyescandataerror_out               : out  std_logic;
    gt13_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt13_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt13_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt13_rxusrclk_in                        : in   std_logic;
    gt13_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt13_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt13_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt13_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt13_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt13_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt13_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt13_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt13_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt13_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt13_rxoutclk_out                       : out  std_logic;
    gt13_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt13_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt13_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt13_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt13_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt13_gttxreset_in                       : in   std_logic;
    gt13_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt13_txusrclk_in                        : in   std_logic;
    gt13_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt13_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt13_gthtxn_out                         : out  std_logic;
    gt13_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt13_txoutclk_out                       : out  std_logic;
    gt13_txoutclkfabric_out                 : out  std_logic;
    gt13_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt13_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt13_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT14  (X1Y18)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt14_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt14_drpclk_in                          : in   std_logic;
    gt14_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt14_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt14_drpen_in                           : in   std_logic;
    gt14_drprdy_out                         : out  std_logic;
    gt14_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt14_eyescanreset_in                    : in   std_logic;
    gt14_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt14_eyescandataerror_out               : out  std_logic;
    gt14_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt14_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt14_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt14_rxusrclk_in                        : in   std_logic;
    gt14_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt14_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt14_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt14_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt14_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt14_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt14_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt14_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt14_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt14_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt14_rxoutclk_out                       : out  std_logic;
    gt14_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt14_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt14_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt14_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt14_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt14_gttxreset_in                       : in   std_logic;
    gt14_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt14_txusrclk_in                        : in   std_logic;
    gt14_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt14_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt14_gthtxn_out                         : out  std_logic;
    gt14_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt14_txoutclk_out                       : out  std_logic;
    gt14_txoutclkfabric_out                 : out  std_logic;
    gt14_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt14_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt14_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT15  (X1Y19)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt15_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt15_drpclk_in                          : in   std_logic;
    gt15_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt15_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt15_drpen_in                           : in   std_logic;
    gt15_drprdy_out                         : out  std_logic;
    gt15_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt15_eyescanreset_in                    : in   std_logic;
    gt15_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt15_eyescandataerror_out               : out  std_logic;
    gt15_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt15_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt15_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt15_rxusrclk_in                        : in   std_logic;
    gt15_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt15_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt15_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt15_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt15_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt15_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt15_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt15_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt15_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt15_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt15_rxoutclk_out                       : out  std_logic;
    gt15_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt15_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt15_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt15_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt15_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt15_gttxreset_in                       : in   std_logic;
    gt15_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt15_txusrclk_in                        : in   std_logic;
    gt15_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt15_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt15_gthtxn_out                         : out  std_logic;
    gt15_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt15_txoutclk_out                       : out  std_logic;
    gt15_txoutclkfabric_out                 : out  std_logic;
    gt15_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt15_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt15_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT16  (X1Y20)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt16_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt16_drpclk_in                          : in   std_logic;
    gt16_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt16_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt16_drpen_in                           : in   std_logic;
    gt16_drprdy_out                         : out  std_logic;
    gt16_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt16_eyescanreset_in                    : in   std_logic;
    gt16_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt16_eyescandataerror_out               : out  std_logic;
    gt16_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt16_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt16_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt16_rxusrclk_in                        : in   std_logic;
    gt16_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt16_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt16_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt16_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt16_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt16_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt16_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt16_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt16_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt16_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt16_rxoutclk_out                       : out  std_logic;
    gt16_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt16_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt16_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt16_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt16_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt16_gttxreset_in                       : in   std_logic;
    gt16_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt16_txusrclk_in                        : in   std_logic;
    gt16_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt16_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt16_gthtxn_out                         : out  std_logic;
    gt16_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt16_txoutclk_out                       : out  std_logic;
    gt16_txoutclkfabric_out                 : out  std_logic;
    gt16_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt16_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt16_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT17  (X1Y21)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt17_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt17_drpclk_in                          : in   std_logic;
    gt17_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt17_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt17_drpen_in                           : in   std_logic;
    gt17_drprdy_out                         : out  std_logic;
    gt17_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt17_eyescanreset_in                    : in   std_logic;
    gt17_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt17_eyescandataerror_out               : out  std_logic;
    gt17_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt17_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt17_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt17_rxusrclk_in                        : in   std_logic;
    gt17_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt17_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt17_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt17_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt17_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt17_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt17_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt17_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt17_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt17_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt17_rxoutclk_out                       : out  std_logic;
    gt17_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt17_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt17_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt17_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt17_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt17_gttxreset_in                       : in   std_logic;
    gt17_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt17_txusrclk_in                        : in   std_logic;
    gt17_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt17_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt17_gthtxn_out                         : out  std_logic;
    gt17_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt17_txoutclk_out                       : out  std_logic;
    gt17_txoutclkfabric_out                 : out  std_logic;
    gt17_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt17_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt17_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT18  (X1Y22)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt18_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt18_drpclk_in                          : in   std_logic;
    gt18_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt18_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt18_drpen_in                           : in   std_logic;
    gt18_drprdy_out                         : out  std_logic;
    gt18_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt18_eyescanreset_in                    : in   std_logic;
    gt18_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt18_eyescandataerror_out               : out  std_logic;
    gt18_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt18_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt18_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt18_rxusrclk_in                        : in   std_logic;
    gt18_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt18_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt18_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt18_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt18_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt18_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt18_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt18_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt18_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt18_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt18_rxoutclk_out                       : out  std_logic;
    gt18_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt18_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt18_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt18_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt18_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt18_gttxreset_in                       : in   std_logic;
    gt18_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt18_txusrclk_in                        : in   std_logic;
    gt18_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt18_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt18_gthtxn_out                         : out  std_logic;
    gt18_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt18_txoutclk_out                       : out  std_logic;
    gt18_txoutclkfabric_out                 : out  std_logic;
    gt18_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt18_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt18_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT19  (X1Y23)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt19_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt19_drpclk_in                          : in   std_logic;
    gt19_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt19_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt19_drpen_in                           : in   std_logic;
    gt19_drprdy_out                         : out  std_logic;
    gt19_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt19_eyescanreset_in                    : in   std_logic;
    gt19_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt19_eyescandataerror_out               : out  std_logic;
    gt19_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt19_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt19_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt19_rxusrclk_in                        : in   std_logic;
    gt19_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt19_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt19_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt19_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt19_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt19_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt19_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt19_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt19_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt19_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt19_rxoutclk_out                       : out  std_logic;
    gt19_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt19_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt19_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt19_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt19_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt19_gttxreset_in                       : in   std_logic;
    gt19_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt19_txusrclk_in                        : in   std_logic;
    gt19_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt19_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt19_gthtxn_out                         : out  std_logic;
    gt19_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt19_txoutclk_out                       : out  std_logic;
    gt19_txoutclkfabric_out                 : out  std_logic;
    gt19_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt19_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt19_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT20  (X1Y24)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt20_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt20_drpclk_in                          : in   std_logic;
    gt20_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt20_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt20_drpen_in                           : in   std_logic;
    gt20_drprdy_out                         : out  std_logic;
    gt20_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt20_eyescanreset_in                    : in   std_logic;
    gt20_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt20_eyescandataerror_out               : out  std_logic;
    gt20_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt20_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt20_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt20_rxusrclk_in                        : in   std_logic;
    gt20_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt20_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt20_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt20_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt20_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt20_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt20_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt20_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt20_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt20_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt20_rxoutclk_out                       : out  std_logic;
    gt20_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt20_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt20_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt20_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt20_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt20_gttxreset_in                       : in   std_logic;
    gt20_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt20_txusrclk_in                        : in   std_logic;
    gt20_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt20_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt20_gthtxn_out                         : out  std_logic;
    gt20_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt20_txoutclk_out                       : out  std_logic;
    gt20_txoutclkfabric_out                 : out  std_logic;
    gt20_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt20_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt20_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT21  (X1Y25)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt21_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt21_drpclk_in                          : in   std_logic;
    gt21_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt21_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt21_drpen_in                           : in   std_logic;
    gt21_drprdy_out                         : out  std_logic;
    gt21_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt21_eyescanreset_in                    : in   std_logic;
    gt21_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt21_eyescandataerror_out               : out  std_logic;
    gt21_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt21_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt21_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt21_rxusrclk_in                        : in   std_logic;
    gt21_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt21_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt21_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt21_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt21_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt21_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt21_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt21_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt21_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt21_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt21_rxoutclk_out                       : out  std_logic;
    gt21_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt21_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt21_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt21_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt21_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt21_gttxreset_in                       : in   std_logic;
    gt21_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt21_txusrclk_in                        : in   std_logic;
    gt21_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt21_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt21_gthtxn_out                         : out  std_logic;
    gt21_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt21_txoutclk_out                       : out  std_logic;
    gt21_txoutclkfabric_out                 : out  std_logic;
    gt21_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt21_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt21_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT22  (X1Y26)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt22_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt22_drpclk_in                          : in   std_logic;
    gt22_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt22_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt22_drpen_in                           : in   std_logic;
    gt22_drprdy_out                         : out  std_logic;
    gt22_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt22_eyescanreset_in                    : in   std_logic;
    gt22_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt22_eyescandataerror_out               : out  std_logic;
    gt22_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt22_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt22_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt22_rxusrclk_in                        : in   std_logic;
    gt22_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt22_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt22_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt22_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt22_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt22_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt22_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt22_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt22_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt22_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt22_rxoutclk_out                       : out  std_logic;
    gt22_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt22_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt22_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt22_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt22_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt22_gttxreset_in                       : in   std_logic;
    gt22_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt22_txusrclk_in                        : in   std_logic;
    gt22_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt22_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt22_gthtxn_out                         : out  std_logic;
    gt22_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt22_txoutclk_out                       : out  std_logic;
    gt22_txoutclkfabric_out                 : out  std_logic;
    gt22_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt22_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt22_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT23  (X1Y27)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt23_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt23_drpclk_in                          : in   std_logic;
    gt23_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt23_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt23_drpen_in                           : in   std_logic;
    gt23_drprdy_out                         : out  std_logic;
    gt23_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt23_eyescanreset_in                    : in   std_logic;
    gt23_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt23_eyescandataerror_out               : out  std_logic;
    gt23_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt23_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt23_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt23_rxusrclk_in                        : in   std_logic;
    gt23_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt23_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt23_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt23_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt23_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt23_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt23_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt23_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt23_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt23_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt23_rxoutclk_out                       : out  std_logic;
    gt23_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt23_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt23_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt23_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt23_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt23_gttxreset_in                       : in   std_logic;
    gt23_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt23_txusrclk_in                        : in   std_logic;
    gt23_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt23_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt23_gthtxn_out                         : out  std_logic;
    gt23_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt23_txoutclk_out                       : out  std_logic;
    gt23_txoutclkfabric_out                 : out  std_logic;
    gt23_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt23_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt23_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT24  (X1Y28)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt24_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt24_drpclk_in                          : in   std_logic;
    gt24_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt24_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt24_drpen_in                           : in   std_logic;
    gt24_drprdy_out                         : out  std_logic;
    gt24_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt24_eyescanreset_in                    : in   std_logic;
    gt24_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt24_eyescandataerror_out               : out  std_logic;
    gt24_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt24_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt24_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt24_rxusrclk_in                        : in   std_logic;
    gt24_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt24_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt24_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt24_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt24_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt24_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt24_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt24_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt24_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt24_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt24_rxoutclk_out                       : out  std_logic;
    gt24_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt24_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt24_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt24_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt24_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt24_gttxreset_in                       : in   std_logic;
    gt24_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt24_txusrclk_in                        : in   std_logic;
    gt24_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt24_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt24_gthtxn_out                         : out  std_logic;
    gt24_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt24_txoutclk_out                       : out  std_logic;
    gt24_txoutclkfabric_out                 : out  std_logic;
    gt24_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt24_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt24_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT25  (X1Y29)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt25_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt25_drpclk_in                          : in   std_logic;
    gt25_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt25_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt25_drpen_in                           : in   std_logic;
    gt25_drprdy_out                         : out  std_logic;
    gt25_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt25_eyescanreset_in                    : in   std_logic;
    gt25_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt25_eyescandataerror_out               : out  std_logic;
    gt25_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt25_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt25_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt25_rxusrclk_in                        : in   std_logic;
    gt25_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt25_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt25_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt25_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt25_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt25_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt25_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt25_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt25_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt25_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt25_rxoutclk_out                       : out  std_logic;
    gt25_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt25_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt25_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt25_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt25_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt25_gttxreset_in                       : in   std_logic;
    gt25_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt25_txusrclk_in                        : in   std_logic;
    gt25_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt25_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt25_gthtxn_out                         : out  std_logic;
    gt25_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt25_txoutclk_out                       : out  std_logic;
    gt25_txoutclkfabric_out                 : out  std_logic;
    gt25_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt25_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt25_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT26  (X1Y30)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt26_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt26_drpclk_in                          : in   std_logic;
    gt26_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt26_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt26_drpen_in                           : in   std_logic;
    gt26_drprdy_out                         : out  std_logic;
    gt26_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt26_eyescanreset_in                    : in   std_logic;
    gt26_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt26_eyescandataerror_out               : out  std_logic;
    gt26_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt26_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt26_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt26_rxusrclk_in                        : in   std_logic;
    gt26_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt26_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt26_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt26_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt26_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt26_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt26_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt26_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt26_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt26_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt26_rxoutclk_out                       : out  std_logic;
    gt26_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt26_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt26_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt26_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt26_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt26_gttxreset_in                       : in   std_logic;
    gt26_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt26_txusrclk_in                        : in   std_logic;
    gt26_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt26_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt26_gthtxn_out                         : out  std_logic;
    gt26_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt26_txoutclk_out                       : out  std_logic;
    gt26_txoutclkfabric_out                 : out  std_logic;
    gt26_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt26_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt26_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT27  (X1Y31)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt27_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt27_drpclk_in                          : in   std_logic;
    gt27_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt27_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt27_drpen_in                           : in   std_logic;
    gt27_drprdy_out                         : out  std_logic;
    gt27_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt27_eyescanreset_in                    : in   std_logic;
    gt27_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt27_eyescandataerror_out               : out  std_logic;
    gt27_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt27_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt27_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt27_rxusrclk_in                        : in   std_logic;
    gt27_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt27_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt27_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt27_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt27_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt27_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt27_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt27_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt27_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt27_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt27_rxoutclk_out                       : out  std_logic;
    gt27_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt27_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt27_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt27_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt27_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt27_gttxreset_in                       : in   std_logic;
    gt27_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt27_txusrclk_in                        : in   std_logic;
    gt27_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt27_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt27_gthtxn_out                         : out  std_logic;
    gt27_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt27_txoutclk_out                       : out  std_logic;
    gt27_txoutclkfabric_out                 : out  std_logic;
    gt27_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt27_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt27_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT28  (X1Y32)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt28_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt28_drpclk_in                          : in   std_logic;
    gt28_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt28_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt28_drpen_in                           : in   std_logic;
    gt28_drprdy_out                         : out  std_logic;
    gt28_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt28_eyescanreset_in                    : in   std_logic;
    gt28_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt28_eyescandataerror_out               : out  std_logic;
    gt28_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt28_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt28_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt28_rxusrclk_in                        : in   std_logic;
    gt28_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt28_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt28_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt28_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt28_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt28_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt28_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt28_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt28_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt28_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt28_rxoutclk_out                       : out  std_logic;
    gt28_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt28_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt28_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt28_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt28_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt28_gttxreset_in                       : in   std_logic;
    gt28_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt28_txusrclk_in                        : in   std_logic;
    gt28_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt28_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt28_gthtxn_out                         : out  std_logic;
    gt28_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt28_txoutclk_out                       : out  std_logic;
    gt28_txoutclkfabric_out                 : out  std_logic;
    gt28_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt28_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt28_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT29  (X1Y33)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt29_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt29_drpclk_in                          : in   std_logic;
    gt29_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt29_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt29_drpen_in                           : in   std_logic;
    gt29_drprdy_out                         : out  std_logic;
    gt29_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt29_eyescanreset_in                    : in   std_logic;
    gt29_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt29_eyescandataerror_out               : out  std_logic;
    gt29_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt29_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt29_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt29_rxusrclk_in                        : in   std_logic;
    gt29_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt29_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt29_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt29_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt29_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt29_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt29_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt29_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt29_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt29_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt29_rxoutclk_out                       : out  std_logic;
    gt29_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt29_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt29_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt29_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt29_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt29_gttxreset_in                       : in   std_logic;
    gt29_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt29_txusrclk_in                        : in   std_logic;
    gt29_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt29_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt29_gthtxn_out                         : out  std_logic;
    gt29_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt29_txoutclk_out                       : out  std_logic;
    gt29_txoutclkfabric_out                 : out  std_logic;
    gt29_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt29_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt29_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT30  (X1Y34)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt30_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt30_drpclk_in                          : in   std_logic;
    gt30_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt30_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt30_drpen_in                           : in   std_logic;
    gt30_drprdy_out                         : out  std_logic;
    gt30_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt30_eyescanreset_in                    : in   std_logic;
    gt30_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt30_eyescandataerror_out               : out  std_logic;
    gt30_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt30_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt30_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt30_rxusrclk_in                        : in   std_logic;
    gt30_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt30_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt30_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt30_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt30_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt30_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt30_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt30_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt30_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt30_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt30_rxoutclk_out                       : out  std_logic;
    gt30_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt30_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt30_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt30_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt30_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt30_gttxreset_in                       : in   std_logic;
    gt30_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt30_txusrclk_in                        : in   std_logic;
    gt30_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt30_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt30_gthtxn_out                         : out  std_logic;
    gt30_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt30_txoutclk_out                       : out  std_logic;
    gt30_txoutclkfabric_out                 : out  std_logic;
    gt30_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt30_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt30_txcharisk_in                       : in   std_logic_vector(7 downto 0);

    --GT31  (X1Y35)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt31_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt31_drpclk_in                          : in   std_logic;
    gt31_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt31_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt31_drpen_in                           : in   std_logic;
    gt31_drprdy_out                         : out  std_logic;
    gt31_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt31_eyescanreset_in                    : in   std_logic;
    gt31_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt31_eyescandataerror_out               : out  std_logic;
    gt31_eyescantrigger_in                  : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt31_rxslide_in                         : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt31_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt31_rxusrclk_in                        : in   std_logic;
    gt31_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt31_rxdata_out                         : out  std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt31_rxdisperr_out                      : out  std_logic_vector(7 downto 0);
    gt31_rxnotintable_out                   : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt31_gthrxn_in                          : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt31_rxphmonitor_out                    : out  std_logic_vector(4 downto 0);
    gt31_rxphslipmonitor_out                : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt31_rxbyteisaligned_out                : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt31_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt31_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt31_rxoutclk_out                       : out  std_logic;
    gt31_rxoutclkfabric_out                 : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt31_gtrxreset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt31_rxcharisk_out                      : out  std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt31_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt31_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt31_gttxreset_in                       : in   std_logic;
    gt31_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt31_txusrclk_in                        : in   std_logic;
    gt31_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt31_txdata_in                          : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt31_gthtxn_out                         : out  std_logic;
    gt31_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt31_txoutclk_out                       : out  std_logic;
    gt31_txoutclkfabric_out                 : out  std_logic;
    gt31_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt31_txresetdone_out                    : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt31_txcharisk_in                       : in   std_logic_vector(7 downto 0);


    --____________________________COMMON PORTS________________________________
    GT0_QPLLLOCK_IN : in std_logic;
    GT0_QPLLREFCLKLOST_IN  : in std_logic;
    GT0_QPLLRESET_OUT  : out std_logic;
     GT0_QPLLOUTCLK_IN  : in std_logic;
     GT0_QPLLOUTREFCLK_IN : in std_logic;
    --____________________________COMMON PORTS________________________________
    GT1_QPLLLOCK_IN : in std_logic;
    GT1_QPLLREFCLKLOST_IN  : in std_logic;
    GT1_QPLLRESET_OUT  : out std_logic;
     GT1_QPLLOUTCLK_IN  : in std_logic;
     GT1_QPLLOUTREFCLK_IN : in std_logic;
    --____________________________COMMON PORTS________________________________
    GT2_QPLLLOCK_IN : in std_logic;
    GT2_QPLLREFCLKLOST_IN  : in std_logic;
    GT2_QPLLRESET_OUT  : out std_logic;
     GT2_QPLLOUTCLK_IN  : in std_logic;
     GT2_QPLLOUTREFCLK_IN : in std_logic;
    --____________________________COMMON PORTS________________________________
    GT3_QPLLLOCK_IN : in std_logic;
    GT3_QPLLREFCLKLOST_IN  : in std_logic;
    GT3_QPLLRESET_OUT  : out std_logic;
     GT3_QPLLOUTCLK_IN  : in std_logic;
     GT3_QPLLOUTREFCLK_IN : in std_logic;
    --____________________________COMMON PORTS________________________________
    GT4_QPLLLOCK_IN : in std_logic;
    GT4_QPLLREFCLKLOST_IN  : in std_logic;
    GT4_QPLLRESET_OUT  : out std_logic;
     GT4_QPLLOUTCLK_IN  : in std_logic;
     GT4_QPLLOUTREFCLK_IN : in std_logic;
    --____________________________COMMON PORTS________________________________
    GT5_QPLLLOCK_IN : in std_logic;
    GT5_QPLLREFCLKLOST_IN  : in std_logic;
    GT5_QPLLRESET_OUT  : out std_logic;
     GT5_QPLLOUTCLK_IN  : in std_logic;
     GT5_QPLLOUTREFCLK_IN : in std_logic;
    --____________________________COMMON PORTS________________________________
    GT6_QPLLLOCK_IN : in std_logic;
    GT6_QPLLREFCLKLOST_IN  : in std_logic;
    GT6_QPLLRESET_OUT  : out std_logic;
     GT6_QPLLOUTCLK_IN  : in std_logic;
     GT6_QPLLOUTREFCLK_IN : in std_logic;
    --____________________________COMMON PORTS________________________________
    GT7_QPLLLOCK_IN : in std_logic;
    GT7_QPLLREFCLKLOST_IN  : in std_logic;
    GT7_QPLLRESET_OUT  : out std_logic;
     GT7_QPLLOUTCLK_IN  : in std_logic;
     GT7_QPLLOUTREFCLK_IN : in std_logic

);

end component;

component gtwizard_0_common_reset  
generic
(
      STABLE_CLOCK_PERIOD      : integer := 8        -- Period of the stable clock driving this state-machine, unit is [ns]
   );
port
   (    
      STABLE_CLOCK             : in std_logic;             --Stable Clock, either a stable clock from the PCB
      SOFT_RESET               : in std_logic;               --User Reset, can be pulled any time
      COMMON_RESET             : out std_logic  --Reset QPLL
   );
end component;

component gtwizard_0_common 
generic
(
    -- Simulation attributes
    WRAPPER_SIM_GTRESET_SPEEDUP     : string     :=  "FALSE" ;       -- Set to "TRUE" to speed up sim reset
    SIM_QPLLREFCLK_SEL              :bit_vector  := "001"
 
);
port
(
    QPLLREFCLKSEL_IN   : in std_logic_vector(2 downto 0);
    GTREFCLK0_IN : in std_logic;
    GTREFCLK1_IN      : in std_logic;
    QPLLLOCK_OUT : out std_logic;
    QPLLLOCKDETCLK_IN : in std_logic;
    QPLLOUTCLK_OUT : out std_logic;
    QPLLOUTREFCLK_OUT : out std_logic;
    QPLLREFCLKLOST_OUT : out std_logic;    
    QPLLRESET_IN : in std_logic

);

end component;

component gtwizard_0_GT_USRCLK_SOURCE 
port
(
    txusrclk2_in : in std_logic;
    txusrclk_in : in std_logic;
    GT0_TXUSRCLK_OUT             : out std_logic;
    GT0_TXUSRCLK2_OUT            : out std_logic;
    GT0_TXOUTCLK_IN              : in  std_logic;
    GT0_TXCLK_LOCK_OUT           : out std_logic;
    GT0_TX_MMCM_RESET_IN         : in std_logic;
    GT0_RXUSRCLK_OUT             : out std_logic;
    GT0_RXUSRCLK2_OUT            : out std_logic;
    GT0_RXOUTCLK_IN              : in  std_logic;
    GT0_RXCLK_LOCK_OUT           : out std_logic;
    GT0_RX_MMCM_RESET_IN         : in std_logic;
 
    GT1_TXUSRCLK_OUT             : out std_logic;
    GT1_TXUSRCLK2_OUT            : out std_logic;
    GT1_TXOUTCLK_IN              : in  std_logic;
    GT1_TXCLK_LOCK_OUT           : out std_logic;
    GT1_TX_MMCM_RESET_IN         : in std_logic;
    GT1_RXUSRCLK_OUT             : out std_logic;
    GT1_RXUSRCLK2_OUT            : out std_logic;
    GT1_RXOUTCLK_IN              : in  std_logic;
    GT1_RXCLK_LOCK_OUT           : out std_logic;
    GT1_RX_MMCM_RESET_IN         : in std_logic;
 
    GT2_TXUSRCLK_OUT             : out std_logic;
    GT2_TXUSRCLK2_OUT            : out std_logic;
    GT2_TXOUTCLK_IN              : in  std_logic;
    GT2_TXCLK_LOCK_OUT           : out std_logic;
    GT2_TX_MMCM_RESET_IN         : in std_logic;
    GT2_RXUSRCLK_OUT             : out std_logic;
    GT2_RXUSRCLK2_OUT            : out std_logic;
    GT2_RXOUTCLK_IN              : in  std_logic;
    GT2_RXCLK_LOCK_OUT           : out std_logic;
    GT2_RX_MMCM_RESET_IN         : in std_logic;
 
    GT3_TXUSRCLK_OUT             : out std_logic;
    GT3_TXUSRCLK2_OUT            : out std_logic;
    GT3_TXOUTCLK_IN              : in  std_logic;
    GT3_TXCLK_LOCK_OUT           : out std_logic;
    GT3_TX_MMCM_RESET_IN         : in std_logic;
    GT3_RXUSRCLK_OUT             : out std_logic;
    GT3_RXUSRCLK2_OUT            : out std_logic;
    GT3_RXOUTCLK_IN              : in  std_logic;
    GT3_RXCLK_LOCK_OUT           : out std_logic;
    GT3_RX_MMCM_RESET_IN         : in std_logic;
 
    GT4_TXUSRCLK_OUT             : out std_logic;
    GT4_TXUSRCLK2_OUT            : out std_logic;
    GT4_TXOUTCLK_IN              : in  std_logic;
    GT4_TXCLK_LOCK_OUT           : out std_logic;
    GT4_TX_MMCM_RESET_IN         : in std_logic;
    GT4_RXUSRCLK_OUT             : out std_logic;
    GT4_RXUSRCLK2_OUT            : out std_logic;
    GT4_RXOUTCLK_IN              : in  std_logic;
    GT4_RXCLK_LOCK_OUT           : out std_logic;
    GT4_RX_MMCM_RESET_IN         : in std_logic;
 
    GT5_TXUSRCLK_OUT             : out std_logic;
    GT5_TXUSRCLK2_OUT            : out std_logic;
    GT5_TXOUTCLK_IN              : in  std_logic;
    GT5_TXCLK_LOCK_OUT           : out std_logic;
    GT5_TX_MMCM_RESET_IN         : in std_logic;
    GT5_RXUSRCLK_OUT             : out std_logic;
    GT5_RXUSRCLK2_OUT            : out std_logic;
    GT5_RXOUTCLK_IN              : in  std_logic;
    GT5_RXCLK_LOCK_OUT           : out std_logic;
    GT5_RX_MMCM_RESET_IN         : in std_logic;
 
    GT6_TXUSRCLK_OUT             : out std_logic;
    GT6_TXUSRCLK2_OUT            : out std_logic;
    GT6_TXOUTCLK_IN              : in  std_logic;
    GT6_TXCLK_LOCK_OUT           : out std_logic;
    GT6_TX_MMCM_RESET_IN         : in std_logic;
    GT6_RXUSRCLK_OUT             : out std_logic;
    GT6_RXUSRCLK2_OUT            : out std_logic;
    GT6_RXOUTCLK_IN              : in  std_logic;
    GT6_RXCLK_LOCK_OUT           : out std_logic;
    GT6_RX_MMCM_RESET_IN         : in std_logic;
 
    GT7_TXUSRCLK_OUT             : out std_logic;
    GT7_TXUSRCLK2_OUT            : out std_logic;
    GT7_TXOUTCLK_IN              : in  std_logic;
    GT7_TXCLK_LOCK_OUT           : out std_logic;
    GT7_TX_MMCM_RESET_IN         : in std_logic;
    GT7_RXUSRCLK_OUT             : out std_logic;
    GT7_RXUSRCLK2_OUT            : out std_logic;
    GT7_RXOUTCLK_IN              : in  std_logic;
    GT7_RXCLK_LOCK_OUT           : out std_logic;
    GT7_RX_MMCM_RESET_IN         : in std_logic;
 
    GT8_TXUSRCLK_OUT             : out std_logic;
    GT8_TXUSRCLK2_OUT            : out std_logic;
    GT8_TXOUTCLK_IN              : in  std_logic;
    GT8_TXCLK_LOCK_OUT           : out std_logic;
    GT8_TX_MMCM_RESET_IN         : in std_logic;
    GT8_RXUSRCLK_OUT             : out std_logic;
    GT8_RXUSRCLK2_OUT            : out std_logic;
    GT8_RXOUTCLK_IN              : in  std_logic;
    GT8_RXCLK_LOCK_OUT           : out std_logic;
    GT8_RX_MMCM_RESET_IN         : in std_logic;
 
    GT9_TXUSRCLK_OUT             : out std_logic;
    GT9_TXUSRCLK2_OUT            : out std_logic;
    GT9_TXOUTCLK_IN              : in  std_logic;
    GT9_TXCLK_LOCK_OUT           : out std_logic;
    GT9_TX_MMCM_RESET_IN         : in std_logic;
    GT9_RXUSRCLK_OUT             : out std_logic;
    GT9_RXUSRCLK2_OUT            : out std_logic;
    GT9_RXOUTCLK_IN              : in  std_logic;
    GT9_RXCLK_LOCK_OUT           : out std_logic;
    GT9_RX_MMCM_RESET_IN         : in std_logic;
 
    GT10_TXUSRCLK_OUT             : out std_logic;
    GT10_TXUSRCLK2_OUT            : out std_logic;
    GT10_TXOUTCLK_IN              : in  std_logic;
    GT10_TXCLK_LOCK_OUT           : out std_logic;
    GT10_TX_MMCM_RESET_IN         : in std_logic;
    GT10_RXUSRCLK_OUT             : out std_logic;
    GT10_RXUSRCLK2_OUT            : out std_logic;
    GT10_RXOUTCLK_IN              : in  std_logic;
    GT10_RXCLK_LOCK_OUT           : out std_logic;
    GT10_RX_MMCM_RESET_IN         : in std_logic;
 
    GT11_TXUSRCLK_OUT             : out std_logic;
    GT11_TXUSRCLK2_OUT            : out std_logic;
    GT11_TXOUTCLK_IN              : in  std_logic;
    GT11_TXCLK_LOCK_OUT           : out std_logic;
    GT11_TX_MMCM_RESET_IN         : in std_logic;
    GT11_RXUSRCLK_OUT             : out std_logic;
    GT11_RXUSRCLK2_OUT            : out std_logic;
    GT11_RXOUTCLK_IN              : in  std_logic;
    GT11_RXCLK_LOCK_OUT           : out std_logic;
    GT11_RX_MMCM_RESET_IN         : in std_logic;
 
    GT12_TXUSRCLK_OUT             : out std_logic;
    GT12_TXUSRCLK2_OUT            : out std_logic;
    GT12_TXOUTCLK_IN              : in  std_logic;
    GT12_TXCLK_LOCK_OUT           : out std_logic;
    GT12_TX_MMCM_RESET_IN         : in std_logic;
    GT12_RXUSRCLK_OUT             : out std_logic;
    GT12_RXUSRCLK2_OUT            : out std_logic;
    GT12_RXOUTCLK_IN              : in  std_logic;
    GT12_RXCLK_LOCK_OUT           : out std_logic;
    GT12_RX_MMCM_RESET_IN         : in std_logic;
 
    GT13_TXUSRCLK_OUT             : out std_logic;
    GT13_TXUSRCLK2_OUT            : out std_logic;
    GT13_TXOUTCLK_IN              : in  std_logic;
    GT13_TXCLK_LOCK_OUT           : out std_logic;
    GT13_TX_MMCM_RESET_IN         : in std_logic;
    GT13_RXUSRCLK_OUT             : out std_logic;
    GT13_RXUSRCLK2_OUT            : out std_logic;
    GT13_RXOUTCLK_IN              : in  std_logic;
    GT13_RXCLK_LOCK_OUT           : out std_logic;
    GT13_RX_MMCM_RESET_IN         : in std_logic;
 
    GT14_TXUSRCLK_OUT             : out std_logic;
    GT14_TXUSRCLK2_OUT            : out std_logic;
    GT14_TXOUTCLK_IN              : in  std_logic;
    GT14_TXCLK_LOCK_OUT           : out std_logic;
    GT14_TX_MMCM_RESET_IN         : in std_logic;
    GT14_RXUSRCLK_OUT             : out std_logic;
    GT14_RXUSRCLK2_OUT            : out std_logic;
    GT14_RXOUTCLK_IN              : in  std_logic;
    GT14_RXCLK_LOCK_OUT           : out std_logic;
    GT14_RX_MMCM_RESET_IN         : in std_logic;
 
    GT15_TXUSRCLK_OUT             : out std_logic;
    GT15_TXUSRCLK2_OUT            : out std_logic;
    GT15_TXOUTCLK_IN              : in  std_logic;
    GT15_TXCLK_LOCK_OUT           : out std_logic;
    GT15_TX_MMCM_RESET_IN         : in std_logic;
    GT15_RXUSRCLK_OUT             : out std_logic;
    GT15_RXUSRCLK2_OUT            : out std_logic;
    GT15_RXOUTCLK_IN              : in  std_logic;
    GT15_RXCLK_LOCK_OUT           : out std_logic;
    GT15_RX_MMCM_RESET_IN         : in std_logic;
 
    GT16_TXUSRCLK_OUT             : out std_logic;
    GT16_TXUSRCLK2_OUT            : out std_logic;
    GT16_TXOUTCLK_IN              : in  std_logic;
    GT16_TXCLK_LOCK_OUT           : out std_logic;
    GT16_TX_MMCM_RESET_IN         : in std_logic;
    GT16_RXUSRCLK_OUT             : out std_logic;
    GT16_RXUSRCLK2_OUT            : out std_logic;
    GT16_RXOUTCLK_IN              : in  std_logic;
    GT16_RXCLK_LOCK_OUT           : out std_logic;
    GT16_RX_MMCM_RESET_IN         : in std_logic;
 
    GT17_TXUSRCLK_OUT             : out std_logic;
    GT17_TXUSRCLK2_OUT            : out std_logic;
    GT17_TXOUTCLK_IN              : in  std_logic;
    GT17_TXCLK_LOCK_OUT           : out std_logic;
    GT17_TX_MMCM_RESET_IN         : in std_logic;
    GT17_RXUSRCLK_OUT             : out std_logic;
    GT17_RXUSRCLK2_OUT            : out std_logic;
    GT17_RXOUTCLK_IN              : in  std_logic;
    GT17_RXCLK_LOCK_OUT           : out std_logic;
    GT17_RX_MMCM_RESET_IN         : in std_logic;
 
    GT18_TXUSRCLK_OUT             : out std_logic;
    GT18_TXUSRCLK2_OUT            : out std_logic;
    GT18_TXOUTCLK_IN              : in  std_logic;
    GT18_TXCLK_LOCK_OUT           : out std_logic;
    GT18_TX_MMCM_RESET_IN         : in std_logic;
    GT18_RXUSRCLK_OUT             : out std_logic;
    GT18_RXUSRCLK2_OUT            : out std_logic;
    GT18_RXOUTCLK_IN              : in  std_logic;
    GT18_RXCLK_LOCK_OUT           : out std_logic;
    GT18_RX_MMCM_RESET_IN         : in std_logic;
 
    GT19_TXUSRCLK_OUT             : out std_logic;
    GT19_TXUSRCLK2_OUT            : out std_logic;
    GT19_TXOUTCLK_IN              : in  std_logic;
    GT19_TXCLK_LOCK_OUT           : out std_logic;
    GT19_TX_MMCM_RESET_IN         : in std_logic;
    GT19_RXUSRCLK_OUT             : out std_logic;
    GT19_RXUSRCLK2_OUT            : out std_logic;
    GT19_RXOUTCLK_IN              : in  std_logic;
    GT19_RXCLK_LOCK_OUT           : out std_logic;
    GT19_RX_MMCM_RESET_IN         : in std_logic;
 
    GT20_TXUSRCLK_OUT             : out std_logic;
    GT20_TXUSRCLK2_OUT            : out std_logic;
    GT20_TXOUTCLK_IN              : in  std_logic;
    GT20_TXCLK_LOCK_OUT           : out std_logic;
    GT20_TX_MMCM_RESET_IN         : in std_logic;
    GT20_RXUSRCLK_OUT             : out std_logic;
    GT20_RXUSRCLK2_OUT            : out std_logic;
    GT20_RXOUTCLK_IN              : in  std_logic;
    GT20_RXCLK_LOCK_OUT           : out std_logic;
    GT20_RX_MMCM_RESET_IN         : in std_logic;
 
    GT21_TXUSRCLK_OUT             : out std_logic;
    GT21_TXUSRCLK2_OUT            : out std_logic;
    GT21_TXOUTCLK_IN              : in  std_logic;
    GT21_TXCLK_LOCK_OUT           : out std_logic;
    GT21_TX_MMCM_RESET_IN         : in std_logic;
    GT21_RXUSRCLK_OUT             : out std_logic;
    GT21_RXUSRCLK2_OUT            : out std_logic;
    GT21_RXOUTCLK_IN              : in  std_logic;
    GT21_RXCLK_LOCK_OUT           : out std_logic;
    GT21_RX_MMCM_RESET_IN         : in std_logic;
 
    GT22_TXUSRCLK_OUT             : out std_logic;
    GT22_TXUSRCLK2_OUT            : out std_logic;
    GT22_TXOUTCLK_IN              : in  std_logic;
    GT22_TXCLK_LOCK_OUT           : out std_logic;
    GT22_TX_MMCM_RESET_IN         : in std_logic;
    GT22_RXUSRCLK_OUT             : out std_logic;
    GT22_RXUSRCLK2_OUT            : out std_logic;
    GT22_RXOUTCLK_IN              : in  std_logic;
    GT22_RXCLK_LOCK_OUT           : out std_logic;
    GT22_RX_MMCM_RESET_IN         : in std_logic;
 
    GT23_TXUSRCLK_OUT             : out std_logic;
    GT23_TXUSRCLK2_OUT            : out std_logic;
    GT23_TXOUTCLK_IN              : in  std_logic;
    GT23_TXCLK_LOCK_OUT           : out std_logic;
    GT23_TX_MMCM_RESET_IN         : in std_logic;
    GT23_RXUSRCLK_OUT             : out std_logic;
    GT23_RXUSRCLK2_OUT            : out std_logic;
    GT23_RXOUTCLK_IN              : in  std_logic;
    GT23_RXCLK_LOCK_OUT           : out std_logic;
    GT23_RX_MMCM_RESET_IN         : in std_logic;
 
    GT24_TXUSRCLK_OUT             : out std_logic;
    GT24_TXUSRCLK2_OUT            : out std_logic;
    GT24_TXOUTCLK_IN              : in  std_logic;
    GT24_TXCLK_LOCK_OUT           : out std_logic;
    GT24_TX_MMCM_RESET_IN         : in std_logic;
    GT24_RXUSRCLK_OUT             : out std_logic;
    GT24_RXUSRCLK2_OUT            : out std_logic;
    GT24_RXOUTCLK_IN              : in  std_logic;
    GT24_RXCLK_LOCK_OUT           : out std_logic;
    GT24_RX_MMCM_RESET_IN         : in std_logic;
 
    GT25_TXUSRCLK_OUT             : out std_logic;
    GT25_TXUSRCLK2_OUT            : out std_logic;
    GT25_TXOUTCLK_IN              : in  std_logic;
    GT25_TXCLK_LOCK_OUT           : out std_logic;
    GT25_TX_MMCM_RESET_IN         : in std_logic;
    GT25_RXUSRCLK_OUT             : out std_logic;
    GT25_RXUSRCLK2_OUT            : out std_logic;
    GT25_RXOUTCLK_IN              : in  std_logic;
    GT25_RXCLK_LOCK_OUT           : out std_logic;
    GT25_RX_MMCM_RESET_IN         : in std_logic;
 
    GT26_TXUSRCLK_OUT             : out std_logic;
    GT26_TXUSRCLK2_OUT            : out std_logic;
    GT26_TXOUTCLK_IN              : in  std_logic;
    GT26_TXCLK_LOCK_OUT           : out std_logic;
    GT26_TX_MMCM_RESET_IN         : in std_logic;
    GT26_RXUSRCLK_OUT             : out std_logic;
    GT26_RXUSRCLK2_OUT            : out std_logic;
    GT26_RXOUTCLK_IN              : in  std_logic;
    GT26_RXCLK_LOCK_OUT           : out std_logic;
    GT26_RX_MMCM_RESET_IN         : in std_logic;
 
    GT27_TXUSRCLK_OUT             : out std_logic;
    GT27_TXUSRCLK2_OUT            : out std_logic;
    GT27_TXOUTCLK_IN              : in  std_logic;
    GT27_TXCLK_LOCK_OUT           : out std_logic;
    GT27_TX_MMCM_RESET_IN         : in std_logic;
    GT27_RXUSRCLK_OUT             : out std_logic;
    GT27_RXUSRCLK2_OUT            : out std_logic;
    GT27_RXOUTCLK_IN              : in  std_logic;
    GT27_RXCLK_LOCK_OUT           : out std_logic;
    GT27_RX_MMCM_RESET_IN         : in std_logic;
 
    GT28_TXUSRCLK_OUT             : out std_logic;
    GT28_TXUSRCLK2_OUT            : out std_logic;
    GT28_TXOUTCLK_IN              : in  std_logic;
    GT28_TXCLK_LOCK_OUT           : out std_logic;
    GT28_TX_MMCM_RESET_IN         : in std_logic;
    GT28_RXUSRCLK_OUT             : out std_logic;
    GT28_RXUSRCLK2_OUT            : out std_logic;
    GT28_RXOUTCLK_IN              : in  std_logic;
    GT28_RXCLK_LOCK_OUT           : out std_logic;
    GT28_RX_MMCM_RESET_IN         : in std_logic;
 
    GT29_TXUSRCLK_OUT             : out std_logic;
    GT29_TXUSRCLK2_OUT            : out std_logic;
    GT29_TXOUTCLK_IN              : in  std_logic;
    GT29_TXCLK_LOCK_OUT           : out std_logic;
    GT29_TX_MMCM_RESET_IN         : in std_logic;
    GT29_RXUSRCLK_OUT             : out std_logic;
    GT29_RXUSRCLK2_OUT            : out std_logic;
    GT29_RXOUTCLK_IN              : in  std_logic;
    GT29_RXCLK_LOCK_OUT           : out std_logic;
    GT29_RX_MMCM_RESET_IN         : in std_logic;
 
    GT30_TXUSRCLK_OUT             : out std_logic;
    GT30_TXUSRCLK2_OUT            : out std_logic;
    GT30_TXOUTCLK_IN              : in  std_logic;
    GT30_TXCLK_LOCK_OUT           : out std_logic;
    GT30_TX_MMCM_RESET_IN         : in std_logic;
    GT30_RXUSRCLK_OUT             : out std_logic;
    GT30_RXUSRCLK2_OUT            : out std_logic;
    GT30_RXOUTCLK_IN              : in  std_logic;
    GT30_RXCLK_LOCK_OUT           : out std_logic;
    GT30_RX_MMCM_RESET_IN         : in std_logic;
 
    GT31_TXUSRCLK_OUT             : out std_logic;
    GT31_TXUSRCLK2_OUT            : out std_logic;
    GT31_TXOUTCLK_IN              : in  std_logic;
    GT31_TXCLK_LOCK_OUT           : out std_logic;
    GT31_TX_MMCM_RESET_IN         : in std_logic;
    GT31_RXUSRCLK_OUT             : out std_logic;
    GT31_RXUSRCLK2_OUT            : out std_logic;
    GT31_RXOUTCLK_IN              : in  std_logic;
    GT31_RXCLK_LOCK_OUT           : out std_logic;
    GT31_RX_MMCM_RESET_IN         : in std_logic;
    Q2_CLK0_GTREFCLK_PAD_N_IN               : in   std_logic;
    Q2_CLK0_GTREFCLK_PAD_P_IN               : in   std_logic;
    Q2_CLK0_GTREFCLK_OUT                    : out  std_logic;
    Q5_CLK0_GTREFCLK_PAD_N_IN               : in   std_logic;
    Q5_CLK0_GTREFCLK_PAD_P_IN               : in   std_logic;
    Q5_CLK0_GTREFCLK_OUT                    : out  std_logic;
    Q7_CLK0_GTREFCLK_PAD_N_IN               : in   std_logic;
    Q7_CLK0_GTREFCLK_PAD_P_IN               : in   std_logic;
    Q7_CLK0_GTREFCLK_OUT                    : out  std_logic
);
end component;

--***********************************Parameter Declarations********************

    constant DLY : time := 1 ns;

--************************** Register Declarations ****************************

    signal   gt0_txfsmresetdone_i            : std_logic;
signal   gt0_rxfsmresetdone_i            : std_logic;
    signal   gt0_txfsmresetdone_r            : std_logic;
    signal   gt0_txfsmresetdone_r2           : std_logic;
signal   gt0_rxresetdone_r               : std_logic;
signal   gt0_rxresetdone_r2              : std_logic;
signal   gt0_rxresetdone_r3              : std_logic;


    signal   gt1_txfsmresetdone_i            : std_logic;
signal   gt1_rxfsmresetdone_i            : std_logic;
    signal   gt1_txfsmresetdone_r            : std_logic;
    signal   gt1_txfsmresetdone_r2           : std_logic;
signal   gt1_rxresetdone_r               : std_logic;
signal   gt1_rxresetdone_r2              : std_logic;
signal   gt1_rxresetdone_r3              : std_logic;


    signal   gt2_txfsmresetdone_i            : std_logic;
signal   gt2_rxfsmresetdone_i            : std_logic;
    signal   gt2_txfsmresetdone_r            : std_logic;
    signal   gt2_txfsmresetdone_r2           : std_logic;
signal   gt2_rxresetdone_r               : std_logic;
signal   gt2_rxresetdone_r2              : std_logic;
signal   gt2_rxresetdone_r3              : std_logic;


    signal   gt3_txfsmresetdone_i            : std_logic;
signal   gt3_rxfsmresetdone_i            : std_logic;
    signal   gt3_txfsmresetdone_r            : std_logic;
    signal   gt3_txfsmresetdone_r2           : std_logic;
signal   gt3_rxresetdone_r               : std_logic;
signal   gt3_rxresetdone_r2              : std_logic;
signal   gt3_rxresetdone_r3              : std_logic;


    signal   gt4_txfsmresetdone_i            : std_logic;
signal   gt4_rxfsmresetdone_i            : std_logic;
    signal   gt4_txfsmresetdone_r            : std_logic;
    signal   gt4_txfsmresetdone_r2           : std_logic;
signal   gt4_rxresetdone_r               : std_logic;
signal   gt4_rxresetdone_r2              : std_logic;
signal   gt4_rxresetdone_r3              : std_logic;


    signal   gt5_txfsmresetdone_i            : std_logic;
signal   gt5_rxfsmresetdone_i            : std_logic;
    signal   gt5_txfsmresetdone_r            : std_logic;
    signal   gt5_txfsmresetdone_r2           : std_logic;
signal   gt5_rxresetdone_r               : std_logic;
signal   gt5_rxresetdone_r2              : std_logic;
signal   gt5_rxresetdone_r3              : std_logic;


    signal   gt6_txfsmresetdone_i            : std_logic;
signal   gt6_rxfsmresetdone_i            : std_logic;
    signal   gt6_txfsmresetdone_r            : std_logic;
    signal   gt6_txfsmresetdone_r2           : std_logic;
signal   gt6_rxresetdone_r               : std_logic;
signal   gt6_rxresetdone_r2              : std_logic;
signal   gt6_rxresetdone_r3              : std_logic;


    signal   gt7_txfsmresetdone_i            : std_logic;
signal   gt7_rxfsmresetdone_i            : std_logic;
    signal   gt7_txfsmresetdone_r            : std_logic;
    signal   gt7_txfsmresetdone_r2           : std_logic;
signal   gt7_rxresetdone_r               : std_logic;
signal   gt7_rxresetdone_r2              : std_logic;
signal   gt7_rxresetdone_r3              : std_logic;


    signal   gt8_txfsmresetdone_i            : std_logic;
signal   gt8_rxfsmresetdone_i            : std_logic;
    signal   gt8_txfsmresetdone_r            : std_logic;
    signal   gt8_txfsmresetdone_r2           : std_logic;
signal   gt8_rxresetdone_r               : std_logic;
signal   gt8_rxresetdone_r2              : std_logic;
signal   gt8_rxresetdone_r3              : std_logic;


    signal   gt9_txfsmresetdone_i            : std_logic;
signal   gt9_rxfsmresetdone_i            : std_logic;
    signal   gt9_txfsmresetdone_r            : std_logic;
    signal   gt9_txfsmresetdone_r2           : std_logic;
signal   gt9_rxresetdone_r               : std_logic;
signal   gt9_rxresetdone_r2              : std_logic;
signal   gt9_rxresetdone_r3              : std_logic;


    signal   gt10_txfsmresetdone_i           : std_logic;
signal   gt10_rxfsmresetdone_i           : std_logic;
    signal   gt10_txfsmresetdone_r           : std_logic;
    signal   gt10_txfsmresetdone_r2          : std_logic;
signal   gt10_rxresetdone_r              : std_logic;
signal   gt10_rxresetdone_r2             : std_logic;
signal   gt10_rxresetdone_r3             : std_logic;


    signal   gt11_txfsmresetdone_i           : std_logic;
signal   gt11_rxfsmresetdone_i           : std_logic;
    signal   gt11_txfsmresetdone_r           : std_logic;
    signal   gt11_txfsmresetdone_r2          : std_logic;
signal   gt11_rxresetdone_r              : std_logic;
signal   gt11_rxresetdone_r2             : std_logic;
signal   gt11_rxresetdone_r3             : std_logic;


    signal   gt12_txfsmresetdone_i           : std_logic;
signal   gt12_rxfsmresetdone_i           : std_logic;
    signal   gt12_txfsmresetdone_r           : std_logic;
    signal   gt12_txfsmresetdone_r2          : std_logic;
signal   gt12_rxresetdone_r              : std_logic;
signal   gt12_rxresetdone_r2             : std_logic;
signal   gt12_rxresetdone_r3             : std_logic;


    signal   gt13_txfsmresetdone_i           : std_logic;
signal   gt13_rxfsmresetdone_i           : std_logic;
    signal   gt13_txfsmresetdone_r           : std_logic;
    signal   gt13_txfsmresetdone_r2          : std_logic;
signal   gt13_rxresetdone_r              : std_logic;
signal   gt13_rxresetdone_r2             : std_logic;
signal   gt13_rxresetdone_r3             : std_logic;


    signal   gt14_txfsmresetdone_i           : std_logic;
signal   gt14_rxfsmresetdone_i           : std_logic;
    signal   gt14_txfsmresetdone_r           : std_logic;
    signal   gt14_txfsmresetdone_r2          : std_logic;
signal   gt14_rxresetdone_r              : std_logic;
signal   gt14_rxresetdone_r2             : std_logic;
signal   gt14_rxresetdone_r3             : std_logic;


    signal   gt15_txfsmresetdone_i           : std_logic;
signal   gt15_rxfsmresetdone_i           : std_logic;
    signal   gt15_txfsmresetdone_r           : std_logic;
    signal   gt15_txfsmresetdone_r2          : std_logic;
signal   gt15_rxresetdone_r              : std_logic;
signal   gt15_rxresetdone_r2             : std_logic;
signal   gt15_rxresetdone_r3             : std_logic;


    signal   gt16_txfsmresetdone_i           : std_logic;
signal   gt16_rxfsmresetdone_i           : std_logic;
    signal   gt16_txfsmresetdone_r           : std_logic;
    signal   gt16_txfsmresetdone_r2          : std_logic;
signal   gt16_rxresetdone_r              : std_logic;
signal   gt16_rxresetdone_r2             : std_logic;
signal   gt16_rxresetdone_r3             : std_logic;


    signal   gt17_txfsmresetdone_i           : std_logic;
signal   gt17_rxfsmresetdone_i           : std_logic;
    signal   gt17_txfsmresetdone_r           : std_logic;
    signal   gt17_txfsmresetdone_r2          : std_logic;
signal   gt17_rxresetdone_r              : std_logic;
signal   gt17_rxresetdone_r2             : std_logic;
signal   gt17_rxresetdone_r3             : std_logic;


    signal   gt18_txfsmresetdone_i           : std_logic;
signal   gt18_rxfsmresetdone_i           : std_logic;
    signal   gt18_txfsmresetdone_r           : std_logic;
    signal   gt18_txfsmresetdone_r2          : std_logic;
signal   gt18_rxresetdone_r              : std_logic;
signal   gt18_rxresetdone_r2             : std_logic;
signal   gt18_rxresetdone_r3             : std_logic;


    signal   gt19_txfsmresetdone_i           : std_logic;
signal   gt19_rxfsmresetdone_i           : std_logic;
    signal   gt19_txfsmresetdone_r           : std_logic;
    signal   gt19_txfsmresetdone_r2          : std_logic;
signal   gt19_rxresetdone_r              : std_logic;
signal   gt19_rxresetdone_r2             : std_logic;
signal   gt19_rxresetdone_r3             : std_logic;


    signal   gt20_txfsmresetdone_i           : std_logic;
signal   gt20_rxfsmresetdone_i           : std_logic;
    signal   gt20_txfsmresetdone_r           : std_logic;
    signal   gt20_txfsmresetdone_r2          : std_logic;
signal   gt20_rxresetdone_r              : std_logic;
signal   gt20_rxresetdone_r2             : std_logic;
signal   gt20_rxresetdone_r3             : std_logic;


    signal   gt21_txfsmresetdone_i           : std_logic;
signal   gt21_rxfsmresetdone_i           : std_logic;
    signal   gt21_txfsmresetdone_r           : std_logic;
    signal   gt21_txfsmresetdone_r2          : std_logic;
signal   gt21_rxresetdone_r              : std_logic;
signal   gt21_rxresetdone_r2             : std_logic;
signal   gt21_rxresetdone_r3             : std_logic;


    signal   gt22_txfsmresetdone_i           : std_logic;
signal   gt22_rxfsmresetdone_i           : std_logic;
    signal   gt22_txfsmresetdone_r           : std_logic;
    signal   gt22_txfsmresetdone_r2          : std_logic;
signal   gt22_rxresetdone_r              : std_logic;
signal   gt22_rxresetdone_r2             : std_logic;
signal   gt22_rxresetdone_r3             : std_logic;


    signal   gt23_txfsmresetdone_i           : std_logic;
signal   gt23_rxfsmresetdone_i           : std_logic;
    signal   gt23_txfsmresetdone_r           : std_logic;
    signal   gt23_txfsmresetdone_r2          : std_logic;
signal   gt23_rxresetdone_r              : std_logic;
signal   gt23_rxresetdone_r2             : std_logic;
signal   gt23_rxresetdone_r3             : std_logic;


    signal   gt24_txfsmresetdone_i           : std_logic;
signal   gt24_rxfsmresetdone_i           : std_logic;
    signal   gt24_txfsmresetdone_r           : std_logic;
    signal   gt24_txfsmresetdone_r2          : std_logic;
signal   gt24_rxresetdone_r              : std_logic;
signal   gt24_rxresetdone_r2             : std_logic;
signal   gt24_rxresetdone_r3             : std_logic;


    signal   gt25_txfsmresetdone_i           : std_logic;
signal   gt25_rxfsmresetdone_i           : std_logic;
    signal   gt25_txfsmresetdone_r           : std_logic;
    signal   gt25_txfsmresetdone_r2          : std_logic;
signal   gt25_rxresetdone_r              : std_logic;
signal   gt25_rxresetdone_r2             : std_logic;
signal   gt25_rxresetdone_r3             : std_logic;


    signal   gt26_txfsmresetdone_i           : std_logic;
signal   gt26_rxfsmresetdone_i           : std_logic;
    signal   gt26_txfsmresetdone_r           : std_logic;
    signal   gt26_txfsmresetdone_r2          : std_logic;
signal   gt26_rxresetdone_r              : std_logic;
signal   gt26_rxresetdone_r2             : std_logic;
signal   gt26_rxresetdone_r3             : std_logic;


    signal   gt27_txfsmresetdone_i           : std_logic;
signal   gt27_rxfsmresetdone_i           : std_logic;
    signal   gt27_txfsmresetdone_r           : std_logic;
    signal   gt27_txfsmresetdone_r2          : std_logic;
signal   gt27_rxresetdone_r              : std_logic;
signal   gt27_rxresetdone_r2             : std_logic;
signal   gt27_rxresetdone_r3             : std_logic;


    signal   gt28_txfsmresetdone_i           : std_logic;
signal   gt28_rxfsmresetdone_i           : std_logic;
    signal   gt28_txfsmresetdone_r           : std_logic;
    signal   gt28_txfsmresetdone_r2          : std_logic;
signal   gt28_rxresetdone_r              : std_logic;
signal   gt28_rxresetdone_r2             : std_logic;
signal   gt28_rxresetdone_r3             : std_logic;


    signal   gt29_txfsmresetdone_i           : std_logic;
signal   gt29_rxfsmresetdone_i           : std_logic;
    signal   gt29_txfsmresetdone_r           : std_logic;
    signal   gt29_txfsmresetdone_r2          : std_logic;
signal   gt29_rxresetdone_r              : std_logic;
signal   gt29_rxresetdone_r2             : std_logic;
signal   gt29_rxresetdone_r3             : std_logic;


    signal   gt30_txfsmresetdone_i           : std_logic;
signal   gt30_rxfsmresetdone_i           : std_logic;
    signal   gt30_txfsmresetdone_r           : std_logic;
    signal   gt30_txfsmresetdone_r2          : std_logic;
signal   gt30_rxresetdone_r              : std_logic;
signal   gt30_rxresetdone_r2             : std_logic;
signal   gt30_rxresetdone_r3             : std_logic;


    signal   gt31_txfsmresetdone_i           : std_logic;
signal   gt31_rxfsmresetdone_i           : std_logic;
    signal   gt31_txfsmresetdone_r           : std_logic;
    signal   gt31_txfsmresetdone_r2          : std_logic;
signal   gt31_rxresetdone_r              : std_logic;
signal   gt31_rxresetdone_r2             : std_logic;
signal   gt31_rxresetdone_r3             : std_logic;


signal   reset_pulse                     : std_logic_vector(3 downto 0);
    signal   reset_counter  :   unsigned(5 downto 0) := "000000";

--**************************** Wire Declarations ******************************
    -------------------------- GT Wrapper Wires ------------------------------
    --________________________________________________________________________
    --________________________________________________________________________
    --GT0  (X1Y4)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt0_drpaddr_i                   : std_logic_vector(8 downto 0);
    signal  gt0_drpdi_i                     : std_logic_vector(15 downto 0);
    signal  gt0_drpdo_i                     : std_logic_vector(15 downto 0);
    signal  gt0_drpen_i                     : std_logic;
    signal  gt0_drprdy_i                    : std_logic;
    signal  gt0_drpwe_i                     : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt0_eyescanreset_i              : std_logic;
    signal  gt0_rxuserrdy_i                 : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt0_eyescandataerror_i          : std_logic;
    signal  gt0_eyescantrigger_i            : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt0_rxslide_i                   : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt0_dmonitorout_i               : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt0_rxdata_i                    : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt0_rxdisperr_i                 : std_logic_vector(7 downto 0);
    signal  gt0_rxnotintable_i              : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt0_gthrxn_i                    : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt0_rxdlyen_i                   : std_logic;
    signal  gt0_rxdlysreset_i               : std_logic;
    signal  gt0_rxdlysresetdone_i           : std_logic;
    signal  gt0_rxphalign_i                 : std_logic;
    signal  gt0_rxphaligndone_i             : std_logic;
    signal  gt0_rxphalignen_i               : std_logic;
    signal  gt0_rxphdlyreset_i              : std_logic;
    signal  gt0_rxphmonitor_i               : std_logic_vector(4 downto 0);
    signal  gt0_rxphslipmonitor_i           : std_logic_vector(4 downto 0);
    signal  gt0_rxsyncallin_i               : std_logic;
    signal  gt0_rxsyncdone_i                : std_logic;
    signal  gt0_rxsyncin_i                  : std_logic;
    signal  gt0_rxsyncmode_i                : std_logic;
    signal  gt0_rxsyncout_i                 : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt0_rxbyteisaligned_i           : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt0_rxlpmhfhold_i               : std_logic;
    signal  gt0_rxlpmlfhold_i               : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt0_rxmonitorout_i              : std_logic_vector(6 downto 0);
    signal  gt0_rxmonitorsel_i              : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt0_rxoutclk_i                  : std_logic;
    signal  gt0_rxoutclkfabric_i            : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt0_gtrxreset_i                 : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt0_rxcharisk_i                 : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt0_gthrxp_i                    : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt0_rxresetdone_i               : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt0_gttxreset_i                 : std_logic;
    signal  gt0_txuserrdy_i                 : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt0_txdlyen_i                   : std_logic;
    signal  gt0_txdlysreset_i               : std_logic;
    signal  gt0_txdlysresetdone_i           : std_logic;
    signal  gt0_txphalign_i                 : std_logic;
    signal  gt0_txphaligndone_i             : std_logic;
    signal  gt0_txphalignen_i               : std_logic;
    signal  gt0_txphdlyreset_i              : std_logic;
    signal  gt0_txphinit_i                  : std_logic;
    signal  gt0_txphinitdone_i              : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt0_txdata_i                    : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt0_gthtxn_i                    : std_logic;
    signal  gt0_gthtxp_i                    : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt0_txoutclk_i                  : std_logic;
    signal  gt0_txoutclkfabric_i            : std_logic;
    signal  gt0_txoutclkpcs_i               : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt0_txresetdone_i               : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt0_txcharisk_i                 : std_logic_vector(7 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT1  (X1Y5)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt1_drpaddr_i                   : std_logic_vector(8 downto 0);
    signal  gt1_drpdi_i                     : std_logic_vector(15 downto 0);
    signal  gt1_drpdo_i                     : std_logic_vector(15 downto 0);
    signal  gt1_drpen_i                     : std_logic;
    signal  gt1_drprdy_i                    : std_logic;
    signal  gt1_drpwe_i                     : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt1_eyescanreset_i              : std_logic;
    signal  gt1_rxuserrdy_i                 : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt1_eyescandataerror_i          : std_logic;
    signal  gt1_eyescantrigger_i            : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt1_rxslide_i                   : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt1_dmonitorout_i               : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt1_rxdata_i                    : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt1_rxdisperr_i                 : std_logic_vector(7 downto 0);
    signal  gt1_rxnotintable_i              : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt1_gthrxn_i                    : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt1_rxdlyen_i                   : std_logic;
    signal  gt1_rxdlysreset_i               : std_logic;
    signal  gt1_rxdlysresetdone_i           : std_logic;
    signal  gt1_rxphalign_i                 : std_logic;
    signal  gt1_rxphaligndone_i             : std_logic;
    signal  gt1_rxphalignen_i               : std_logic;
    signal  gt1_rxphdlyreset_i              : std_logic;
    signal  gt1_rxphmonitor_i               : std_logic_vector(4 downto 0);
    signal  gt1_rxphslipmonitor_i           : std_logic_vector(4 downto 0);
    signal  gt1_rxsyncallin_i               : std_logic;
    signal  gt1_rxsyncdone_i                : std_logic;
    signal  gt1_rxsyncin_i                  : std_logic;
    signal  gt1_rxsyncmode_i                : std_logic;
    signal  gt1_rxsyncout_i                 : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt1_rxbyteisaligned_i           : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt1_rxlpmhfhold_i               : std_logic;
    signal  gt1_rxlpmlfhold_i               : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt1_rxmonitorout_i              : std_logic_vector(6 downto 0);
    signal  gt1_rxmonitorsel_i              : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt1_rxoutclk_i                  : std_logic;
    signal  gt1_rxoutclkfabric_i            : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt1_gtrxreset_i                 : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt1_rxcharisk_i                 : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt1_gthrxp_i                    : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt1_rxresetdone_i               : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt1_gttxreset_i                 : std_logic;
    signal  gt1_txuserrdy_i                 : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt1_txdlyen_i                   : std_logic;
    signal  gt1_txdlysreset_i               : std_logic;
    signal  gt1_txdlysresetdone_i           : std_logic;
    signal  gt1_txphalign_i                 : std_logic;
    signal  gt1_txphaligndone_i             : std_logic;
    signal  gt1_txphalignen_i               : std_logic;
    signal  gt1_txphdlyreset_i              : std_logic;
    signal  gt1_txphinit_i                  : std_logic;
    signal  gt1_txphinitdone_i              : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt1_txdata_i                    : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt1_gthtxn_i                    : std_logic;
    signal  gt1_gthtxp_i                    : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt1_txoutclk_i                  : std_logic;
    signal  gt1_txoutclkfabric_i            : std_logic;
    signal  gt1_txoutclkpcs_i               : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt1_txresetdone_i               : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt1_txcharisk_i                 : std_logic_vector(7 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT2  (X1Y6)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt2_drpaddr_i                   : std_logic_vector(8 downto 0);
    signal  gt2_drpdi_i                     : std_logic_vector(15 downto 0);
    signal  gt2_drpdo_i                     : std_logic_vector(15 downto 0);
    signal  gt2_drpen_i                     : std_logic;
    signal  gt2_drprdy_i                    : std_logic;
    signal  gt2_drpwe_i                     : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt2_eyescanreset_i              : std_logic;
    signal  gt2_rxuserrdy_i                 : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt2_eyescandataerror_i          : std_logic;
    signal  gt2_eyescantrigger_i            : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt2_rxslide_i                   : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt2_dmonitorout_i               : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt2_rxdata_i                    : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt2_rxdisperr_i                 : std_logic_vector(7 downto 0);
    signal  gt2_rxnotintable_i              : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt2_gthrxn_i                    : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt2_rxdlyen_i                   : std_logic;
    signal  gt2_rxdlysreset_i               : std_logic;
    signal  gt2_rxdlysresetdone_i           : std_logic;
    signal  gt2_rxphalign_i                 : std_logic;
    signal  gt2_rxphaligndone_i             : std_logic;
    signal  gt2_rxphalignen_i               : std_logic;
    signal  gt2_rxphdlyreset_i              : std_logic;
    signal  gt2_rxphmonitor_i               : std_logic_vector(4 downto 0);
    signal  gt2_rxphslipmonitor_i           : std_logic_vector(4 downto 0);
    signal  gt2_rxsyncallin_i               : std_logic;
    signal  gt2_rxsyncdone_i                : std_logic;
    signal  gt2_rxsyncin_i                  : std_logic;
    signal  gt2_rxsyncmode_i                : std_logic;
    signal  gt2_rxsyncout_i                 : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt2_rxbyteisaligned_i           : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt2_rxlpmhfhold_i               : std_logic;
    signal  gt2_rxlpmlfhold_i               : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt2_rxmonitorout_i              : std_logic_vector(6 downto 0);
    signal  gt2_rxmonitorsel_i              : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt2_rxoutclk_i                  : std_logic;
    signal  gt2_rxoutclkfabric_i            : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt2_gtrxreset_i                 : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt2_rxcharisk_i                 : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt2_gthrxp_i                    : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt2_rxresetdone_i               : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt2_gttxreset_i                 : std_logic;
    signal  gt2_txuserrdy_i                 : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt2_txdlyen_i                   : std_logic;
    signal  gt2_txdlysreset_i               : std_logic;
    signal  gt2_txdlysresetdone_i           : std_logic;
    signal  gt2_txphalign_i                 : std_logic;
    signal  gt2_txphaligndone_i             : std_logic;
    signal  gt2_txphalignen_i               : std_logic;
    signal  gt2_txphdlyreset_i              : std_logic;
    signal  gt2_txphinit_i                  : std_logic;
    signal  gt2_txphinitdone_i              : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt2_txdata_i                    : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt2_gthtxn_i                    : std_logic;
    signal  gt2_gthtxp_i                    : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt2_txoutclk_i                  : std_logic;
    signal  gt2_txoutclkfabric_i            : std_logic;
    signal  gt2_txoutclkpcs_i               : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt2_txresetdone_i               : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt2_txcharisk_i                 : std_logic_vector(7 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT3  (X1Y7)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt3_drpaddr_i                   : std_logic_vector(8 downto 0);
    signal  gt3_drpdi_i                     : std_logic_vector(15 downto 0);
    signal  gt3_drpdo_i                     : std_logic_vector(15 downto 0);
    signal  gt3_drpen_i                     : std_logic;
    signal  gt3_drprdy_i                    : std_logic;
    signal  gt3_drpwe_i                     : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt3_eyescanreset_i              : std_logic;
    signal  gt3_rxuserrdy_i                 : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt3_eyescandataerror_i          : std_logic;
    signal  gt3_eyescantrigger_i            : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt3_rxslide_i                   : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt3_dmonitorout_i               : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt3_rxdata_i                    : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt3_rxdisperr_i                 : std_logic_vector(7 downto 0);
    signal  gt3_rxnotintable_i              : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt3_gthrxn_i                    : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt3_rxdlyen_i                   : std_logic;
    signal  gt3_rxdlysreset_i               : std_logic;
    signal  gt3_rxdlysresetdone_i           : std_logic;
    signal  gt3_rxphalign_i                 : std_logic;
    signal  gt3_rxphaligndone_i             : std_logic;
    signal  gt3_rxphalignen_i               : std_logic;
    signal  gt3_rxphdlyreset_i              : std_logic;
    signal  gt3_rxphmonitor_i               : std_logic_vector(4 downto 0);
    signal  gt3_rxphslipmonitor_i           : std_logic_vector(4 downto 0);
    signal  gt3_rxsyncallin_i               : std_logic;
    signal  gt3_rxsyncdone_i                : std_logic;
    signal  gt3_rxsyncin_i                  : std_logic;
    signal  gt3_rxsyncmode_i                : std_logic;
    signal  gt3_rxsyncout_i                 : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt3_rxbyteisaligned_i           : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt3_rxlpmhfhold_i               : std_logic;
    signal  gt3_rxlpmlfhold_i               : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt3_rxmonitorout_i              : std_logic_vector(6 downto 0);
    signal  gt3_rxmonitorsel_i              : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt3_rxoutclk_i                  : std_logic;
    signal  gt3_rxoutclkfabric_i            : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt3_gtrxreset_i                 : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt3_rxcharisk_i                 : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt3_gthrxp_i                    : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt3_rxresetdone_i               : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt3_gttxreset_i                 : std_logic;
    signal  gt3_txuserrdy_i                 : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt3_txdlyen_i                   : std_logic;
    signal  gt3_txdlysreset_i               : std_logic;
    signal  gt3_txdlysresetdone_i           : std_logic;
    signal  gt3_txphalign_i                 : std_logic;
    signal  gt3_txphaligndone_i             : std_logic;
    signal  gt3_txphalignen_i               : std_logic;
    signal  gt3_txphdlyreset_i              : std_logic;
    signal  gt3_txphinit_i                  : std_logic;
    signal  gt3_txphinitdone_i              : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt3_txdata_i                    : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt3_gthtxn_i                    : std_logic;
    signal  gt3_gthtxp_i                    : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt3_txoutclk_i                  : std_logic;
    signal  gt3_txoutclkfabric_i            : std_logic;
    signal  gt3_txoutclkpcs_i               : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt3_txresetdone_i               : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt3_txcharisk_i                 : std_logic_vector(7 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT4  (X1Y8)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt4_drpaddr_i                   : std_logic_vector(8 downto 0);
    signal  gt4_drpdi_i                     : std_logic_vector(15 downto 0);
    signal  gt4_drpdo_i                     : std_logic_vector(15 downto 0);
    signal  gt4_drpen_i                     : std_logic;
    signal  gt4_drprdy_i                    : std_logic;
    signal  gt4_drpwe_i                     : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt4_eyescanreset_i              : std_logic;
    signal  gt4_rxuserrdy_i                 : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt4_eyescandataerror_i          : std_logic;
    signal  gt4_eyescantrigger_i            : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt4_rxslide_i                   : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt4_dmonitorout_i               : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt4_rxdata_i                    : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt4_rxdisperr_i                 : std_logic_vector(7 downto 0);
    signal  gt4_rxnotintable_i              : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt4_gthrxn_i                    : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt4_rxdlyen_i                   : std_logic;
    signal  gt4_rxdlysreset_i               : std_logic;
    signal  gt4_rxdlysresetdone_i           : std_logic;
    signal  gt4_rxphalign_i                 : std_logic;
    signal  gt4_rxphaligndone_i             : std_logic;
    signal  gt4_rxphalignen_i               : std_logic;
    signal  gt4_rxphdlyreset_i              : std_logic;
    signal  gt4_rxphmonitor_i               : std_logic_vector(4 downto 0);
    signal  gt4_rxphslipmonitor_i           : std_logic_vector(4 downto 0);
    signal  gt4_rxsyncallin_i               : std_logic;
    signal  gt4_rxsyncdone_i                : std_logic;
    signal  gt4_rxsyncin_i                  : std_logic;
    signal  gt4_rxsyncmode_i                : std_logic;
    signal  gt4_rxsyncout_i                 : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt4_rxbyteisaligned_i           : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt4_rxlpmhfhold_i               : std_logic;
    signal  gt4_rxlpmlfhold_i               : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt4_rxmonitorout_i              : std_logic_vector(6 downto 0);
    signal  gt4_rxmonitorsel_i              : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt4_rxoutclk_i                  : std_logic;
    signal  gt4_rxoutclkfabric_i            : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt4_gtrxreset_i                 : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt4_rxcharisk_i                 : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt4_gthrxp_i                    : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt4_rxresetdone_i               : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt4_gttxreset_i                 : std_logic;
    signal  gt4_txuserrdy_i                 : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt4_txdlyen_i                   : std_logic;
    signal  gt4_txdlysreset_i               : std_logic;
    signal  gt4_txdlysresetdone_i           : std_logic;
    signal  gt4_txphalign_i                 : std_logic;
    signal  gt4_txphaligndone_i             : std_logic;
    signal  gt4_txphalignen_i               : std_logic;
    signal  gt4_txphdlyreset_i              : std_logic;
    signal  gt4_txphinit_i                  : std_logic;
    signal  gt4_txphinitdone_i              : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt4_txdata_i                    : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt4_gthtxn_i                    : std_logic;
    signal  gt4_gthtxp_i                    : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt4_txoutclk_i                  : std_logic;
    signal  gt4_txoutclkfabric_i            : std_logic;
    signal  gt4_txoutclkpcs_i               : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt4_txresetdone_i               : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt4_txcharisk_i                 : std_logic_vector(7 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT5  (X1Y9)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt5_drpaddr_i                   : std_logic_vector(8 downto 0);
    signal  gt5_drpdi_i                     : std_logic_vector(15 downto 0);
    signal  gt5_drpdo_i                     : std_logic_vector(15 downto 0);
    signal  gt5_drpen_i                     : std_logic;
    signal  gt5_drprdy_i                    : std_logic;
    signal  gt5_drpwe_i                     : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt5_eyescanreset_i              : std_logic;
    signal  gt5_rxuserrdy_i                 : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt5_eyescandataerror_i          : std_logic;
    signal  gt5_eyescantrigger_i            : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt5_rxslide_i                   : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt5_dmonitorout_i               : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt5_rxdata_i                    : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt5_rxdisperr_i                 : std_logic_vector(7 downto 0);
    signal  gt5_rxnotintable_i              : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt5_gthrxn_i                    : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt5_rxdlyen_i                   : std_logic;
    signal  gt5_rxdlysreset_i               : std_logic;
    signal  gt5_rxdlysresetdone_i           : std_logic;
    signal  gt5_rxphalign_i                 : std_logic;
    signal  gt5_rxphaligndone_i             : std_logic;
    signal  gt5_rxphalignen_i               : std_logic;
    signal  gt5_rxphdlyreset_i              : std_logic;
    signal  gt5_rxphmonitor_i               : std_logic_vector(4 downto 0);
    signal  gt5_rxphslipmonitor_i           : std_logic_vector(4 downto 0);
    signal  gt5_rxsyncallin_i               : std_logic;
    signal  gt5_rxsyncdone_i                : std_logic;
    signal  gt5_rxsyncin_i                  : std_logic;
    signal  gt5_rxsyncmode_i                : std_logic;
    signal  gt5_rxsyncout_i                 : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt5_rxbyteisaligned_i           : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt5_rxlpmhfhold_i               : std_logic;
    signal  gt5_rxlpmlfhold_i               : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt5_rxmonitorout_i              : std_logic_vector(6 downto 0);
    signal  gt5_rxmonitorsel_i              : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt5_rxoutclk_i                  : std_logic;
    signal  gt5_rxoutclkfabric_i            : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt5_gtrxreset_i                 : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt5_rxcharisk_i                 : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt5_gthrxp_i                    : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt5_rxresetdone_i               : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt5_gttxreset_i                 : std_logic;
    signal  gt5_txuserrdy_i                 : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt5_txdlyen_i                   : std_logic;
    signal  gt5_txdlysreset_i               : std_logic;
    signal  gt5_txdlysresetdone_i           : std_logic;
    signal  gt5_txphalign_i                 : std_logic;
    signal  gt5_txphaligndone_i             : std_logic;
    signal  gt5_txphalignen_i               : std_logic;
    signal  gt5_txphdlyreset_i              : std_logic;
    signal  gt5_txphinit_i                  : std_logic;
    signal  gt5_txphinitdone_i              : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt5_txdata_i                    : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt5_gthtxn_i                    : std_logic;
    signal  gt5_gthtxp_i                    : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt5_txoutclk_i                  : std_logic;
    signal  gt5_txoutclkfabric_i            : std_logic;
    signal  gt5_txoutclkpcs_i               : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt5_txresetdone_i               : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt5_txcharisk_i                 : std_logic_vector(7 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT6  (X1Y10)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt6_drpaddr_i                   : std_logic_vector(8 downto 0);
    signal  gt6_drpdi_i                     : std_logic_vector(15 downto 0);
    signal  gt6_drpdo_i                     : std_logic_vector(15 downto 0);
    signal  gt6_drpen_i                     : std_logic;
    signal  gt6_drprdy_i                    : std_logic;
    signal  gt6_drpwe_i                     : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt6_eyescanreset_i              : std_logic;
    signal  gt6_rxuserrdy_i                 : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt6_eyescandataerror_i          : std_logic;
    signal  gt6_eyescantrigger_i            : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt6_rxslide_i                   : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt6_dmonitorout_i               : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt6_rxdata_i                    : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt6_rxdisperr_i                 : std_logic_vector(7 downto 0);
    signal  gt6_rxnotintable_i              : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt6_gthrxn_i                    : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt6_rxdlyen_i                   : std_logic;
    signal  gt6_rxdlysreset_i               : std_logic;
    signal  gt6_rxdlysresetdone_i           : std_logic;
    signal  gt6_rxphalign_i                 : std_logic;
    signal  gt6_rxphaligndone_i             : std_logic;
    signal  gt6_rxphalignen_i               : std_logic;
    signal  gt6_rxphdlyreset_i              : std_logic;
    signal  gt6_rxphmonitor_i               : std_logic_vector(4 downto 0);
    signal  gt6_rxphslipmonitor_i           : std_logic_vector(4 downto 0);
    signal  gt6_rxsyncallin_i               : std_logic;
    signal  gt6_rxsyncdone_i                : std_logic;
    signal  gt6_rxsyncin_i                  : std_logic;
    signal  gt6_rxsyncmode_i                : std_logic;
    signal  gt6_rxsyncout_i                 : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt6_rxbyteisaligned_i           : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt6_rxlpmhfhold_i               : std_logic;
    signal  gt6_rxlpmlfhold_i               : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt6_rxmonitorout_i              : std_logic_vector(6 downto 0);
    signal  gt6_rxmonitorsel_i              : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt6_rxoutclk_i                  : std_logic;
    signal  gt6_rxoutclkfabric_i            : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt6_gtrxreset_i                 : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt6_rxcharisk_i                 : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt6_gthrxp_i                    : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt6_rxresetdone_i               : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt6_gttxreset_i                 : std_logic;
    signal  gt6_txuserrdy_i                 : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt6_txdlyen_i                   : std_logic;
    signal  gt6_txdlysreset_i               : std_logic;
    signal  gt6_txdlysresetdone_i           : std_logic;
    signal  gt6_txphalign_i                 : std_logic;
    signal  gt6_txphaligndone_i             : std_logic;
    signal  gt6_txphalignen_i               : std_logic;
    signal  gt6_txphdlyreset_i              : std_logic;
    signal  gt6_txphinit_i                  : std_logic;
    signal  gt6_txphinitdone_i              : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt6_txdata_i                    : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt6_gthtxn_i                    : std_logic;
    signal  gt6_gthtxp_i                    : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt6_txoutclk_i                  : std_logic;
    signal  gt6_txoutclkfabric_i            : std_logic;
    signal  gt6_txoutclkpcs_i               : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt6_txresetdone_i               : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt6_txcharisk_i                 : std_logic_vector(7 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT7  (X1Y11)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt7_drpaddr_i                   : std_logic_vector(8 downto 0);
    signal  gt7_drpdi_i                     : std_logic_vector(15 downto 0);
    signal  gt7_drpdo_i                     : std_logic_vector(15 downto 0);
    signal  gt7_drpen_i                     : std_logic;
    signal  gt7_drprdy_i                    : std_logic;
    signal  gt7_drpwe_i                     : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt7_eyescanreset_i              : std_logic;
    signal  gt7_rxuserrdy_i                 : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt7_eyescandataerror_i          : std_logic;
    signal  gt7_eyescantrigger_i            : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt7_rxslide_i                   : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt7_dmonitorout_i               : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt7_rxdata_i                    : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt7_rxdisperr_i                 : std_logic_vector(7 downto 0);
    signal  gt7_rxnotintable_i              : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt7_gthrxn_i                    : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt7_rxdlyen_i                   : std_logic;
    signal  gt7_rxdlysreset_i               : std_logic;
    signal  gt7_rxdlysresetdone_i           : std_logic;
    signal  gt7_rxphalign_i                 : std_logic;
    signal  gt7_rxphaligndone_i             : std_logic;
    signal  gt7_rxphalignen_i               : std_logic;
    signal  gt7_rxphdlyreset_i              : std_logic;
    signal  gt7_rxphmonitor_i               : std_logic_vector(4 downto 0);
    signal  gt7_rxphslipmonitor_i           : std_logic_vector(4 downto 0);
    signal  gt7_rxsyncallin_i               : std_logic;
    signal  gt7_rxsyncdone_i                : std_logic;
    signal  gt7_rxsyncin_i                  : std_logic;
    signal  gt7_rxsyncmode_i                : std_logic;
    signal  gt7_rxsyncout_i                 : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt7_rxbyteisaligned_i           : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt7_rxlpmhfhold_i               : std_logic;
    signal  gt7_rxlpmlfhold_i               : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt7_rxmonitorout_i              : std_logic_vector(6 downto 0);
    signal  gt7_rxmonitorsel_i              : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt7_rxoutclk_i                  : std_logic;
    signal  gt7_rxoutclkfabric_i            : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt7_gtrxreset_i                 : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt7_rxcharisk_i                 : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt7_gthrxp_i                    : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt7_rxresetdone_i               : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt7_gttxreset_i                 : std_logic;
    signal  gt7_txuserrdy_i                 : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt7_txdlyen_i                   : std_logic;
    signal  gt7_txdlysreset_i               : std_logic;
    signal  gt7_txdlysresetdone_i           : std_logic;
    signal  gt7_txphalign_i                 : std_logic;
    signal  gt7_txphaligndone_i             : std_logic;
    signal  gt7_txphalignen_i               : std_logic;
    signal  gt7_txphdlyreset_i              : std_logic;
    signal  gt7_txphinit_i                  : std_logic;
    signal  gt7_txphinitdone_i              : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt7_txdata_i                    : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt7_gthtxn_i                    : std_logic;
    signal  gt7_gthtxp_i                    : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt7_txoutclk_i                  : std_logic;
    signal  gt7_txoutclkfabric_i            : std_logic;
    signal  gt7_txoutclkpcs_i               : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt7_txresetdone_i               : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt7_txcharisk_i                 : std_logic_vector(7 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT8  (X1Y12)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt8_drpaddr_i                   : std_logic_vector(8 downto 0);
    signal  gt8_drpdi_i                     : std_logic_vector(15 downto 0);
    signal  gt8_drpdo_i                     : std_logic_vector(15 downto 0);
    signal  gt8_drpen_i                     : std_logic;
    signal  gt8_drprdy_i                    : std_logic;
    signal  gt8_drpwe_i                     : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt8_eyescanreset_i              : std_logic;
    signal  gt8_rxuserrdy_i                 : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt8_eyescandataerror_i          : std_logic;
    signal  gt8_eyescantrigger_i            : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt8_rxslide_i                   : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt8_dmonitorout_i               : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt8_rxdata_i                    : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt8_rxdisperr_i                 : std_logic_vector(7 downto 0);
    signal  gt8_rxnotintable_i              : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt8_gthrxn_i                    : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt8_rxdlyen_i                   : std_logic;
    signal  gt8_rxdlysreset_i               : std_logic;
    signal  gt8_rxdlysresetdone_i           : std_logic;
    signal  gt8_rxphalign_i                 : std_logic;
    signal  gt8_rxphaligndone_i             : std_logic;
    signal  gt8_rxphalignen_i               : std_logic;
    signal  gt8_rxphdlyreset_i              : std_logic;
    signal  gt8_rxphmonitor_i               : std_logic_vector(4 downto 0);
    signal  gt8_rxphslipmonitor_i           : std_logic_vector(4 downto 0);
    signal  gt8_rxsyncallin_i               : std_logic;
    signal  gt8_rxsyncdone_i                : std_logic;
    signal  gt8_rxsyncin_i                  : std_logic;
    signal  gt8_rxsyncmode_i                : std_logic;
    signal  gt8_rxsyncout_i                 : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt8_rxbyteisaligned_i           : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt8_rxlpmhfhold_i               : std_logic;
    signal  gt8_rxlpmlfhold_i               : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt8_rxmonitorout_i              : std_logic_vector(6 downto 0);
    signal  gt8_rxmonitorsel_i              : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt8_rxoutclk_i                  : std_logic;
    signal  gt8_rxoutclkfabric_i            : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt8_gtrxreset_i                 : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt8_rxcharisk_i                 : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt8_gthrxp_i                    : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt8_rxresetdone_i               : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt8_gttxreset_i                 : std_logic;
    signal  gt8_txuserrdy_i                 : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt8_txdlyen_i                   : std_logic;
    signal  gt8_txdlysreset_i               : std_logic;
    signal  gt8_txdlysresetdone_i           : std_logic;
    signal  gt8_txphalign_i                 : std_logic;
    signal  gt8_txphaligndone_i             : std_logic;
    signal  gt8_txphalignen_i               : std_logic;
    signal  gt8_txphdlyreset_i              : std_logic;
    signal  gt8_txphinit_i                  : std_logic;
    signal  gt8_txphinitdone_i              : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt8_txdata_i                    : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt8_gthtxn_i                    : std_logic;
    signal  gt8_gthtxp_i                    : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt8_txoutclk_i                  : std_logic;
    signal  gt8_txoutclkfabric_i            : std_logic;
    signal  gt8_txoutclkpcs_i               : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt8_txresetdone_i               : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt8_txcharisk_i                 : std_logic_vector(7 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT9  (X1Y13)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt9_drpaddr_i                   : std_logic_vector(8 downto 0);
    signal  gt9_drpdi_i                     : std_logic_vector(15 downto 0);
    signal  gt9_drpdo_i                     : std_logic_vector(15 downto 0);
    signal  gt9_drpen_i                     : std_logic;
    signal  gt9_drprdy_i                    : std_logic;
    signal  gt9_drpwe_i                     : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt9_eyescanreset_i              : std_logic;
    signal  gt9_rxuserrdy_i                 : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt9_eyescandataerror_i          : std_logic;
    signal  gt9_eyescantrigger_i            : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt9_rxslide_i                   : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt9_dmonitorout_i               : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt9_rxdata_i                    : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt9_rxdisperr_i                 : std_logic_vector(7 downto 0);
    signal  gt9_rxnotintable_i              : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt9_gthrxn_i                    : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt9_rxdlyen_i                   : std_logic;
    signal  gt9_rxdlysreset_i               : std_logic;
    signal  gt9_rxdlysresetdone_i           : std_logic;
    signal  gt9_rxphalign_i                 : std_logic;
    signal  gt9_rxphaligndone_i             : std_logic;
    signal  gt9_rxphalignen_i               : std_logic;
    signal  gt9_rxphdlyreset_i              : std_logic;
    signal  gt9_rxphmonitor_i               : std_logic_vector(4 downto 0);
    signal  gt9_rxphslipmonitor_i           : std_logic_vector(4 downto 0);
    signal  gt9_rxsyncallin_i               : std_logic;
    signal  gt9_rxsyncdone_i                : std_logic;
    signal  gt9_rxsyncin_i                  : std_logic;
    signal  gt9_rxsyncmode_i                : std_logic;
    signal  gt9_rxsyncout_i                 : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt9_rxbyteisaligned_i           : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt9_rxlpmhfhold_i               : std_logic;
    signal  gt9_rxlpmlfhold_i               : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt9_rxmonitorout_i              : std_logic_vector(6 downto 0);
    signal  gt9_rxmonitorsel_i              : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt9_rxoutclk_i                  : std_logic;
    signal  gt9_rxoutclkfabric_i            : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt9_gtrxreset_i                 : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt9_rxcharisk_i                 : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt9_gthrxp_i                    : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt9_rxresetdone_i               : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt9_gttxreset_i                 : std_logic;
    signal  gt9_txuserrdy_i                 : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt9_txdlyen_i                   : std_logic;
    signal  gt9_txdlysreset_i               : std_logic;
    signal  gt9_txdlysresetdone_i           : std_logic;
    signal  gt9_txphalign_i                 : std_logic;
    signal  gt9_txphaligndone_i             : std_logic;
    signal  gt9_txphalignen_i               : std_logic;
    signal  gt9_txphdlyreset_i              : std_logic;
    signal  gt9_txphinit_i                  : std_logic;
    signal  gt9_txphinitdone_i              : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt9_txdata_i                    : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt9_gthtxn_i                    : std_logic;
    signal  gt9_gthtxp_i                    : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt9_txoutclk_i                  : std_logic;
    signal  gt9_txoutclkfabric_i            : std_logic;
    signal  gt9_txoutclkpcs_i               : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt9_txresetdone_i               : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt9_txcharisk_i                 : std_logic_vector(7 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT10  (X1Y14)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt10_drpaddr_i                  : std_logic_vector(8 downto 0);
    signal  gt10_drpdi_i                    : std_logic_vector(15 downto 0);
    signal  gt10_drpdo_i                    : std_logic_vector(15 downto 0);
    signal  gt10_drpen_i                    : std_logic;
    signal  gt10_drprdy_i                   : std_logic;
    signal  gt10_drpwe_i                    : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt10_eyescanreset_i             : std_logic;
    signal  gt10_rxuserrdy_i                : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt10_eyescandataerror_i         : std_logic;
    signal  gt10_eyescantrigger_i           : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt10_rxslide_i                  : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt10_dmonitorout_i              : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt10_rxdata_i                   : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt10_rxdisperr_i                : std_logic_vector(7 downto 0);
    signal  gt10_rxnotintable_i             : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt10_gthrxn_i                   : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt10_rxdlyen_i                  : std_logic;
    signal  gt10_rxdlysreset_i              : std_logic;
    signal  gt10_rxdlysresetdone_i          : std_logic;
    signal  gt10_rxphalign_i                : std_logic;
    signal  gt10_rxphaligndone_i            : std_logic;
    signal  gt10_rxphalignen_i              : std_logic;
    signal  gt10_rxphdlyreset_i             : std_logic;
    signal  gt10_rxphmonitor_i              : std_logic_vector(4 downto 0);
    signal  gt10_rxphslipmonitor_i          : std_logic_vector(4 downto 0);
    signal  gt10_rxsyncallin_i              : std_logic;
    signal  gt10_rxsyncdone_i               : std_logic;
    signal  gt10_rxsyncin_i                 : std_logic;
    signal  gt10_rxsyncmode_i               : std_logic;
    signal  gt10_rxsyncout_i                : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt10_rxbyteisaligned_i          : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt10_rxlpmhfhold_i              : std_logic;
    signal  gt10_rxlpmlfhold_i              : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt10_rxmonitorout_i             : std_logic_vector(6 downto 0);
    signal  gt10_rxmonitorsel_i             : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt10_rxoutclk_i                 : std_logic;
    signal  gt10_rxoutclkfabric_i           : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt10_gtrxreset_i                : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt10_rxcharisk_i                : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt10_gthrxp_i                   : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt10_rxresetdone_i              : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt10_gttxreset_i                : std_logic;
    signal  gt10_txuserrdy_i                : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt10_txdlyen_i                  : std_logic;
    signal  gt10_txdlysreset_i              : std_logic;
    signal  gt10_txdlysresetdone_i          : std_logic;
    signal  gt10_txphalign_i                : std_logic;
    signal  gt10_txphaligndone_i            : std_logic;
    signal  gt10_txphalignen_i              : std_logic;
    signal  gt10_txphdlyreset_i             : std_logic;
    signal  gt10_txphinit_i                 : std_logic;
    signal  gt10_txphinitdone_i             : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt10_txdata_i                   : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt10_gthtxn_i                   : std_logic;
    signal  gt10_gthtxp_i                   : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt10_txoutclk_i                 : std_logic;
    signal  gt10_txoutclkfabric_i           : std_logic;
    signal  gt10_txoutclkpcs_i              : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt10_txresetdone_i              : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt10_txcharisk_i                : std_logic_vector(7 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT11  (X1Y15)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt11_drpaddr_i                  : std_logic_vector(8 downto 0);
    signal  gt11_drpdi_i                    : std_logic_vector(15 downto 0);
    signal  gt11_drpdo_i                    : std_logic_vector(15 downto 0);
    signal  gt11_drpen_i                    : std_logic;
    signal  gt11_drprdy_i                   : std_logic;
    signal  gt11_drpwe_i                    : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt11_eyescanreset_i             : std_logic;
    signal  gt11_rxuserrdy_i                : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt11_eyescandataerror_i         : std_logic;
    signal  gt11_eyescantrigger_i           : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt11_rxslide_i                  : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt11_dmonitorout_i              : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt11_rxdata_i                   : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt11_rxdisperr_i                : std_logic_vector(7 downto 0);
    signal  gt11_rxnotintable_i             : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt11_gthrxn_i                   : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt11_rxdlyen_i                  : std_logic;
    signal  gt11_rxdlysreset_i              : std_logic;
    signal  gt11_rxdlysresetdone_i          : std_logic;
    signal  gt11_rxphalign_i                : std_logic;
    signal  gt11_rxphaligndone_i            : std_logic;
    signal  gt11_rxphalignen_i              : std_logic;
    signal  gt11_rxphdlyreset_i             : std_logic;
    signal  gt11_rxphmonitor_i              : std_logic_vector(4 downto 0);
    signal  gt11_rxphslipmonitor_i          : std_logic_vector(4 downto 0);
    signal  gt11_rxsyncallin_i              : std_logic;
    signal  gt11_rxsyncdone_i               : std_logic;
    signal  gt11_rxsyncin_i                 : std_logic;
    signal  gt11_rxsyncmode_i               : std_logic;
    signal  gt11_rxsyncout_i                : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt11_rxbyteisaligned_i          : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt11_rxlpmhfhold_i              : std_logic;
    signal  gt11_rxlpmlfhold_i              : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt11_rxmonitorout_i             : std_logic_vector(6 downto 0);
    signal  gt11_rxmonitorsel_i             : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt11_rxoutclk_i                 : std_logic;
    signal  gt11_rxoutclkfabric_i           : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt11_gtrxreset_i                : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt11_rxcharisk_i                : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt11_gthrxp_i                   : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt11_rxresetdone_i              : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt11_gttxreset_i                : std_logic;
    signal  gt11_txuserrdy_i                : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt11_txdlyen_i                  : std_logic;
    signal  gt11_txdlysreset_i              : std_logic;
    signal  gt11_txdlysresetdone_i          : std_logic;
    signal  gt11_txphalign_i                : std_logic;
    signal  gt11_txphaligndone_i            : std_logic;
    signal  gt11_txphalignen_i              : std_logic;
    signal  gt11_txphdlyreset_i             : std_logic;
    signal  gt11_txphinit_i                 : std_logic;
    signal  gt11_txphinitdone_i             : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt11_txdata_i                   : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt11_gthtxn_i                   : std_logic;
    signal  gt11_gthtxp_i                   : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt11_txoutclk_i                 : std_logic;
    signal  gt11_txoutclkfabric_i           : std_logic;
    signal  gt11_txoutclkpcs_i              : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt11_txresetdone_i              : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt11_txcharisk_i                : std_logic_vector(7 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT12  (X1Y16)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt12_drpaddr_i                  : std_logic_vector(8 downto 0);
    signal  gt12_drpdi_i                    : std_logic_vector(15 downto 0);
    signal  gt12_drpdo_i                    : std_logic_vector(15 downto 0);
    signal  gt12_drpen_i                    : std_logic;
    signal  gt12_drprdy_i                   : std_logic;
    signal  gt12_drpwe_i                    : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt12_eyescanreset_i             : std_logic;
    signal  gt12_rxuserrdy_i                : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt12_eyescandataerror_i         : std_logic;
    signal  gt12_eyescantrigger_i           : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt12_rxslide_i                  : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt12_dmonitorout_i              : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt12_rxdata_i                   : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt12_rxdisperr_i                : std_logic_vector(7 downto 0);
    signal  gt12_rxnotintable_i             : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt12_gthrxn_i                   : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt12_rxdlyen_i                  : std_logic;
    signal  gt12_rxdlysreset_i              : std_logic;
    signal  gt12_rxdlysresetdone_i          : std_logic;
    signal  gt12_rxphalign_i                : std_logic;
    signal  gt12_rxphaligndone_i            : std_logic;
    signal  gt12_rxphalignen_i              : std_logic;
    signal  gt12_rxphdlyreset_i             : std_logic;
    signal  gt12_rxphmonitor_i              : std_logic_vector(4 downto 0);
    signal  gt12_rxphslipmonitor_i          : std_logic_vector(4 downto 0);
    signal  gt12_rxsyncallin_i              : std_logic;
    signal  gt12_rxsyncdone_i               : std_logic;
    signal  gt12_rxsyncin_i                 : std_logic;
    signal  gt12_rxsyncmode_i               : std_logic;
    signal  gt12_rxsyncout_i                : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt12_rxbyteisaligned_i          : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt12_rxlpmhfhold_i              : std_logic;
    signal  gt12_rxlpmlfhold_i              : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt12_rxmonitorout_i             : std_logic_vector(6 downto 0);
    signal  gt12_rxmonitorsel_i             : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt12_rxoutclk_i                 : std_logic;
    signal  gt12_rxoutclkfabric_i           : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt12_gtrxreset_i                : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt12_rxcharisk_i                : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt12_gthrxp_i                   : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt12_rxresetdone_i              : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt12_gttxreset_i                : std_logic;
    signal  gt12_txuserrdy_i                : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt12_txdlyen_i                  : std_logic;
    signal  gt12_txdlysreset_i              : std_logic;
    signal  gt12_txdlysresetdone_i          : std_logic;
    signal  gt12_txphalign_i                : std_logic;
    signal  gt12_txphaligndone_i            : std_logic;
    signal  gt12_txphalignen_i              : std_logic;
    signal  gt12_txphdlyreset_i             : std_logic;
    signal  gt12_txphinit_i                 : std_logic;
    signal  gt12_txphinitdone_i             : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt12_txdata_i                   : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt12_gthtxn_i                   : std_logic;
    signal  gt12_gthtxp_i                   : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt12_txoutclk_i                 : std_logic;
    signal  gt12_txoutclkfabric_i           : std_logic;
    signal  gt12_txoutclkpcs_i              : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt12_txresetdone_i              : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt12_txcharisk_i                : std_logic_vector(7 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT13  (X1Y17)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt13_drpaddr_i                  : std_logic_vector(8 downto 0);
    signal  gt13_drpdi_i                    : std_logic_vector(15 downto 0);
    signal  gt13_drpdo_i                    : std_logic_vector(15 downto 0);
    signal  gt13_drpen_i                    : std_logic;
    signal  gt13_drprdy_i                   : std_logic;
    signal  gt13_drpwe_i                    : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt13_eyescanreset_i             : std_logic;
    signal  gt13_rxuserrdy_i                : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt13_eyescandataerror_i         : std_logic;
    signal  gt13_eyescantrigger_i           : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt13_rxslide_i                  : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt13_dmonitorout_i              : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt13_rxdata_i                   : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt13_rxdisperr_i                : std_logic_vector(7 downto 0);
    signal  gt13_rxnotintable_i             : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt13_gthrxn_i                   : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt13_rxdlyen_i                  : std_logic;
    signal  gt13_rxdlysreset_i              : std_logic;
    signal  gt13_rxdlysresetdone_i          : std_logic;
    signal  gt13_rxphalign_i                : std_logic;
    signal  gt13_rxphaligndone_i            : std_logic;
    signal  gt13_rxphalignen_i              : std_logic;
    signal  gt13_rxphdlyreset_i             : std_logic;
    signal  gt13_rxphmonitor_i              : std_logic_vector(4 downto 0);
    signal  gt13_rxphslipmonitor_i          : std_logic_vector(4 downto 0);
    signal  gt13_rxsyncallin_i              : std_logic;
    signal  gt13_rxsyncdone_i               : std_logic;
    signal  gt13_rxsyncin_i                 : std_logic;
    signal  gt13_rxsyncmode_i               : std_logic;
    signal  gt13_rxsyncout_i                : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt13_rxbyteisaligned_i          : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt13_rxlpmhfhold_i              : std_logic;
    signal  gt13_rxlpmlfhold_i              : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt13_rxmonitorout_i             : std_logic_vector(6 downto 0);
    signal  gt13_rxmonitorsel_i             : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt13_rxoutclk_i                 : std_logic;
    signal  gt13_rxoutclkfabric_i           : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt13_gtrxreset_i                : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt13_rxcharisk_i                : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt13_gthrxp_i                   : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt13_rxresetdone_i              : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt13_gttxreset_i                : std_logic;
    signal  gt13_txuserrdy_i                : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt13_txdlyen_i                  : std_logic;
    signal  gt13_txdlysreset_i              : std_logic;
    signal  gt13_txdlysresetdone_i          : std_logic;
    signal  gt13_txphalign_i                : std_logic;
    signal  gt13_txphaligndone_i            : std_logic;
    signal  gt13_txphalignen_i              : std_logic;
    signal  gt13_txphdlyreset_i             : std_logic;
    signal  gt13_txphinit_i                 : std_logic;
    signal  gt13_txphinitdone_i             : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt13_txdata_i                   : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt13_gthtxn_i                   : std_logic;
    signal  gt13_gthtxp_i                   : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt13_txoutclk_i                 : std_logic;
    signal  gt13_txoutclkfabric_i           : std_logic;
    signal  gt13_txoutclkpcs_i              : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt13_txresetdone_i              : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt13_txcharisk_i                : std_logic_vector(7 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT14  (X1Y18)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt14_drpaddr_i                  : std_logic_vector(8 downto 0);
    signal  gt14_drpdi_i                    : std_logic_vector(15 downto 0);
    signal  gt14_drpdo_i                    : std_logic_vector(15 downto 0);
    signal  gt14_drpen_i                    : std_logic;
    signal  gt14_drprdy_i                   : std_logic;
    signal  gt14_drpwe_i                    : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt14_eyescanreset_i             : std_logic;
    signal  gt14_rxuserrdy_i                : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt14_eyescandataerror_i         : std_logic;
    signal  gt14_eyescantrigger_i           : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt14_rxslide_i                  : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt14_dmonitorout_i              : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt14_rxdata_i                   : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt14_rxdisperr_i                : std_logic_vector(7 downto 0);
    signal  gt14_rxnotintable_i             : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt14_gthrxn_i                   : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt14_rxdlyen_i                  : std_logic;
    signal  gt14_rxdlysreset_i              : std_logic;
    signal  gt14_rxdlysresetdone_i          : std_logic;
    signal  gt14_rxphalign_i                : std_logic;
    signal  gt14_rxphaligndone_i            : std_logic;
    signal  gt14_rxphalignen_i              : std_logic;
    signal  gt14_rxphdlyreset_i             : std_logic;
    signal  gt14_rxphmonitor_i              : std_logic_vector(4 downto 0);
    signal  gt14_rxphslipmonitor_i          : std_logic_vector(4 downto 0);
    signal  gt14_rxsyncallin_i              : std_logic;
    signal  gt14_rxsyncdone_i               : std_logic;
    signal  gt14_rxsyncin_i                 : std_logic;
    signal  gt14_rxsyncmode_i               : std_logic;
    signal  gt14_rxsyncout_i                : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt14_rxbyteisaligned_i          : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt14_rxlpmhfhold_i              : std_logic;
    signal  gt14_rxlpmlfhold_i              : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt14_rxmonitorout_i             : std_logic_vector(6 downto 0);
    signal  gt14_rxmonitorsel_i             : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt14_rxoutclk_i                 : std_logic;
    signal  gt14_rxoutclkfabric_i           : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt14_gtrxreset_i                : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt14_rxcharisk_i                : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt14_gthrxp_i                   : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt14_rxresetdone_i              : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt14_gttxreset_i                : std_logic;
    signal  gt14_txuserrdy_i                : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt14_txdlyen_i                  : std_logic;
    signal  gt14_txdlysreset_i              : std_logic;
    signal  gt14_txdlysresetdone_i          : std_logic;
    signal  gt14_txphalign_i                : std_logic;
    signal  gt14_txphaligndone_i            : std_logic;
    signal  gt14_txphalignen_i              : std_logic;
    signal  gt14_txphdlyreset_i             : std_logic;
    signal  gt14_txphinit_i                 : std_logic;
    signal  gt14_txphinitdone_i             : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt14_txdata_i                   : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt14_gthtxn_i                   : std_logic;
    signal  gt14_gthtxp_i                   : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt14_txoutclk_i                 : std_logic;
    signal  gt14_txoutclkfabric_i           : std_logic;
    signal  gt14_txoutclkpcs_i              : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt14_txresetdone_i              : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt14_txcharisk_i                : std_logic_vector(7 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT15  (X1Y19)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt15_drpaddr_i                  : std_logic_vector(8 downto 0);
    signal  gt15_drpdi_i                    : std_logic_vector(15 downto 0);
    signal  gt15_drpdo_i                    : std_logic_vector(15 downto 0);
    signal  gt15_drpen_i                    : std_logic;
    signal  gt15_drprdy_i                   : std_logic;
    signal  gt15_drpwe_i                    : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt15_eyescanreset_i             : std_logic;
    signal  gt15_rxuserrdy_i                : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt15_eyescandataerror_i         : std_logic;
    signal  gt15_eyescantrigger_i           : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt15_rxslide_i                  : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt15_dmonitorout_i              : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt15_rxdata_i                   : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt15_rxdisperr_i                : std_logic_vector(7 downto 0);
    signal  gt15_rxnotintable_i             : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt15_gthrxn_i                   : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt15_rxdlyen_i                  : std_logic;
    signal  gt15_rxdlysreset_i              : std_logic;
    signal  gt15_rxdlysresetdone_i          : std_logic;
    signal  gt15_rxphalign_i                : std_logic;
    signal  gt15_rxphaligndone_i            : std_logic;
    signal  gt15_rxphalignen_i              : std_logic;
    signal  gt15_rxphdlyreset_i             : std_logic;
    signal  gt15_rxphmonitor_i              : std_logic_vector(4 downto 0);
    signal  gt15_rxphslipmonitor_i          : std_logic_vector(4 downto 0);
    signal  gt15_rxsyncallin_i              : std_logic;
    signal  gt15_rxsyncdone_i               : std_logic;
    signal  gt15_rxsyncin_i                 : std_logic;
    signal  gt15_rxsyncmode_i               : std_logic;
    signal  gt15_rxsyncout_i                : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt15_rxbyteisaligned_i          : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt15_rxlpmhfhold_i              : std_logic;
    signal  gt15_rxlpmlfhold_i              : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt15_rxmonitorout_i             : std_logic_vector(6 downto 0);
    signal  gt15_rxmonitorsel_i             : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt15_rxoutclk_i                 : std_logic;
    signal  gt15_rxoutclkfabric_i           : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt15_gtrxreset_i                : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt15_rxcharisk_i                : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt15_gthrxp_i                   : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt15_rxresetdone_i              : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt15_gttxreset_i                : std_logic;
    signal  gt15_txuserrdy_i                : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt15_txdlyen_i                  : std_logic;
    signal  gt15_txdlysreset_i              : std_logic;
    signal  gt15_txdlysresetdone_i          : std_logic;
    signal  gt15_txphalign_i                : std_logic;
    signal  gt15_txphaligndone_i            : std_logic;
    signal  gt15_txphalignen_i              : std_logic;
    signal  gt15_txphdlyreset_i             : std_logic;
    signal  gt15_txphinit_i                 : std_logic;
    signal  gt15_txphinitdone_i             : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt15_txdata_i                   : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt15_gthtxn_i                   : std_logic;
    signal  gt15_gthtxp_i                   : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt15_txoutclk_i                 : std_logic;
    signal  gt15_txoutclkfabric_i           : std_logic;
    signal  gt15_txoutclkpcs_i              : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt15_txresetdone_i              : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt15_txcharisk_i                : std_logic_vector(7 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT16  (X1Y20)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt16_drpaddr_i                  : std_logic_vector(8 downto 0);
    signal  gt16_drpdi_i                    : std_logic_vector(15 downto 0);
    signal  gt16_drpdo_i                    : std_logic_vector(15 downto 0);
    signal  gt16_drpen_i                    : std_logic;
    signal  gt16_drprdy_i                   : std_logic;
    signal  gt16_drpwe_i                    : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt16_eyescanreset_i             : std_logic;
    signal  gt16_rxuserrdy_i                : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt16_eyescandataerror_i         : std_logic;
    signal  gt16_eyescantrigger_i           : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt16_rxslide_i                  : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt16_dmonitorout_i              : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt16_rxdata_i                   : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt16_rxdisperr_i                : std_logic_vector(7 downto 0);
    signal  gt16_rxnotintable_i             : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt16_gthrxn_i                   : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt16_rxdlyen_i                  : std_logic;
    signal  gt16_rxdlysreset_i              : std_logic;
    signal  gt16_rxdlysresetdone_i          : std_logic;
    signal  gt16_rxphalign_i                : std_logic;
    signal  gt16_rxphaligndone_i            : std_logic;
    signal  gt16_rxphalignen_i              : std_logic;
    signal  gt16_rxphdlyreset_i             : std_logic;
    signal  gt16_rxphmonitor_i              : std_logic_vector(4 downto 0);
    signal  gt16_rxphslipmonitor_i          : std_logic_vector(4 downto 0);
    signal  gt16_rxsyncallin_i              : std_logic;
    signal  gt16_rxsyncdone_i               : std_logic;
    signal  gt16_rxsyncin_i                 : std_logic;
    signal  gt16_rxsyncmode_i               : std_logic;
    signal  gt16_rxsyncout_i                : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt16_rxbyteisaligned_i          : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt16_rxlpmhfhold_i              : std_logic;
    signal  gt16_rxlpmlfhold_i              : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt16_rxmonitorout_i             : std_logic_vector(6 downto 0);
    signal  gt16_rxmonitorsel_i             : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt16_rxoutclk_i                 : std_logic;
    signal  gt16_rxoutclkfabric_i           : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt16_gtrxreset_i                : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt16_rxcharisk_i                : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt16_gthrxp_i                   : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt16_rxresetdone_i              : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt16_gttxreset_i                : std_logic;
    signal  gt16_txuserrdy_i                : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt16_txdlyen_i                  : std_logic;
    signal  gt16_txdlysreset_i              : std_logic;
    signal  gt16_txdlysresetdone_i          : std_logic;
    signal  gt16_txphalign_i                : std_logic;
    signal  gt16_txphaligndone_i            : std_logic;
    signal  gt16_txphalignen_i              : std_logic;
    signal  gt16_txphdlyreset_i             : std_logic;
    signal  gt16_txphinit_i                 : std_logic;
    signal  gt16_txphinitdone_i             : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt16_txdata_i                   : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt16_gthtxn_i                   : std_logic;
    signal  gt16_gthtxp_i                   : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt16_txoutclk_i                 : std_logic;
    signal  gt16_txoutclkfabric_i           : std_logic;
    signal  gt16_txoutclkpcs_i              : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt16_txresetdone_i              : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt16_txcharisk_i                : std_logic_vector(7 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT17  (X1Y21)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt17_drpaddr_i                  : std_logic_vector(8 downto 0);
    signal  gt17_drpdi_i                    : std_logic_vector(15 downto 0);
    signal  gt17_drpdo_i                    : std_logic_vector(15 downto 0);
    signal  gt17_drpen_i                    : std_logic;
    signal  gt17_drprdy_i                   : std_logic;
    signal  gt17_drpwe_i                    : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt17_eyescanreset_i             : std_logic;
    signal  gt17_rxuserrdy_i                : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt17_eyescandataerror_i         : std_logic;
    signal  gt17_eyescantrigger_i           : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt17_rxslide_i                  : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt17_dmonitorout_i              : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt17_rxdata_i                   : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt17_rxdisperr_i                : std_logic_vector(7 downto 0);
    signal  gt17_rxnotintable_i             : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt17_gthrxn_i                   : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt17_rxdlyen_i                  : std_logic;
    signal  gt17_rxdlysreset_i              : std_logic;
    signal  gt17_rxdlysresetdone_i          : std_logic;
    signal  gt17_rxphalign_i                : std_logic;
    signal  gt17_rxphaligndone_i            : std_logic;
    signal  gt17_rxphalignen_i              : std_logic;
    signal  gt17_rxphdlyreset_i             : std_logic;
    signal  gt17_rxphmonitor_i              : std_logic_vector(4 downto 0);
    signal  gt17_rxphslipmonitor_i          : std_logic_vector(4 downto 0);
    signal  gt17_rxsyncallin_i              : std_logic;
    signal  gt17_rxsyncdone_i               : std_logic;
    signal  gt17_rxsyncin_i                 : std_logic;
    signal  gt17_rxsyncmode_i               : std_logic;
    signal  gt17_rxsyncout_i                : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt17_rxbyteisaligned_i          : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt17_rxlpmhfhold_i              : std_logic;
    signal  gt17_rxlpmlfhold_i              : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt17_rxmonitorout_i             : std_logic_vector(6 downto 0);
    signal  gt17_rxmonitorsel_i             : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt17_rxoutclk_i                 : std_logic;
    signal  gt17_rxoutclkfabric_i           : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt17_gtrxreset_i                : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt17_rxcharisk_i                : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt17_gthrxp_i                   : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt17_rxresetdone_i              : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt17_gttxreset_i                : std_logic;
    signal  gt17_txuserrdy_i                : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt17_txdlyen_i                  : std_logic;
    signal  gt17_txdlysreset_i              : std_logic;
    signal  gt17_txdlysresetdone_i          : std_logic;
    signal  gt17_txphalign_i                : std_logic;
    signal  gt17_txphaligndone_i            : std_logic;
    signal  gt17_txphalignen_i              : std_logic;
    signal  gt17_txphdlyreset_i             : std_logic;
    signal  gt17_txphinit_i                 : std_logic;
    signal  gt17_txphinitdone_i             : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt17_txdata_i                   : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt17_gthtxn_i                   : std_logic;
    signal  gt17_gthtxp_i                   : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt17_txoutclk_i                 : std_logic;
    signal  gt17_txoutclkfabric_i           : std_logic;
    signal  gt17_txoutclkpcs_i              : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt17_txresetdone_i              : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt17_txcharisk_i                : std_logic_vector(7 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT18  (X1Y22)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt18_drpaddr_i                  : std_logic_vector(8 downto 0);
    signal  gt18_drpdi_i                    : std_logic_vector(15 downto 0);
    signal  gt18_drpdo_i                    : std_logic_vector(15 downto 0);
    signal  gt18_drpen_i                    : std_logic;
    signal  gt18_drprdy_i                   : std_logic;
    signal  gt18_drpwe_i                    : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt18_eyescanreset_i             : std_logic;
    signal  gt18_rxuserrdy_i                : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt18_eyescandataerror_i         : std_logic;
    signal  gt18_eyescantrigger_i           : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt18_rxslide_i                  : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt18_dmonitorout_i              : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt18_rxdata_i                   : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt18_rxdisperr_i                : std_logic_vector(7 downto 0);
    signal  gt18_rxnotintable_i             : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt18_gthrxn_i                   : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt18_rxdlyen_i                  : std_logic;
    signal  gt18_rxdlysreset_i              : std_logic;
    signal  gt18_rxdlysresetdone_i          : std_logic;
    signal  gt18_rxphalign_i                : std_logic;
    signal  gt18_rxphaligndone_i            : std_logic;
    signal  gt18_rxphalignen_i              : std_logic;
    signal  gt18_rxphdlyreset_i             : std_logic;
    signal  gt18_rxphmonitor_i              : std_logic_vector(4 downto 0);
    signal  gt18_rxphslipmonitor_i          : std_logic_vector(4 downto 0);
    signal  gt18_rxsyncallin_i              : std_logic;
    signal  gt18_rxsyncdone_i               : std_logic;
    signal  gt18_rxsyncin_i                 : std_logic;
    signal  gt18_rxsyncmode_i               : std_logic;
    signal  gt18_rxsyncout_i                : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt18_rxbyteisaligned_i          : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt18_rxlpmhfhold_i              : std_logic;
    signal  gt18_rxlpmlfhold_i              : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt18_rxmonitorout_i             : std_logic_vector(6 downto 0);
    signal  gt18_rxmonitorsel_i             : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt18_rxoutclk_i                 : std_logic;
    signal  gt18_rxoutclkfabric_i           : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt18_gtrxreset_i                : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt18_rxcharisk_i                : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt18_gthrxp_i                   : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt18_rxresetdone_i              : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt18_gttxreset_i                : std_logic;
    signal  gt18_txuserrdy_i                : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt18_txdlyen_i                  : std_logic;
    signal  gt18_txdlysreset_i              : std_logic;
    signal  gt18_txdlysresetdone_i          : std_logic;
    signal  gt18_txphalign_i                : std_logic;
    signal  gt18_txphaligndone_i            : std_logic;
    signal  gt18_txphalignen_i              : std_logic;
    signal  gt18_txphdlyreset_i             : std_logic;
    signal  gt18_txphinit_i                 : std_logic;
    signal  gt18_txphinitdone_i             : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt18_txdata_i                   : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt18_gthtxn_i                   : std_logic;
    signal  gt18_gthtxp_i                   : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt18_txoutclk_i                 : std_logic;
    signal  gt18_txoutclkfabric_i           : std_logic;
    signal  gt18_txoutclkpcs_i              : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt18_txresetdone_i              : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt18_txcharisk_i                : std_logic_vector(7 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT19  (X1Y23)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt19_drpaddr_i                  : std_logic_vector(8 downto 0);
    signal  gt19_drpdi_i                    : std_logic_vector(15 downto 0);
    signal  gt19_drpdo_i                    : std_logic_vector(15 downto 0);
    signal  gt19_drpen_i                    : std_logic;
    signal  gt19_drprdy_i                   : std_logic;
    signal  gt19_drpwe_i                    : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt19_eyescanreset_i             : std_logic;
    signal  gt19_rxuserrdy_i                : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt19_eyescandataerror_i         : std_logic;
    signal  gt19_eyescantrigger_i           : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt19_rxslide_i                  : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt19_dmonitorout_i              : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt19_rxdata_i                   : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt19_rxdisperr_i                : std_logic_vector(7 downto 0);
    signal  gt19_rxnotintable_i             : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt19_gthrxn_i                   : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt19_rxdlyen_i                  : std_logic;
    signal  gt19_rxdlysreset_i              : std_logic;
    signal  gt19_rxdlysresetdone_i          : std_logic;
    signal  gt19_rxphalign_i                : std_logic;
    signal  gt19_rxphaligndone_i            : std_logic;
    signal  gt19_rxphalignen_i              : std_logic;
    signal  gt19_rxphdlyreset_i             : std_logic;
    signal  gt19_rxphmonitor_i              : std_logic_vector(4 downto 0);
    signal  gt19_rxphslipmonitor_i          : std_logic_vector(4 downto 0);
    signal  gt19_rxsyncallin_i              : std_logic;
    signal  gt19_rxsyncdone_i               : std_logic;
    signal  gt19_rxsyncin_i                 : std_logic;
    signal  gt19_rxsyncmode_i               : std_logic;
    signal  gt19_rxsyncout_i                : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt19_rxbyteisaligned_i          : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt19_rxlpmhfhold_i              : std_logic;
    signal  gt19_rxlpmlfhold_i              : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt19_rxmonitorout_i             : std_logic_vector(6 downto 0);
    signal  gt19_rxmonitorsel_i             : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt19_rxoutclk_i                 : std_logic;
    signal  gt19_rxoutclkfabric_i           : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt19_gtrxreset_i                : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt19_rxcharisk_i                : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt19_gthrxp_i                   : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt19_rxresetdone_i              : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt19_gttxreset_i                : std_logic;
    signal  gt19_txuserrdy_i                : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt19_txdlyen_i                  : std_logic;
    signal  gt19_txdlysreset_i              : std_logic;
    signal  gt19_txdlysresetdone_i          : std_logic;
    signal  gt19_txphalign_i                : std_logic;
    signal  gt19_txphaligndone_i            : std_logic;
    signal  gt19_txphalignen_i              : std_logic;
    signal  gt19_txphdlyreset_i             : std_logic;
    signal  gt19_txphinit_i                 : std_logic;
    signal  gt19_txphinitdone_i             : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt19_txdata_i                   : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt19_gthtxn_i                   : std_logic;
    signal  gt19_gthtxp_i                   : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt19_txoutclk_i                 : std_logic;
    signal  gt19_txoutclkfabric_i           : std_logic;
    signal  gt19_txoutclkpcs_i              : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt19_txresetdone_i              : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt19_txcharisk_i                : std_logic_vector(7 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT20  (X1Y24)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt20_drpaddr_i                  : std_logic_vector(8 downto 0);
    signal  gt20_drpdi_i                    : std_logic_vector(15 downto 0);
    signal  gt20_drpdo_i                    : std_logic_vector(15 downto 0);
    signal  gt20_drpen_i                    : std_logic;
    signal  gt20_drprdy_i                   : std_logic;
    signal  gt20_drpwe_i                    : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt20_eyescanreset_i             : std_logic;
    signal  gt20_rxuserrdy_i                : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt20_eyescandataerror_i         : std_logic;
    signal  gt20_eyescantrigger_i           : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt20_rxslide_i                  : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt20_dmonitorout_i              : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt20_rxdata_i                   : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt20_rxdisperr_i                : std_logic_vector(7 downto 0);
    signal  gt20_rxnotintable_i             : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt20_gthrxn_i                   : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt20_rxdlyen_i                  : std_logic;
    signal  gt20_rxdlysreset_i              : std_logic;
    signal  gt20_rxdlysresetdone_i          : std_logic;
    signal  gt20_rxphalign_i                : std_logic;
    signal  gt20_rxphaligndone_i            : std_logic;
    signal  gt20_rxphalignen_i              : std_logic;
    signal  gt20_rxphdlyreset_i             : std_logic;
    signal  gt20_rxphmonitor_i              : std_logic_vector(4 downto 0);
    signal  gt20_rxphslipmonitor_i          : std_logic_vector(4 downto 0);
    signal  gt20_rxsyncallin_i              : std_logic;
    signal  gt20_rxsyncdone_i               : std_logic;
    signal  gt20_rxsyncin_i                 : std_logic;
    signal  gt20_rxsyncmode_i               : std_logic;
    signal  gt20_rxsyncout_i                : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt20_rxbyteisaligned_i          : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt20_rxlpmhfhold_i              : std_logic;
    signal  gt20_rxlpmlfhold_i              : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt20_rxmonitorout_i             : std_logic_vector(6 downto 0);
    signal  gt20_rxmonitorsel_i             : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt20_rxoutclk_i                 : std_logic;
    signal  gt20_rxoutclkfabric_i           : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt20_gtrxreset_i                : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt20_rxcharisk_i                : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt20_gthrxp_i                   : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt20_rxresetdone_i              : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt20_gttxreset_i                : std_logic;
    signal  gt20_txuserrdy_i                : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt20_txdlyen_i                  : std_logic;
    signal  gt20_txdlysreset_i              : std_logic;
    signal  gt20_txdlysresetdone_i          : std_logic;
    signal  gt20_txphalign_i                : std_logic;
    signal  gt20_txphaligndone_i            : std_logic;
    signal  gt20_txphalignen_i              : std_logic;
    signal  gt20_txphdlyreset_i             : std_logic;
    signal  gt20_txphinit_i                 : std_logic;
    signal  gt20_txphinitdone_i             : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt20_txdata_i                   : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt20_gthtxn_i                   : std_logic;
    signal  gt20_gthtxp_i                   : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt20_txoutclk_i                 : std_logic;
    signal  gt20_txoutclkfabric_i           : std_logic;
    signal  gt20_txoutclkpcs_i              : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt20_txresetdone_i              : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt20_txcharisk_i                : std_logic_vector(7 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT21  (X1Y25)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt21_drpaddr_i                  : std_logic_vector(8 downto 0);
    signal  gt21_drpdi_i                    : std_logic_vector(15 downto 0);
    signal  gt21_drpdo_i                    : std_logic_vector(15 downto 0);
    signal  gt21_drpen_i                    : std_logic;
    signal  gt21_drprdy_i                   : std_logic;
    signal  gt21_drpwe_i                    : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt21_eyescanreset_i             : std_logic;
    signal  gt21_rxuserrdy_i                : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt21_eyescandataerror_i         : std_logic;
    signal  gt21_eyescantrigger_i           : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt21_rxslide_i                  : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt21_dmonitorout_i              : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt21_rxdata_i                   : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt21_rxdisperr_i                : std_logic_vector(7 downto 0);
    signal  gt21_rxnotintable_i             : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt21_gthrxn_i                   : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt21_rxdlyen_i                  : std_logic;
    signal  gt21_rxdlysreset_i              : std_logic;
    signal  gt21_rxdlysresetdone_i          : std_logic;
    signal  gt21_rxphalign_i                : std_logic;
    signal  gt21_rxphaligndone_i            : std_logic;
    signal  gt21_rxphalignen_i              : std_logic;
    signal  gt21_rxphdlyreset_i             : std_logic;
    signal  gt21_rxphmonitor_i              : std_logic_vector(4 downto 0);
    signal  gt21_rxphslipmonitor_i          : std_logic_vector(4 downto 0);
    signal  gt21_rxsyncallin_i              : std_logic;
    signal  gt21_rxsyncdone_i               : std_logic;
    signal  gt21_rxsyncin_i                 : std_logic;
    signal  gt21_rxsyncmode_i               : std_logic;
    signal  gt21_rxsyncout_i                : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt21_rxbyteisaligned_i          : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt21_rxlpmhfhold_i              : std_logic;
    signal  gt21_rxlpmlfhold_i              : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt21_rxmonitorout_i             : std_logic_vector(6 downto 0);
    signal  gt21_rxmonitorsel_i             : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt21_rxoutclk_i                 : std_logic;
    signal  gt21_rxoutclkfabric_i           : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt21_gtrxreset_i                : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt21_rxcharisk_i                : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt21_gthrxp_i                   : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt21_rxresetdone_i              : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt21_gttxreset_i                : std_logic;
    signal  gt21_txuserrdy_i                : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt21_txdlyen_i                  : std_logic;
    signal  gt21_txdlysreset_i              : std_logic;
    signal  gt21_txdlysresetdone_i          : std_logic;
    signal  gt21_txphalign_i                : std_logic;
    signal  gt21_txphaligndone_i            : std_logic;
    signal  gt21_txphalignen_i              : std_logic;
    signal  gt21_txphdlyreset_i             : std_logic;
    signal  gt21_txphinit_i                 : std_logic;
    signal  gt21_txphinitdone_i             : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt21_txdata_i                   : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt21_gthtxn_i                   : std_logic;
    signal  gt21_gthtxp_i                   : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt21_txoutclk_i                 : std_logic;
    signal  gt21_txoutclkfabric_i           : std_logic;
    signal  gt21_txoutclkpcs_i              : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt21_txresetdone_i              : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt21_txcharisk_i                : std_logic_vector(7 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT22  (X1Y26)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt22_drpaddr_i                  : std_logic_vector(8 downto 0);
    signal  gt22_drpdi_i                    : std_logic_vector(15 downto 0);
    signal  gt22_drpdo_i                    : std_logic_vector(15 downto 0);
    signal  gt22_drpen_i                    : std_logic;
    signal  gt22_drprdy_i                   : std_logic;
    signal  gt22_drpwe_i                    : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt22_eyescanreset_i             : std_logic;
    signal  gt22_rxuserrdy_i                : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt22_eyescandataerror_i         : std_logic;
    signal  gt22_eyescantrigger_i           : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt22_rxslide_i                  : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt22_dmonitorout_i              : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt22_rxdata_i                   : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt22_rxdisperr_i                : std_logic_vector(7 downto 0);
    signal  gt22_rxnotintable_i             : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt22_gthrxn_i                   : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt22_rxdlyen_i                  : std_logic;
    signal  gt22_rxdlysreset_i              : std_logic;
    signal  gt22_rxdlysresetdone_i          : std_logic;
    signal  gt22_rxphalign_i                : std_logic;
    signal  gt22_rxphaligndone_i            : std_logic;
    signal  gt22_rxphalignen_i              : std_logic;
    signal  gt22_rxphdlyreset_i             : std_logic;
    signal  gt22_rxphmonitor_i              : std_logic_vector(4 downto 0);
    signal  gt22_rxphslipmonitor_i          : std_logic_vector(4 downto 0);
    signal  gt22_rxsyncallin_i              : std_logic;
    signal  gt22_rxsyncdone_i               : std_logic;
    signal  gt22_rxsyncin_i                 : std_logic;
    signal  gt22_rxsyncmode_i               : std_logic;
    signal  gt22_rxsyncout_i                : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt22_rxbyteisaligned_i          : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt22_rxlpmhfhold_i              : std_logic;
    signal  gt22_rxlpmlfhold_i              : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt22_rxmonitorout_i             : std_logic_vector(6 downto 0);
    signal  gt22_rxmonitorsel_i             : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt22_rxoutclk_i                 : std_logic;
    signal  gt22_rxoutclkfabric_i           : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt22_gtrxreset_i                : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt22_rxcharisk_i                : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt22_gthrxp_i                   : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt22_rxresetdone_i              : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt22_gttxreset_i                : std_logic;
    signal  gt22_txuserrdy_i                : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt22_txdlyen_i                  : std_logic;
    signal  gt22_txdlysreset_i              : std_logic;
    signal  gt22_txdlysresetdone_i          : std_logic;
    signal  gt22_txphalign_i                : std_logic;
    signal  gt22_txphaligndone_i            : std_logic;
    signal  gt22_txphalignen_i              : std_logic;
    signal  gt22_txphdlyreset_i             : std_logic;
    signal  gt22_txphinit_i                 : std_logic;
    signal  gt22_txphinitdone_i             : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt22_txdata_i                   : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt22_gthtxn_i                   : std_logic;
    signal  gt22_gthtxp_i                   : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt22_txoutclk_i                 : std_logic;
    signal  gt22_txoutclkfabric_i           : std_logic;
    signal  gt22_txoutclkpcs_i              : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt22_txresetdone_i              : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt22_txcharisk_i                : std_logic_vector(7 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT23  (X1Y27)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt23_drpaddr_i                  : std_logic_vector(8 downto 0);
    signal  gt23_drpdi_i                    : std_logic_vector(15 downto 0);
    signal  gt23_drpdo_i                    : std_logic_vector(15 downto 0);
    signal  gt23_drpen_i                    : std_logic;
    signal  gt23_drprdy_i                   : std_logic;
    signal  gt23_drpwe_i                    : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt23_eyescanreset_i             : std_logic;
    signal  gt23_rxuserrdy_i                : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt23_eyescandataerror_i         : std_logic;
    signal  gt23_eyescantrigger_i           : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt23_rxslide_i                  : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt23_dmonitorout_i              : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt23_rxdata_i                   : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt23_rxdisperr_i                : std_logic_vector(7 downto 0);
    signal  gt23_rxnotintable_i             : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt23_gthrxn_i                   : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt23_rxdlyen_i                  : std_logic;
    signal  gt23_rxdlysreset_i              : std_logic;
    signal  gt23_rxdlysresetdone_i          : std_logic;
    signal  gt23_rxphalign_i                : std_logic;
    signal  gt23_rxphaligndone_i            : std_logic;
    signal  gt23_rxphalignen_i              : std_logic;
    signal  gt23_rxphdlyreset_i             : std_logic;
    signal  gt23_rxphmonitor_i              : std_logic_vector(4 downto 0);
    signal  gt23_rxphslipmonitor_i          : std_logic_vector(4 downto 0);
    signal  gt23_rxsyncallin_i              : std_logic;
    signal  gt23_rxsyncdone_i               : std_logic;
    signal  gt23_rxsyncin_i                 : std_logic;
    signal  gt23_rxsyncmode_i               : std_logic;
    signal  gt23_rxsyncout_i                : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt23_rxbyteisaligned_i          : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt23_rxlpmhfhold_i              : std_logic;
    signal  gt23_rxlpmlfhold_i              : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt23_rxmonitorout_i             : std_logic_vector(6 downto 0);
    signal  gt23_rxmonitorsel_i             : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt23_rxoutclk_i                 : std_logic;
    signal  gt23_rxoutclkfabric_i           : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt23_gtrxreset_i                : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt23_rxcharisk_i                : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt23_gthrxp_i                   : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt23_rxresetdone_i              : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt23_gttxreset_i                : std_logic;
    signal  gt23_txuserrdy_i                : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt23_txdlyen_i                  : std_logic;
    signal  gt23_txdlysreset_i              : std_logic;
    signal  gt23_txdlysresetdone_i          : std_logic;
    signal  gt23_txphalign_i                : std_logic;
    signal  gt23_txphaligndone_i            : std_logic;
    signal  gt23_txphalignen_i              : std_logic;
    signal  gt23_txphdlyreset_i             : std_logic;
    signal  gt23_txphinit_i                 : std_logic;
    signal  gt23_txphinitdone_i             : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt23_txdata_i                   : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt23_gthtxn_i                   : std_logic;
    signal  gt23_gthtxp_i                   : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt23_txoutclk_i                 : std_logic;
    signal  gt23_txoutclkfabric_i           : std_logic;
    signal  gt23_txoutclkpcs_i              : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt23_txresetdone_i              : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt23_txcharisk_i                : std_logic_vector(7 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT24  (X1Y28)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt24_drpaddr_i                  : std_logic_vector(8 downto 0);
    signal  gt24_drpdi_i                    : std_logic_vector(15 downto 0);
    signal  gt24_drpdo_i                    : std_logic_vector(15 downto 0);
    signal  gt24_drpen_i                    : std_logic;
    signal  gt24_drprdy_i                   : std_logic;
    signal  gt24_drpwe_i                    : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt24_eyescanreset_i             : std_logic;
    signal  gt24_rxuserrdy_i                : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt24_eyescandataerror_i         : std_logic;
    signal  gt24_eyescantrigger_i           : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt24_rxslide_i                  : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt24_dmonitorout_i              : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt24_rxdata_i                   : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt24_rxdisperr_i                : std_logic_vector(7 downto 0);
    signal  gt24_rxnotintable_i             : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt24_gthrxn_i                   : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt24_rxdlyen_i                  : std_logic;
    signal  gt24_rxdlysreset_i              : std_logic;
    signal  gt24_rxdlysresetdone_i          : std_logic;
    signal  gt24_rxphalign_i                : std_logic;
    signal  gt24_rxphaligndone_i            : std_logic;
    signal  gt24_rxphalignen_i              : std_logic;
    signal  gt24_rxphdlyreset_i             : std_logic;
    signal  gt24_rxphmonitor_i              : std_logic_vector(4 downto 0);
    signal  gt24_rxphslipmonitor_i          : std_logic_vector(4 downto 0);
    signal  gt24_rxsyncallin_i              : std_logic;
    signal  gt24_rxsyncdone_i               : std_logic;
    signal  gt24_rxsyncin_i                 : std_logic;
    signal  gt24_rxsyncmode_i               : std_logic;
    signal  gt24_rxsyncout_i                : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt24_rxbyteisaligned_i          : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt24_rxlpmhfhold_i              : std_logic;
    signal  gt24_rxlpmlfhold_i              : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt24_rxmonitorout_i             : std_logic_vector(6 downto 0);
    signal  gt24_rxmonitorsel_i             : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt24_rxoutclk_i                 : std_logic;
    signal  gt24_rxoutclkfabric_i           : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt24_gtrxreset_i                : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt24_rxcharisk_i                : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt24_gthrxp_i                   : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt24_rxresetdone_i              : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt24_gttxreset_i                : std_logic;
    signal  gt24_txuserrdy_i                : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt24_txdlyen_i                  : std_logic;
    signal  gt24_txdlysreset_i              : std_logic;
    signal  gt24_txdlysresetdone_i          : std_logic;
    signal  gt24_txphalign_i                : std_logic;
    signal  gt24_txphaligndone_i            : std_logic;
    signal  gt24_txphalignen_i              : std_logic;
    signal  gt24_txphdlyreset_i             : std_logic;
    signal  gt24_txphinit_i                 : std_logic;
    signal  gt24_txphinitdone_i             : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt24_txdata_i                   : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt24_gthtxn_i                   : std_logic;
    signal  gt24_gthtxp_i                   : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt24_txoutclk_i                 : std_logic;
    signal  gt24_txoutclkfabric_i           : std_logic;
    signal  gt24_txoutclkpcs_i              : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt24_txresetdone_i              : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt24_txcharisk_i                : std_logic_vector(7 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT25  (X1Y29)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt25_drpaddr_i                  : std_logic_vector(8 downto 0);
    signal  gt25_drpdi_i                    : std_logic_vector(15 downto 0);
    signal  gt25_drpdo_i                    : std_logic_vector(15 downto 0);
    signal  gt25_drpen_i                    : std_logic;
    signal  gt25_drprdy_i                   : std_logic;
    signal  gt25_drpwe_i                    : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt25_eyescanreset_i             : std_logic;
    signal  gt25_rxuserrdy_i                : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt25_eyescandataerror_i         : std_logic;
    signal  gt25_eyescantrigger_i           : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt25_rxslide_i                  : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt25_dmonitorout_i              : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt25_rxdata_i                   : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt25_rxdisperr_i                : std_logic_vector(7 downto 0);
    signal  gt25_rxnotintable_i             : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt25_gthrxn_i                   : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt25_rxdlyen_i                  : std_logic;
    signal  gt25_rxdlysreset_i              : std_logic;
    signal  gt25_rxdlysresetdone_i          : std_logic;
    signal  gt25_rxphalign_i                : std_logic;
    signal  gt25_rxphaligndone_i            : std_logic;
    signal  gt25_rxphalignen_i              : std_logic;
    signal  gt25_rxphdlyreset_i             : std_logic;
    signal  gt25_rxphmonitor_i              : std_logic_vector(4 downto 0);
    signal  gt25_rxphslipmonitor_i          : std_logic_vector(4 downto 0);
    signal  gt25_rxsyncallin_i              : std_logic;
    signal  gt25_rxsyncdone_i               : std_logic;
    signal  gt25_rxsyncin_i                 : std_logic;
    signal  gt25_rxsyncmode_i               : std_logic;
    signal  gt25_rxsyncout_i                : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt25_rxbyteisaligned_i          : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt25_rxlpmhfhold_i              : std_logic;
    signal  gt25_rxlpmlfhold_i              : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt25_rxmonitorout_i             : std_logic_vector(6 downto 0);
    signal  gt25_rxmonitorsel_i             : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt25_rxoutclk_i                 : std_logic;
    signal  gt25_rxoutclkfabric_i           : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt25_gtrxreset_i                : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt25_rxcharisk_i                : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt25_gthrxp_i                   : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt25_rxresetdone_i              : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt25_gttxreset_i                : std_logic;
    signal  gt25_txuserrdy_i                : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt25_txdlyen_i                  : std_logic;
    signal  gt25_txdlysreset_i              : std_logic;
    signal  gt25_txdlysresetdone_i          : std_logic;
    signal  gt25_txphalign_i                : std_logic;
    signal  gt25_txphaligndone_i            : std_logic;
    signal  gt25_txphalignen_i              : std_logic;
    signal  gt25_txphdlyreset_i             : std_logic;
    signal  gt25_txphinit_i                 : std_logic;
    signal  gt25_txphinitdone_i             : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt25_txdata_i                   : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt25_gthtxn_i                   : std_logic;
    signal  gt25_gthtxp_i                   : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt25_txoutclk_i                 : std_logic;
    signal  gt25_txoutclkfabric_i           : std_logic;
    signal  gt25_txoutclkpcs_i              : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt25_txresetdone_i              : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt25_txcharisk_i                : std_logic_vector(7 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT26  (X1Y30)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt26_drpaddr_i                  : std_logic_vector(8 downto 0);
    signal  gt26_drpdi_i                    : std_logic_vector(15 downto 0);
    signal  gt26_drpdo_i                    : std_logic_vector(15 downto 0);
    signal  gt26_drpen_i                    : std_logic;
    signal  gt26_drprdy_i                   : std_logic;
    signal  gt26_drpwe_i                    : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt26_eyescanreset_i             : std_logic;
    signal  gt26_rxuserrdy_i                : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt26_eyescandataerror_i         : std_logic;
    signal  gt26_eyescantrigger_i           : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt26_rxslide_i                  : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt26_dmonitorout_i              : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt26_rxdata_i                   : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt26_rxdisperr_i                : std_logic_vector(7 downto 0);
    signal  gt26_rxnotintable_i             : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt26_gthrxn_i                   : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt26_rxdlyen_i                  : std_logic;
    signal  gt26_rxdlysreset_i              : std_logic;
    signal  gt26_rxdlysresetdone_i          : std_logic;
    signal  gt26_rxphalign_i                : std_logic;
    signal  gt26_rxphaligndone_i            : std_logic;
    signal  gt26_rxphalignen_i              : std_logic;
    signal  gt26_rxphdlyreset_i             : std_logic;
    signal  gt26_rxphmonitor_i              : std_logic_vector(4 downto 0);
    signal  gt26_rxphslipmonitor_i          : std_logic_vector(4 downto 0);
    signal  gt26_rxsyncallin_i              : std_logic;
    signal  gt26_rxsyncdone_i               : std_logic;
    signal  gt26_rxsyncin_i                 : std_logic;
    signal  gt26_rxsyncmode_i               : std_logic;
    signal  gt26_rxsyncout_i                : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt26_rxbyteisaligned_i          : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt26_rxlpmhfhold_i              : std_logic;
    signal  gt26_rxlpmlfhold_i              : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt26_rxmonitorout_i             : std_logic_vector(6 downto 0);
    signal  gt26_rxmonitorsel_i             : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt26_rxoutclk_i                 : std_logic;
    signal  gt26_rxoutclkfabric_i           : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt26_gtrxreset_i                : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt26_rxcharisk_i                : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt26_gthrxp_i                   : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt26_rxresetdone_i              : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt26_gttxreset_i                : std_logic;
    signal  gt26_txuserrdy_i                : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt26_txdlyen_i                  : std_logic;
    signal  gt26_txdlysreset_i              : std_logic;
    signal  gt26_txdlysresetdone_i          : std_logic;
    signal  gt26_txphalign_i                : std_logic;
    signal  gt26_txphaligndone_i            : std_logic;
    signal  gt26_txphalignen_i              : std_logic;
    signal  gt26_txphdlyreset_i             : std_logic;
    signal  gt26_txphinit_i                 : std_logic;
    signal  gt26_txphinitdone_i             : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt26_txdata_i                   : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt26_gthtxn_i                   : std_logic;
    signal  gt26_gthtxp_i                   : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt26_txoutclk_i                 : std_logic;
    signal  gt26_txoutclkfabric_i           : std_logic;
    signal  gt26_txoutclkpcs_i              : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt26_txresetdone_i              : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt26_txcharisk_i                : std_logic_vector(7 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT27  (X1Y31)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt27_drpaddr_i                  : std_logic_vector(8 downto 0);
    signal  gt27_drpdi_i                    : std_logic_vector(15 downto 0);
    signal  gt27_drpdo_i                    : std_logic_vector(15 downto 0);
    signal  gt27_drpen_i                    : std_logic;
    signal  gt27_drprdy_i                   : std_logic;
    signal  gt27_drpwe_i                    : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt27_eyescanreset_i             : std_logic;
    signal  gt27_rxuserrdy_i                : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt27_eyescandataerror_i         : std_logic;
    signal  gt27_eyescantrigger_i           : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt27_rxslide_i                  : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt27_dmonitorout_i              : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt27_rxdata_i                   : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt27_rxdisperr_i                : std_logic_vector(7 downto 0);
    signal  gt27_rxnotintable_i             : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt27_gthrxn_i                   : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt27_rxdlyen_i                  : std_logic;
    signal  gt27_rxdlysreset_i              : std_logic;
    signal  gt27_rxdlysresetdone_i          : std_logic;
    signal  gt27_rxphalign_i                : std_logic;
    signal  gt27_rxphaligndone_i            : std_logic;
    signal  gt27_rxphalignen_i              : std_logic;
    signal  gt27_rxphdlyreset_i             : std_logic;
    signal  gt27_rxphmonitor_i              : std_logic_vector(4 downto 0);
    signal  gt27_rxphslipmonitor_i          : std_logic_vector(4 downto 0);
    signal  gt27_rxsyncallin_i              : std_logic;
    signal  gt27_rxsyncdone_i               : std_logic;
    signal  gt27_rxsyncin_i                 : std_logic;
    signal  gt27_rxsyncmode_i               : std_logic;
    signal  gt27_rxsyncout_i                : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt27_rxbyteisaligned_i          : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt27_rxlpmhfhold_i              : std_logic;
    signal  gt27_rxlpmlfhold_i              : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt27_rxmonitorout_i             : std_logic_vector(6 downto 0);
    signal  gt27_rxmonitorsel_i             : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt27_rxoutclk_i                 : std_logic;
    signal  gt27_rxoutclkfabric_i           : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt27_gtrxreset_i                : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt27_rxcharisk_i                : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt27_gthrxp_i                   : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt27_rxresetdone_i              : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt27_gttxreset_i                : std_logic;
    signal  gt27_txuserrdy_i                : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt27_txdlyen_i                  : std_logic;
    signal  gt27_txdlysreset_i              : std_logic;
    signal  gt27_txdlysresetdone_i          : std_logic;
    signal  gt27_txphalign_i                : std_logic;
    signal  gt27_txphaligndone_i            : std_logic;
    signal  gt27_txphalignen_i              : std_logic;
    signal  gt27_txphdlyreset_i             : std_logic;
    signal  gt27_txphinit_i                 : std_logic;
    signal  gt27_txphinitdone_i             : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt27_txdata_i                   : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt27_gthtxn_i                   : std_logic;
    signal  gt27_gthtxp_i                   : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt27_txoutclk_i                 : std_logic;
    signal  gt27_txoutclkfabric_i           : std_logic;
    signal  gt27_txoutclkpcs_i              : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt27_txresetdone_i              : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt27_txcharisk_i                : std_logic_vector(7 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT28  (X1Y32)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt28_drpaddr_i                  : std_logic_vector(8 downto 0);
    signal  gt28_drpdi_i                    : std_logic_vector(15 downto 0);
    signal  gt28_drpdo_i                    : std_logic_vector(15 downto 0);
    signal  gt28_drpen_i                    : std_logic;
    signal  gt28_drprdy_i                   : std_logic;
    signal  gt28_drpwe_i                    : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt28_eyescanreset_i             : std_logic;
    signal  gt28_rxuserrdy_i                : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt28_eyescandataerror_i         : std_logic;
    signal  gt28_eyescantrigger_i           : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt28_rxslide_i                  : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt28_dmonitorout_i              : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt28_rxdata_i                   : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt28_rxdisperr_i                : std_logic_vector(7 downto 0);
    signal  gt28_rxnotintable_i             : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt28_gthrxn_i                   : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt28_rxdlyen_i                  : std_logic;
    signal  gt28_rxdlysreset_i              : std_logic;
    signal  gt28_rxdlysresetdone_i          : std_logic;
    signal  gt28_rxphalign_i                : std_logic;
    signal  gt28_rxphaligndone_i            : std_logic;
    signal  gt28_rxphalignen_i              : std_logic;
    signal  gt28_rxphdlyreset_i             : std_logic;
    signal  gt28_rxphmonitor_i              : std_logic_vector(4 downto 0);
    signal  gt28_rxphslipmonitor_i          : std_logic_vector(4 downto 0);
    signal  gt28_rxsyncallin_i              : std_logic;
    signal  gt28_rxsyncdone_i               : std_logic;
    signal  gt28_rxsyncin_i                 : std_logic;
    signal  gt28_rxsyncmode_i               : std_logic;
    signal  gt28_rxsyncout_i                : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt28_rxbyteisaligned_i          : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt28_rxlpmhfhold_i              : std_logic;
    signal  gt28_rxlpmlfhold_i              : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt28_rxmonitorout_i             : std_logic_vector(6 downto 0);
    signal  gt28_rxmonitorsel_i             : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt28_rxoutclk_i                 : std_logic;
    signal  gt28_rxoutclkfabric_i           : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt28_gtrxreset_i                : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt28_rxcharisk_i                : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt28_gthrxp_i                   : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt28_rxresetdone_i              : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt28_gttxreset_i                : std_logic;
    signal  gt28_txuserrdy_i                : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt28_txdlyen_i                  : std_logic;
    signal  gt28_txdlysreset_i              : std_logic;
    signal  gt28_txdlysresetdone_i          : std_logic;
    signal  gt28_txphalign_i                : std_logic;
    signal  gt28_txphaligndone_i            : std_logic;
    signal  gt28_txphalignen_i              : std_logic;
    signal  gt28_txphdlyreset_i             : std_logic;
    signal  gt28_txphinit_i                 : std_logic;
    signal  gt28_txphinitdone_i             : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt28_txdata_i                   : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt28_gthtxn_i                   : std_logic;
    signal  gt28_gthtxp_i                   : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt28_txoutclk_i                 : std_logic;
    signal  gt28_txoutclkfabric_i           : std_logic;
    signal  gt28_txoutclkpcs_i              : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt28_txresetdone_i              : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt28_txcharisk_i                : std_logic_vector(7 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT29  (X1Y33)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt29_drpaddr_i                  : std_logic_vector(8 downto 0);
    signal  gt29_drpdi_i                    : std_logic_vector(15 downto 0);
    signal  gt29_drpdo_i                    : std_logic_vector(15 downto 0);
    signal  gt29_drpen_i                    : std_logic;
    signal  gt29_drprdy_i                   : std_logic;
    signal  gt29_drpwe_i                    : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt29_eyescanreset_i             : std_logic;
    signal  gt29_rxuserrdy_i                : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt29_eyescandataerror_i         : std_logic;
    signal  gt29_eyescantrigger_i           : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt29_rxslide_i                  : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt29_dmonitorout_i              : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt29_rxdata_i                   : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt29_rxdisperr_i                : std_logic_vector(7 downto 0);
    signal  gt29_rxnotintable_i             : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt29_gthrxn_i                   : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt29_rxdlyen_i                  : std_logic;
    signal  gt29_rxdlysreset_i              : std_logic;
    signal  gt29_rxdlysresetdone_i          : std_logic;
    signal  gt29_rxphalign_i                : std_logic;
    signal  gt29_rxphaligndone_i            : std_logic;
    signal  gt29_rxphalignen_i              : std_logic;
    signal  gt29_rxphdlyreset_i             : std_logic;
    signal  gt29_rxphmonitor_i              : std_logic_vector(4 downto 0);
    signal  gt29_rxphslipmonitor_i          : std_logic_vector(4 downto 0);
    signal  gt29_rxsyncallin_i              : std_logic;
    signal  gt29_rxsyncdone_i               : std_logic;
    signal  gt29_rxsyncin_i                 : std_logic;
    signal  gt29_rxsyncmode_i               : std_logic;
    signal  gt29_rxsyncout_i                : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt29_rxbyteisaligned_i          : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt29_rxlpmhfhold_i              : std_logic;
    signal  gt29_rxlpmlfhold_i              : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt29_rxmonitorout_i             : std_logic_vector(6 downto 0);
    signal  gt29_rxmonitorsel_i             : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt29_rxoutclk_i                 : std_logic;
    signal  gt29_rxoutclkfabric_i           : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt29_gtrxreset_i                : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt29_rxcharisk_i                : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt29_gthrxp_i                   : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt29_rxresetdone_i              : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt29_gttxreset_i                : std_logic;
    signal  gt29_txuserrdy_i                : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt29_txdlyen_i                  : std_logic;
    signal  gt29_txdlysreset_i              : std_logic;
    signal  gt29_txdlysresetdone_i          : std_logic;
    signal  gt29_txphalign_i                : std_logic;
    signal  gt29_txphaligndone_i            : std_logic;
    signal  gt29_txphalignen_i              : std_logic;
    signal  gt29_txphdlyreset_i             : std_logic;
    signal  gt29_txphinit_i                 : std_logic;
    signal  gt29_txphinitdone_i             : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt29_txdata_i                   : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt29_gthtxn_i                   : std_logic;
    signal  gt29_gthtxp_i                   : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt29_txoutclk_i                 : std_logic;
    signal  gt29_txoutclkfabric_i           : std_logic;
    signal  gt29_txoutclkpcs_i              : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt29_txresetdone_i              : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt29_txcharisk_i                : std_logic_vector(7 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT30  (X1Y34)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt30_drpaddr_i                  : std_logic_vector(8 downto 0);
    signal  gt30_drpdi_i                    : std_logic_vector(15 downto 0);
    signal  gt30_drpdo_i                    : std_logic_vector(15 downto 0);
    signal  gt30_drpen_i                    : std_logic;
    signal  gt30_drprdy_i                   : std_logic;
    signal  gt30_drpwe_i                    : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt30_eyescanreset_i             : std_logic;
    signal  gt30_rxuserrdy_i                : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt30_eyescandataerror_i         : std_logic;
    signal  gt30_eyescantrigger_i           : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt30_rxslide_i                  : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt30_dmonitorout_i              : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt30_rxdata_i                   : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt30_rxdisperr_i                : std_logic_vector(7 downto 0);
    signal  gt30_rxnotintable_i             : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt30_gthrxn_i                   : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt30_rxdlyen_i                  : std_logic;
    signal  gt30_rxdlysreset_i              : std_logic;
    signal  gt30_rxdlysresetdone_i          : std_logic;
    signal  gt30_rxphalign_i                : std_logic;
    signal  gt30_rxphaligndone_i            : std_logic;
    signal  gt30_rxphalignen_i              : std_logic;
    signal  gt30_rxphdlyreset_i             : std_logic;
    signal  gt30_rxphmonitor_i              : std_logic_vector(4 downto 0);
    signal  gt30_rxphslipmonitor_i          : std_logic_vector(4 downto 0);
    signal  gt30_rxsyncallin_i              : std_logic;
    signal  gt30_rxsyncdone_i               : std_logic;
    signal  gt30_rxsyncin_i                 : std_logic;
    signal  gt30_rxsyncmode_i               : std_logic;
    signal  gt30_rxsyncout_i                : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt30_rxbyteisaligned_i          : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt30_rxlpmhfhold_i              : std_logic;
    signal  gt30_rxlpmlfhold_i              : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt30_rxmonitorout_i             : std_logic_vector(6 downto 0);
    signal  gt30_rxmonitorsel_i             : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt30_rxoutclk_i                 : std_logic;
    signal  gt30_rxoutclkfabric_i           : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt30_gtrxreset_i                : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt30_rxcharisk_i                : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt30_gthrxp_i                   : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt30_rxresetdone_i              : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt30_gttxreset_i                : std_logic;
    signal  gt30_txuserrdy_i                : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt30_txdlyen_i                  : std_logic;
    signal  gt30_txdlysreset_i              : std_logic;
    signal  gt30_txdlysresetdone_i          : std_logic;
    signal  gt30_txphalign_i                : std_logic;
    signal  gt30_txphaligndone_i            : std_logic;
    signal  gt30_txphalignen_i              : std_logic;
    signal  gt30_txphdlyreset_i             : std_logic;
    signal  gt30_txphinit_i                 : std_logic;
    signal  gt30_txphinitdone_i             : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt30_txdata_i                   : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt30_gthtxn_i                   : std_logic;
    signal  gt30_gthtxp_i                   : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt30_txoutclk_i                 : std_logic;
    signal  gt30_txoutclkfabric_i           : std_logic;
    signal  gt30_txoutclkpcs_i              : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt30_txresetdone_i              : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt30_txcharisk_i                : std_logic_vector(7 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT31  (X1Y35)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt31_drpaddr_i                  : std_logic_vector(8 downto 0);
    signal  gt31_drpdi_i                    : std_logic_vector(15 downto 0);
    signal  gt31_drpdo_i                    : std_logic_vector(15 downto 0);
    signal  gt31_drpen_i                    : std_logic;
    signal  gt31_drprdy_i                   : std_logic;
    signal  gt31_drpwe_i                    : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt31_eyescanreset_i             : std_logic;
    signal  gt31_rxuserrdy_i                : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt31_eyescandataerror_i         : std_logic;
    signal  gt31_eyescantrigger_i           : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt31_rxslide_i                  : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt31_dmonitorout_i              : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt31_rxdata_i                   : std_logic_vector(63 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt31_rxdisperr_i                : std_logic_vector(7 downto 0);
    signal  gt31_rxnotintable_i             : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt31_gthrxn_i                   : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt31_rxdlyen_i                  : std_logic;
    signal  gt31_rxdlysreset_i              : std_logic;
    signal  gt31_rxdlysresetdone_i          : std_logic;
    signal  gt31_rxphalign_i                : std_logic;
    signal  gt31_rxphaligndone_i            : std_logic;
    signal  gt31_rxphalignen_i              : std_logic;
    signal  gt31_rxphdlyreset_i             : std_logic;
    signal  gt31_rxphmonitor_i              : std_logic_vector(4 downto 0);
    signal  gt31_rxphslipmonitor_i          : std_logic_vector(4 downto 0);
    signal  gt31_rxsyncallin_i              : std_logic;
    signal  gt31_rxsyncdone_i               : std_logic;
    signal  gt31_rxsyncin_i                 : std_logic;
    signal  gt31_rxsyncmode_i               : std_logic;
    signal  gt31_rxsyncout_i                : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt31_rxbyteisaligned_i          : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt31_rxlpmhfhold_i              : std_logic;
    signal  gt31_rxlpmlfhold_i              : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt31_rxmonitorout_i             : std_logic_vector(6 downto 0);
    signal  gt31_rxmonitorsel_i             : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt31_rxoutclk_i                 : std_logic;
    signal  gt31_rxoutclkfabric_i           : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt31_gtrxreset_i                : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt31_rxcharisk_i                : std_logic_vector(7 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt31_gthrxp_i                   : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt31_rxresetdone_i              : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt31_gttxreset_i                : std_logic;
    signal  gt31_txuserrdy_i                : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt31_txdlyen_i                  : std_logic;
    signal  gt31_txdlysreset_i              : std_logic;
    signal  gt31_txdlysresetdone_i          : std_logic;
    signal  gt31_txphalign_i                : std_logic;
    signal  gt31_txphaligndone_i            : std_logic;
    signal  gt31_txphalignen_i              : std_logic;
    signal  gt31_txphdlyreset_i             : std_logic;
    signal  gt31_txphinit_i                 : std_logic;
    signal  gt31_txphinitdone_i             : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt31_txdata_i                   : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt31_gthtxn_i                   : std_logic;
    signal  gt31_gthtxp_i                   : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt31_txoutclk_i                 : std_logic;
    signal  gt31_txoutclkfabric_i           : std_logic;
    signal  gt31_txoutclkpcs_i              : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt31_txresetdone_i              : std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt31_txcharisk_i                : std_logic_vector(7 downto 0);

    --____________________________COMMON PORTS________________________________
    signal gt0_qplllock_i : std_logic;
    signal gt0_qpllrefclklost_i  : std_logic;
    signal gt0_qpllreset_i  : std_logic;
    signal gt0_qpllreset_t  : std_logic;
     signal gt0_qplloutclk_i  : std_logic;
     signal gt0_qplloutrefclk_i : std_logic;
    --____________________________COMMON PORTS________________________________
    signal gt1_qplllock_i : std_logic;
    signal gt1_qpllrefclklost_i  : std_logic;
    signal gt1_qpllreset_i  : std_logic;
    signal gt1_qpllreset_t  : std_logic;
     signal gt1_qplloutclk_i  : std_logic;
     signal gt1_qplloutrefclk_i : std_logic;
    --____________________________COMMON PORTS________________________________
    signal gt2_qplllock_i : std_logic;
    signal gt2_qpllrefclklost_i  : std_logic;
    signal gt2_qpllreset_i  : std_logic;
    signal gt2_qpllreset_t  : std_logic;
     signal gt2_qplloutclk_i  : std_logic;
     signal gt2_qplloutrefclk_i : std_logic;
    --____________________________COMMON PORTS________________________________
    signal gt3_qplllock_i : std_logic;
    signal gt3_qpllrefclklost_i  : std_logic;
    signal gt3_qpllreset_i  : std_logic;
    signal gt3_qpllreset_t  : std_logic;
     signal gt3_qplloutclk_i  : std_logic;
     signal gt3_qplloutrefclk_i : std_logic;
    --____________________________COMMON PORTS________________________________
    signal gt4_qplllock_i : std_logic;
    signal gt4_qpllrefclklost_i  : std_logic;
    signal gt4_qpllreset_i  : std_logic;
    signal gt4_qpllreset_t  : std_logic;
     signal gt4_qplloutclk_i  : std_logic;
     signal gt4_qplloutrefclk_i : std_logic;
    --____________________________COMMON PORTS________________________________
    signal gt5_qplllock_i : std_logic;
    signal gt5_qpllrefclklost_i  : std_logic;
    signal gt5_qpllreset_i  : std_logic;
    signal gt5_qpllreset_t  : std_logic;
     signal gt5_qplloutclk_i  : std_logic;
     signal gt5_qplloutrefclk_i : std_logic;
    --____________________________COMMON PORTS________________________________
    signal gt6_qplllock_i : std_logic;
    signal gt6_qpllrefclklost_i  : std_logic;
    signal gt6_qpllreset_i  : std_logic;
    signal gt6_qpllreset_t  : std_logic;
     signal gt6_qplloutclk_i  : std_logic;
     signal gt6_qplloutrefclk_i : std_logic;
    --____________________________COMMON PORTS________________________________
    signal gt7_qplllock_i : std_logic;
    signal gt7_qpllrefclklost_i  : std_logic;
    signal gt7_qpllreset_i  : std_logic;
    signal gt7_qpllreset_t  : std_logic;
     signal gt7_qplloutclk_i  : std_logic;
     signal gt7_qplloutrefclk_i : std_logic;

    ------------------------------- Global Signals -----------------------------
    signal  gt0_tx_system_reset_c           : std_logic;
    signal  gt0_rx_system_reset_c           : std_logic;
    signal  gt1_tx_system_reset_c           : std_logic;
    signal  gt1_rx_system_reset_c           : std_logic;
    signal  gt2_tx_system_reset_c           : std_logic;
    signal  gt2_rx_system_reset_c           : std_logic;
    signal  gt3_tx_system_reset_c           : std_logic;
    signal  gt3_rx_system_reset_c           : std_logic;
    signal  gt4_tx_system_reset_c           : std_logic;
    signal  gt4_rx_system_reset_c           : std_logic;
    signal  gt5_tx_system_reset_c           : std_logic;
    signal  gt5_rx_system_reset_c           : std_logic;
    signal  gt6_tx_system_reset_c           : std_logic;
    signal  gt6_rx_system_reset_c           : std_logic;
    signal  gt7_tx_system_reset_c           : std_logic;
    signal  gt7_rx_system_reset_c           : std_logic;
    signal  gt8_tx_system_reset_c           : std_logic;
    signal  gt8_rx_system_reset_c           : std_logic;
    signal  gt9_tx_system_reset_c           : std_logic;
    signal  gt9_rx_system_reset_c           : std_logic;
    signal  gt10_tx_system_reset_c          : std_logic;
    signal  gt10_rx_system_reset_c          : std_logic;
    signal  gt11_tx_system_reset_c          : std_logic;
    signal  gt11_rx_system_reset_c          : std_logic;
    signal  gt12_tx_system_reset_c          : std_logic;
    signal  gt12_rx_system_reset_c          : std_logic;
    signal  gt13_tx_system_reset_c          : std_logic;
    signal  gt13_rx_system_reset_c          : std_logic;
    signal  gt14_tx_system_reset_c          : std_logic;
    signal  gt14_rx_system_reset_c          : std_logic;
    signal  gt15_tx_system_reset_c          : std_logic;
    signal  gt15_rx_system_reset_c          : std_logic;
    signal  gt16_tx_system_reset_c          : std_logic;
    signal  gt16_rx_system_reset_c          : std_logic;
    signal  gt17_tx_system_reset_c          : std_logic;
    signal  gt17_rx_system_reset_c          : std_logic;
    signal  gt18_tx_system_reset_c          : std_logic;
    signal  gt18_rx_system_reset_c          : std_logic;
    signal  gt19_tx_system_reset_c          : std_logic;
    signal  gt19_rx_system_reset_c          : std_logic;
    signal  gt20_tx_system_reset_c          : std_logic;
    signal  gt20_rx_system_reset_c          : std_logic;
    signal  gt21_tx_system_reset_c          : std_logic;
    signal  gt21_rx_system_reset_c          : std_logic;
    signal  gt22_tx_system_reset_c          : std_logic;
    signal  gt22_rx_system_reset_c          : std_logic;
    signal  gt23_tx_system_reset_c          : std_logic;
    signal  gt23_rx_system_reset_c          : std_logic;
    signal  gt24_tx_system_reset_c          : std_logic;
    signal  gt24_rx_system_reset_c          : std_logic;
    signal  gt25_tx_system_reset_c          : std_logic;
    signal  gt25_rx_system_reset_c          : std_logic;
    signal  gt26_tx_system_reset_c          : std_logic;
    signal  gt26_rx_system_reset_c          : std_logic;
    signal  gt27_tx_system_reset_c          : std_logic;
    signal  gt27_rx_system_reset_c          : std_logic;
    signal  gt28_tx_system_reset_c          : std_logic;
    signal  gt28_rx_system_reset_c          : std_logic;
    signal  gt29_tx_system_reset_c          : std_logic;
    signal  gt29_rx_system_reset_c          : std_logic;
    signal  gt30_tx_system_reset_c          : std_logic;
    signal  gt30_rx_system_reset_c          : std_logic;
    signal  gt31_tx_system_reset_c          : std_logic;
    signal  gt31_rx_system_reset_c          : std_logic;
    signal  tied_to_ground_i                : std_logic;
    signal  tied_to_ground_vec_i            : std_logic_vector(63 downto 0);
    signal  tied_to_vcc_i                   : std_logic;
    signal  tied_to_vcc_vec_i               : std_logic_vector(7 downto 0);
    signal  drpclk_in_i                     : std_logic;
    signal  sysclk_in_i                     : std_logic;
    signal  GTTXRESET_IN                    : std_logic;
    signal  GTRXRESET_IN                    : std_logic;
    signal  QPLLRESET_IN                    : std_logic;

    attribute keep: string;
   ------------------------------- User Clocks ---------------------------------
    signal    gt0_txusrclk_i                  : std_logic; 
    signal    gt0_txusrclk2_i                 : std_logic; 
    signal    gt0_rxusrclk_i                  : std_logic; 
    signal    gt0_rxusrclk2_i                 : std_logic; 
    
    
    
    
    signal    gt1_txusrclk_i                  : std_logic; 
    signal    gt1_txusrclk2_i                 : std_logic; 
    signal    gt1_rxusrclk_i                  : std_logic; 
    signal    gt1_rxusrclk2_i                 : std_logic; 
    
    
    
    
    signal    gt2_txusrclk_i                  : std_logic; 
    signal    gt2_txusrclk2_i                 : std_logic; 
    signal    gt2_rxusrclk_i                  : std_logic; 
    signal    gt2_rxusrclk2_i                 : std_logic; 
    
    
    
    
    signal    gt3_txusrclk_i                  : std_logic; 
    signal    gt3_txusrclk2_i                 : std_logic; 
    signal    gt3_rxusrclk_i                  : std_logic; 
    signal    gt3_rxusrclk2_i                 : std_logic; 
    
    
    
    
    signal    gt4_txusrclk_i                  : std_logic; 
    signal    gt4_txusrclk2_i                 : std_logic; 
    signal    gt4_rxusrclk_i                  : std_logic; 
    signal    gt4_rxusrclk2_i                 : std_logic; 
    
    
    
    
    signal    gt5_txusrclk_i                  : std_logic; 
    signal    gt5_txusrclk2_i                 : std_logic; 
    signal    gt5_rxusrclk_i                  : std_logic; 
    signal    gt5_rxusrclk2_i                 : std_logic; 
    
    
    
    
    signal    gt6_txusrclk_i                  : std_logic; 
    signal    gt6_txusrclk2_i                 : std_logic; 
    signal    gt6_rxusrclk_i                  : std_logic; 
    signal    gt6_rxusrclk2_i                 : std_logic; 
    
    
    
    
    signal    gt7_txusrclk_i                  : std_logic; 
    signal    gt7_txusrclk2_i                 : std_logic; 
    signal    gt7_rxusrclk_i                  : std_logic; 
    signal    gt7_rxusrclk2_i                 : std_logic; 
    
    
    
    
    signal    gt8_txusrclk_i                  : std_logic; 
    signal    gt8_txusrclk2_i                 : std_logic; 
    signal    gt8_rxusrclk_i                  : std_logic; 
    signal    gt8_rxusrclk2_i                 : std_logic; 
    
    
    
    
    signal    gt9_txusrclk_i                  : std_logic; 
    signal    gt9_txusrclk2_i                 : std_logic; 
    signal    gt9_rxusrclk_i                  : std_logic; 
    signal    gt9_rxusrclk2_i                 : std_logic; 
    
    
    
    
    signal    gt10_txusrclk_i                 : std_logic; 
    signal    gt10_txusrclk2_i                : std_logic; 
    signal    gt10_rxusrclk_i                 : std_logic; 
    signal    gt10_rxusrclk2_i                : std_logic; 
    
    
    
    
    signal    gt11_txusrclk_i                 : std_logic; 
    signal    gt11_txusrclk2_i                : std_logic; 
    signal    gt11_rxusrclk_i                 : std_logic; 
    signal    gt11_rxusrclk2_i                : std_logic; 
    
    
    
    
    signal    gt12_txusrclk_i                 : std_logic; 
    signal    gt12_txusrclk2_i                : std_logic; 
    signal    gt12_rxusrclk_i                 : std_logic; 
    signal    gt12_rxusrclk2_i                : std_logic; 
    
    
    
    
    signal    gt13_txusrclk_i                 : std_logic; 
    signal    gt13_txusrclk2_i                : std_logic; 
    signal    gt13_rxusrclk_i                 : std_logic; 
    signal    gt13_rxusrclk2_i                : std_logic; 
    
    
    
    
    signal    gt14_txusrclk_i                 : std_logic; 
    signal    gt14_txusrclk2_i                : std_logic; 
    signal    gt14_rxusrclk_i                 : std_logic; 
    signal    gt14_rxusrclk2_i                : std_logic; 
    
    
    
    
    signal    gt15_txusrclk_i                 : std_logic; 
    signal    gt15_txusrclk2_i                : std_logic; 
    signal    gt15_rxusrclk_i                 : std_logic; 
    signal    gt15_rxusrclk2_i                : std_logic; 
    
    
    
    
    signal    gt16_txusrclk_i                 : std_logic; 
    signal    gt16_txusrclk2_i                : std_logic; 
    signal    gt16_rxusrclk_i                 : std_logic; 
    signal    gt16_rxusrclk2_i                : std_logic; 
    
    
    
    
    signal    gt17_txusrclk_i                 : std_logic; 
    signal    gt17_txusrclk2_i                : std_logic; 
    signal    gt17_rxusrclk_i                 : std_logic; 
    signal    gt17_rxusrclk2_i                : std_logic; 
    
    
    
    
    signal    gt18_txusrclk_i                 : std_logic; 
    signal    gt18_txusrclk2_i                : std_logic; 
    signal    gt18_rxusrclk_i                 : std_logic; 
    signal    gt18_rxusrclk2_i                : std_logic; 
    
    
    
    
    signal    gt19_txusrclk_i                 : std_logic; 
    signal    gt19_txusrclk2_i                : std_logic; 
    signal    gt19_rxusrclk_i                 : std_logic; 
    signal    gt19_rxusrclk2_i                : std_logic; 
    
    
    
    
    signal    gt20_txusrclk_i                 : std_logic; 
    signal    gt20_txusrclk2_i                : std_logic; 
    signal    gt20_rxusrclk_i                 : std_logic; 
    signal    gt20_rxusrclk2_i                : std_logic; 
    
    
    
    
    signal    gt21_txusrclk_i                 : std_logic; 
    signal    gt21_txusrclk2_i                : std_logic; 
    signal    gt21_rxusrclk_i                 : std_logic; 
    signal    gt21_rxusrclk2_i                : std_logic; 
    
    
    
    
    signal    gt22_txusrclk_i                 : std_logic; 
    signal    gt22_txusrclk2_i                : std_logic; 
    signal    gt22_rxusrclk_i                 : std_logic; 
    signal    gt22_rxusrclk2_i                : std_logic; 
    
    
    
    
    signal    gt23_txusrclk_i                 : std_logic; 
    signal    gt23_txusrclk2_i                : std_logic; 
    signal    gt23_rxusrclk_i                 : std_logic; 
    signal    gt23_rxusrclk2_i                : std_logic; 
    
    
    
    
    signal    gt24_txusrclk_i                 : std_logic; 
    signal    gt24_txusrclk2_i                : std_logic; 
    signal    gt24_rxusrclk_i                 : std_logic; 
    signal    gt24_rxusrclk2_i                : std_logic; 
    
    
    
    
    signal    gt25_txusrclk_i                 : std_logic; 
    signal    gt25_txusrclk2_i                : std_logic; 
    signal    gt25_rxusrclk_i                 : std_logic; 
    signal    gt25_rxusrclk2_i                : std_logic; 
    
    
    
    
    signal    gt26_txusrclk_i                 : std_logic; 
    signal    gt26_txusrclk2_i                : std_logic; 
    signal    gt26_rxusrclk_i                 : std_logic; 
    signal    gt26_rxusrclk2_i                : std_logic; 
    
    
    
    
    signal    gt27_txusrclk_i                 : std_logic; 
    signal    gt27_txusrclk2_i                : std_logic; 
    signal    gt27_rxusrclk_i                 : std_logic; 
    signal    gt27_rxusrclk2_i                : std_logic; 
    
    
    
    
    signal    gt28_txusrclk_i                 : std_logic; 
    signal    gt28_txusrclk2_i                : std_logic; 
    signal    gt28_rxusrclk_i                 : std_logic; 
    signal    gt28_rxusrclk2_i                : std_logic; 
    
    
    
    
    signal    gt29_txusrclk_i                 : std_logic; 
    signal    gt29_txusrclk2_i                : std_logic; 
    signal    gt29_rxusrclk_i                 : std_logic; 
    signal    gt29_rxusrclk2_i                : std_logic; 
    
    
    
    
    signal    gt30_txusrclk_i                 : std_logic; 
    signal    gt30_txusrclk2_i                : std_logic; 
    signal    gt30_rxusrclk_i                 : std_logic; 
    signal    gt30_rxusrclk2_i                : std_logic; 
    
    
    
    
    signal    gt31_txusrclk_i                 : std_logic; 
    signal    gt31_txusrclk2_i                : std_logic; 
    signal    gt31_rxusrclk_i                 : std_logic; 
    signal    gt31_rxusrclk2_i                : std_logic; 
    
    
    
    
    signal    gt0_txmmcm_lock_i               : std_logic;
    signal    gt0_txmmcm_reset_i              : std_logic;
    signal    gt0_rxmmcm_lock_i               : std_logic; 
    signal    gt0_rxmmcm_reset_i              : std_logic;
    signal    gt1_txmmcm_lock_i               : std_logic;
    signal    gt1_txmmcm_reset_i              : std_logic;
    signal    gt1_rxmmcm_lock_i               : std_logic; 
    signal    gt1_rxmmcm_reset_i              : std_logic;
    signal    gt2_txmmcm_lock_i               : std_logic;
    signal    gt2_txmmcm_reset_i              : std_logic;
    signal    gt2_rxmmcm_lock_i               : std_logic; 
    signal    gt2_rxmmcm_reset_i              : std_logic;
    signal    gt3_txmmcm_lock_i               : std_logic;
    signal    gt3_txmmcm_reset_i              : std_logic;
    signal    gt3_rxmmcm_lock_i               : std_logic; 
    signal    gt3_rxmmcm_reset_i              : std_logic;
    signal    gt4_txmmcm_lock_i               : std_logic;
    signal    gt4_txmmcm_reset_i              : std_logic;
    signal    gt4_rxmmcm_lock_i               : std_logic; 
    signal    gt4_rxmmcm_reset_i              : std_logic;
    signal    gt5_txmmcm_lock_i               : std_logic;
    signal    gt5_txmmcm_reset_i              : std_logic;
    signal    gt5_rxmmcm_lock_i               : std_logic; 
    signal    gt5_rxmmcm_reset_i              : std_logic;
    signal    gt6_txmmcm_lock_i               : std_logic;
    signal    gt6_txmmcm_reset_i              : std_logic;
    signal    gt6_rxmmcm_lock_i               : std_logic; 
    signal    gt6_rxmmcm_reset_i              : std_logic;
    signal    gt7_txmmcm_lock_i               : std_logic;
    signal    gt7_txmmcm_reset_i              : std_logic;
    signal    gt7_rxmmcm_lock_i               : std_logic; 
    signal    gt7_rxmmcm_reset_i              : std_logic;
    signal    gt8_txmmcm_lock_i               : std_logic;
    signal    gt8_txmmcm_reset_i              : std_logic;
    signal    gt8_rxmmcm_lock_i               : std_logic; 
    signal    gt8_rxmmcm_reset_i              : std_logic;
    signal    gt9_txmmcm_lock_i               : std_logic;
    signal    gt9_txmmcm_reset_i              : std_logic;
    signal    gt9_rxmmcm_lock_i               : std_logic; 
    signal    gt9_rxmmcm_reset_i              : std_logic;
    signal    gt10_txmmcm_lock_i              : std_logic;
    signal    gt10_txmmcm_reset_i             : std_logic;
    signal    gt10_rxmmcm_lock_i              : std_logic; 
    signal    gt10_rxmmcm_reset_i             : std_logic;
    signal    gt11_txmmcm_lock_i              : std_logic;
    signal    gt11_txmmcm_reset_i             : std_logic;
    signal    gt11_rxmmcm_lock_i              : std_logic; 
    signal    gt11_rxmmcm_reset_i             : std_logic;
    signal    gt12_txmmcm_lock_i              : std_logic;
    signal    gt12_txmmcm_reset_i             : std_logic;
    signal    gt12_rxmmcm_lock_i              : std_logic; 
    signal    gt12_rxmmcm_reset_i             : std_logic;
    signal    gt13_txmmcm_lock_i              : std_logic;
    signal    gt13_txmmcm_reset_i             : std_logic;
    signal    gt13_rxmmcm_lock_i              : std_logic; 
    signal    gt13_rxmmcm_reset_i             : std_logic;
    signal    gt14_txmmcm_lock_i              : std_logic;
    signal    gt14_txmmcm_reset_i             : std_logic;
    signal    gt14_rxmmcm_lock_i              : std_logic; 
    signal    gt14_rxmmcm_reset_i             : std_logic;
    signal    gt15_txmmcm_lock_i              : std_logic;
    signal    gt15_txmmcm_reset_i             : std_logic;
    signal    gt15_rxmmcm_lock_i              : std_logic; 
    signal    gt15_rxmmcm_reset_i             : std_logic;
    signal    gt16_txmmcm_lock_i              : std_logic;
    signal    gt16_txmmcm_reset_i             : std_logic;
    signal    gt16_rxmmcm_lock_i              : std_logic; 
    signal    gt16_rxmmcm_reset_i             : std_logic;
    signal    gt17_txmmcm_lock_i              : std_logic;
    signal    gt17_txmmcm_reset_i             : std_logic;
    signal    gt17_rxmmcm_lock_i              : std_logic; 
    signal    gt17_rxmmcm_reset_i             : std_logic;
    signal    gt18_txmmcm_lock_i              : std_logic;
    signal    gt18_txmmcm_reset_i             : std_logic;
    signal    gt18_rxmmcm_lock_i              : std_logic; 
    signal    gt18_rxmmcm_reset_i             : std_logic;
    signal    gt19_txmmcm_lock_i              : std_logic;
    signal    gt19_txmmcm_reset_i             : std_logic;
    signal    gt19_rxmmcm_lock_i              : std_logic; 
    signal    gt19_rxmmcm_reset_i             : std_logic;
    signal    gt20_txmmcm_lock_i              : std_logic;
    signal    gt20_txmmcm_reset_i             : std_logic;
    signal    gt20_rxmmcm_lock_i              : std_logic; 
    signal    gt20_rxmmcm_reset_i             : std_logic;
    signal    gt21_txmmcm_lock_i              : std_logic;
    signal    gt21_txmmcm_reset_i             : std_logic;
    signal    gt21_rxmmcm_lock_i              : std_logic; 
    signal    gt21_rxmmcm_reset_i             : std_logic;
    signal    gt22_txmmcm_lock_i              : std_logic;
    signal    gt22_txmmcm_reset_i             : std_logic;
    signal    gt22_rxmmcm_lock_i              : std_logic; 
    signal    gt22_rxmmcm_reset_i             : std_logic;
    signal    gt23_txmmcm_lock_i              : std_logic;
    signal    gt23_txmmcm_reset_i             : std_logic;
    signal    gt23_rxmmcm_lock_i              : std_logic; 
    signal    gt23_rxmmcm_reset_i             : std_logic;
    signal    gt24_txmmcm_lock_i              : std_logic;
    signal    gt24_txmmcm_reset_i             : std_logic;
    signal    gt24_rxmmcm_lock_i              : std_logic; 
    signal    gt24_rxmmcm_reset_i             : std_logic;
    signal    gt25_txmmcm_lock_i              : std_logic;
    signal    gt25_txmmcm_reset_i             : std_logic;
    signal    gt25_rxmmcm_lock_i              : std_logic; 
    signal    gt25_rxmmcm_reset_i             : std_logic;
    signal    gt26_txmmcm_lock_i              : std_logic;
    signal    gt26_txmmcm_reset_i             : std_logic;
    signal    gt26_rxmmcm_lock_i              : std_logic; 
    signal    gt26_rxmmcm_reset_i             : std_logic;
    signal    gt27_txmmcm_lock_i              : std_logic;
    signal    gt27_txmmcm_reset_i             : std_logic;
    signal    gt27_rxmmcm_lock_i              : std_logic; 
    signal    gt27_rxmmcm_reset_i             : std_logic;
    signal    gt28_txmmcm_lock_i              : std_logic;
    signal    gt28_txmmcm_reset_i             : std_logic;
    signal    gt28_rxmmcm_lock_i              : std_logic; 
    signal    gt28_rxmmcm_reset_i             : std_logic;
    signal    gt29_txmmcm_lock_i              : std_logic;
    signal    gt29_txmmcm_reset_i             : std_logic;
    signal    gt29_rxmmcm_lock_i              : std_logic; 
    signal    gt29_rxmmcm_reset_i             : std_logic;
    signal    gt30_txmmcm_lock_i              : std_logic;
    signal    gt30_txmmcm_reset_i             : std_logic;
    signal    gt30_rxmmcm_lock_i              : std_logic; 
    signal    gt30_rxmmcm_reset_i             : std_logic;
    signal    gt31_txmmcm_lock_i              : std_logic;
    signal    gt31_txmmcm_reset_i             : std_logic;
    signal    gt31_rxmmcm_lock_i              : std_logic; 
    signal    gt31_rxmmcm_reset_i             : std_logic;
    ----------------------------- Reference Clocks ----------------------------
    
signal    q2_clk0_refclk_i                : std_logic;
    
signal    q5_clk0_refclk_i                : std_logic;
    
signal    q7_clk0_refclk_i                : std_logic;

signal commonreset_i : std_logic;
--**************************** Main Body of Code *******************************
begin

    --  Static signal Assigments
tied_to_ground_i                             <= '0';
tied_to_ground_vec_i                         <= x"0000000000000000";
tied_to_vcc_i                                <= '1';
tied_to_vcc_vec_i                            <= "11111111";

     GT0_TX_MMCM_LOCK_OUT <= gt0_txmmcm_lock_i;
    GT0_RX_MMCM_LOCK_OUT <= gt0_rxmmcm_lock_i;
     GT1_TX_MMCM_LOCK_OUT <= gt1_txmmcm_lock_i;
    GT1_RX_MMCM_LOCK_OUT <= gt1_rxmmcm_lock_i;
     GT2_TX_MMCM_LOCK_OUT <= gt2_txmmcm_lock_i;
    GT2_RX_MMCM_LOCK_OUT <= gt2_rxmmcm_lock_i;
     GT3_TX_MMCM_LOCK_OUT <= gt3_txmmcm_lock_i;
    GT3_RX_MMCM_LOCK_OUT <= gt3_rxmmcm_lock_i;
     GT4_TX_MMCM_LOCK_OUT <= gt4_txmmcm_lock_i;
    GT4_RX_MMCM_LOCK_OUT <= gt4_rxmmcm_lock_i;
     GT5_TX_MMCM_LOCK_OUT <= gt5_txmmcm_lock_i;
    GT5_RX_MMCM_LOCK_OUT <= gt5_rxmmcm_lock_i;
     GT6_TX_MMCM_LOCK_OUT <= gt6_txmmcm_lock_i;
    GT6_RX_MMCM_LOCK_OUT <= gt6_rxmmcm_lock_i;
     GT7_TX_MMCM_LOCK_OUT <= gt7_txmmcm_lock_i;
    GT7_RX_MMCM_LOCK_OUT <= gt7_rxmmcm_lock_i;
     GT8_TX_MMCM_LOCK_OUT <= gt8_txmmcm_lock_i;
    GT8_RX_MMCM_LOCK_OUT <= gt8_rxmmcm_lock_i;
     GT9_TX_MMCM_LOCK_OUT <= gt9_txmmcm_lock_i;
    GT9_RX_MMCM_LOCK_OUT <= gt9_rxmmcm_lock_i;
     GT10_TX_MMCM_LOCK_OUT <= gt10_txmmcm_lock_i;
    GT10_RX_MMCM_LOCK_OUT <= gt10_rxmmcm_lock_i;
     GT11_TX_MMCM_LOCK_OUT <= gt11_txmmcm_lock_i;
    GT11_RX_MMCM_LOCK_OUT <= gt11_rxmmcm_lock_i;
     GT12_TX_MMCM_LOCK_OUT <= gt12_txmmcm_lock_i;
    GT12_RX_MMCM_LOCK_OUT <= gt12_rxmmcm_lock_i;
     GT13_TX_MMCM_LOCK_OUT <= gt13_txmmcm_lock_i;
    GT13_RX_MMCM_LOCK_OUT <= gt13_rxmmcm_lock_i;
     GT14_TX_MMCM_LOCK_OUT <= gt14_txmmcm_lock_i;
    GT14_RX_MMCM_LOCK_OUT <= gt14_rxmmcm_lock_i;
     GT15_TX_MMCM_LOCK_OUT <= gt15_txmmcm_lock_i;
    GT15_RX_MMCM_LOCK_OUT <= gt15_rxmmcm_lock_i;
     GT16_TX_MMCM_LOCK_OUT <= gt16_txmmcm_lock_i;
    GT16_RX_MMCM_LOCK_OUT <= gt16_rxmmcm_lock_i;
     GT17_TX_MMCM_LOCK_OUT <= gt17_txmmcm_lock_i;
    GT17_RX_MMCM_LOCK_OUT <= gt17_rxmmcm_lock_i;
     GT18_TX_MMCM_LOCK_OUT <= gt18_txmmcm_lock_i;
    GT18_RX_MMCM_LOCK_OUT <= gt18_rxmmcm_lock_i;
     GT19_TX_MMCM_LOCK_OUT <= gt19_txmmcm_lock_i;
    GT19_RX_MMCM_LOCK_OUT <= gt19_rxmmcm_lock_i;
     GT20_TX_MMCM_LOCK_OUT <= gt20_txmmcm_lock_i;
    GT20_RX_MMCM_LOCK_OUT <= gt20_rxmmcm_lock_i;
     GT21_TX_MMCM_LOCK_OUT <= gt21_txmmcm_lock_i;
    GT21_RX_MMCM_LOCK_OUT <= gt21_rxmmcm_lock_i;
     GT22_TX_MMCM_LOCK_OUT <= gt22_txmmcm_lock_i;
    GT22_RX_MMCM_LOCK_OUT <= gt22_rxmmcm_lock_i;
     GT23_TX_MMCM_LOCK_OUT <= gt23_txmmcm_lock_i;
    GT23_RX_MMCM_LOCK_OUT <= gt23_rxmmcm_lock_i;
     GT24_TX_MMCM_LOCK_OUT <= gt24_txmmcm_lock_i;
    GT24_RX_MMCM_LOCK_OUT <= gt24_rxmmcm_lock_i;
     GT25_TX_MMCM_LOCK_OUT <= gt25_txmmcm_lock_i;
    GT25_RX_MMCM_LOCK_OUT <= gt25_rxmmcm_lock_i;
     GT26_TX_MMCM_LOCK_OUT <= gt26_txmmcm_lock_i;
    GT26_RX_MMCM_LOCK_OUT <= gt26_rxmmcm_lock_i;
     GT27_TX_MMCM_LOCK_OUT <= gt27_txmmcm_lock_i;
    GT27_RX_MMCM_LOCK_OUT <= gt27_rxmmcm_lock_i;
     GT28_TX_MMCM_LOCK_OUT <= gt28_txmmcm_lock_i;
    GT28_RX_MMCM_LOCK_OUT <= gt28_rxmmcm_lock_i;
     GT29_TX_MMCM_LOCK_OUT <= gt29_txmmcm_lock_i;
    GT29_RX_MMCM_LOCK_OUT <= gt29_rxmmcm_lock_i;
     GT30_TX_MMCM_LOCK_OUT <= gt30_txmmcm_lock_i;
    GT30_RX_MMCM_LOCK_OUT <= gt30_rxmmcm_lock_i;
     GT31_TX_MMCM_LOCK_OUT <= gt31_txmmcm_lock_i;
    GT31_RX_MMCM_LOCK_OUT <= gt31_rxmmcm_lock_i;
 
      gt0_qplllock_out  <= gt0_qplllock_i;
      gt0_qpllrefclklost_out <= gt0_qpllrefclklost_i;
     gt0_qpllreset_t <= commonreset_i or gt0_qpllreset_i;
     gt0_qpllreset_out <= commonreset_i or gt0_qpllreset_i;
     gt0_qplloutclk_out <= gt0_qplloutclk_i;
     gt0_qplloutrefclk_out <= gt0_qplloutrefclk_i;
      gt1_qplllock_out  <= gt1_qplllock_i;
      gt1_qpllrefclklost_out <= gt1_qpllrefclklost_i;
     gt1_qpllreset_t <= commonreset_i or gt1_qpllreset_i;
     gt1_qpllreset_out <= commonreset_i or gt1_qpllreset_i;
     gt1_qplloutclk_out <= gt1_qplloutclk_i;
     gt1_qplloutrefclk_out <= gt1_qplloutrefclk_i;
      gt2_qplllock_out  <= gt2_qplllock_i;
      gt2_qpllrefclklost_out <= gt2_qpllrefclklost_i;
     gt2_qpllreset_t <= commonreset_i or gt2_qpllreset_i;
     gt2_qpllreset_out <= commonreset_i or gt2_qpllreset_i;
     gt2_qplloutclk_out <= gt2_qplloutclk_i;
     gt2_qplloutrefclk_out <= gt2_qplloutrefclk_i;
      gt3_qplllock_out  <= gt3_qplllock_i;
      gt3_qpllrefclklost_out <= gt3_qpllrefclklost_i;
     gt3_qpllreset_t <= commonreset_i or gt3_qpllreset_i;
     gt3_qpllreset_out <= commonreset_i or gt3_qpllreset_i;
     gt3_qplloutclk_out <= gt3_qplloutclk_i;
     gt3_qplloutrefclk_out <= gt3_qplloutrefclk_i;
      gt4_qplllock_out  <= gt4_qplllock_i;
      gt4_qpllrefclklost_out <= gt4_qpllrefclklost_i;
     gt4_qpllreset_t <= commonreset_i or gt4_qpllreset_i;
     gt4_qpllreset_out <= commonreset_i or gt4_qpllreset_i;
     gt4_qplloutclk_out <= gt4_qplloutclk_i;
     gt4_qplloutrefclk_out <= gt4_qplloutrefclk_i;
      gt5_qplllock_out  <= gt5_qplllock_i;
      gt5_qpllrefclklost_out <= gt5_qpllrefclklost_i;
     gt5_qpllreset_t <= commonreset_i or gt5_qpllreset_i;
     gt5_qpllreset_out <= commonreset_i or gt5_qpllreset_i;
     gt5_qplloutclk_out <= gt5_qplloutclk_i;
     gt5_qplloutrefclk_out <= gt5_qplloutrefclk_i;
      gt6_qplllock_out  <= gt6_qplllock_i;
      gt6_qpllrefclklost_out <= gt6_qpllrefclklost_i;
     gt6_qpllreset_t <= commonreset_i or gt6_qpllreset_i;
     gt6_qpllreset_out <= commonreset_i or gt6_qpllreset_i;
     gt6_qplloutclk_out <= gt6_qplloutclk_i;
     gt6_qplloutrefclk_out <= gt6_qplloutrefclk_i;
      gt7_qplllock_out  <= gt7_qplllock_i;
      gt7_qpllrefclklost_out <= gt7_qpllrefclklost_i;
     gt7_qpllreset_t <= commonreset_i or gt7_qpllreset_i;
     gt7_qpllreset_out <= commonreset_i or gt7_qpllreset_i;
     gt7_qplloutclk_out <= gt7_qplloutclk_i;
     gt7_qplloutrefclk_out <= gt7_qplloutrefclk_i;


 
      GT0_TXUSRCLK_OUT <= gt0_txusrclk_i; 
      GT0_TXUSRCLK2_OUT <= gt0_txusrclk2_i;
      GT0_RXUSRCLK_OUT <= gt0_rxusrclk_i;
      GT0_RXUSRCLK2_OUT <= gt0_rxusrclk2_i;
 
      GT1_TXUSRCLK_OUT <= gt1_txusrclk_i; 
      GT1_TXUSRCLK2_OUT <= gt1_txusrclk2_i;
      GT1_RXUSRCLK_OUT <= gt1_rxusrclk_i;
      GT1_RXUSRCLK2_OUT <= gt1_rxusrclk2_i;
 
      GT2_TXUSRCLK_OUT <= gt2_txusrclk_i; 
      GT2_TXUSRCLK2_OUT <= gt2_txusrclk2_i;
      GT2_RXUSRCLK_OUT <= gt2_rxusrclk_i;
      GT2_RXUSRCLK2_OUT <= gt2_rxusrclk2_i;
 
      GT3_TXUSRCLK_OUT <= gt3_txusrclk_i; 
      GT3_TXUSRCLK2_OUT <= gt3_txusrclk2_i;
      GT3_RXUSRCLK_OUT <= gt3_rxusrclk_i;
      GT3_RXUSRCLK2_OUT <= gt3_rxusrclk2_i;
 
      GT4_TXUSRCLK_OUT <= gt4_txusrclk_i; 
      GT4_TXUSRCLK2_OUT <= gt4_txusrclk2_i;
      GT4_RXUSRCLK_OUT <= gt4_rxusrclk_i;
      GT4_RXUSRCLK2_OUT <= gt4_rxusrclk2_i;
 
      GT5_TXUSRCLK_OUT <= gt5_txusrclk_i; 
      GT5_TXUSRCLK2_OUT <= gt5_txusrclk2_i;
      GT5_RXUSRCLK_OUT <= gt5_rxusrclk_i;
      GT5_RXUSRCLK2_OUT <= gt5_rxusrclk2_i;
 
      GT6_TXUSRCLK_OUT <= gt6_txusrclk_i; 
      GT6_TXUSRCLK2_OUT <= gt6_txusrclk2_i;
      GT6_RXUSRCLK_OUT <= gt6_rxusrclk_i;
      GT6_RXUSRCLK2_OUT <= gt6_rxusrclk2_i;
 
      GT7_TXUSRCLK_OUT <= gt7_txusrclk_i; 
      GT7_TXUSRCLK2_OUT <= gt7_txusrclk2_i;
      GT7_RXUSRCLK_OUT <= gt7_rxusrclk_i;
      GT7_RXUSRCLK2_OUT <= gt7_rxusrclk2_i;
 
      GT8_TXUSRCLK_OUT <= gt8_txusrclk_i; 
      GT8_TXUSRCLK2_OUT <= gt8_txusrclk2_i;
      GT8_RXUSRCLK_OUT <= gt8_rxusrclk_i;
      GT8_RXUSRCLK2_OUT <= gt8_rxusrclk2_i;
 
      GT9_TXUSRCLK_OUT <= gt9_txusrclk_i; 
      GT9_TXUSRCLK2_OUT <= gt9_txusrclk2_i;
      GT9_RXUSRCLK_OUT <= gt9_rxusrclk_i;
      GT9_RXUSRCLK2_OUT <= gt9_rxusrclk2_i;
 
      GT10_TXUSRCLK_OUT <= gt10_txusrclk_i; 
      GT10_TXUSRCLK2_OUT <= gt10_txusrclk2_i;
      GT10_RXUSRCLK_OUT <= gt10_rxusrclk_i;
      GT10_RXUSRCLK2_OUT <= gt10_rxusrclk2_i;
 
      GT11_TXUSRCLK_OUT <= gt11_txusrclk_i; 
      GT11_TXUSRCLK2_OUT <= gt11_txusrclk2_i;
      GT11_RXUSRCLK_OUT <= gt11_rxusrclk_i;
      GT11_RXUSRCLK2_OUT <= gt11_rxusrclk2_i;
 
      GT12_TXUSRCLK_OUT <= gt12_txusrclk_i; 
      GT12_TXUSRCLK2_OUT <= gt12_txusrclk2_i;
      GT12_RXUSRCLK_OUT <= gt12_rxusrclk_i;
      GT12_RXUSRCLK2_OUT <= gt12_rxusrclk2_i;
 
      GT13_TXUSRCLK_OUT <= gt13_txusrclk_i; 
      GT13_TXUSRCLK2_OUT <= gt13_txusrclk2_i;
      GT13_RXUSRCLK_OUT <= gt13_rxusrclk_i;
      GT13_RXUSRCLK2_OUT <= gt13_rxusrclk2_i;
 
      GT14_TXUSRCLK_OUT <= gt14_txusrclk_i; 
      GT14_TXUSRCLK2_OUT <= gt14_txusrclk2_i;
      GT14_RXUSRCLK_OUT <= gt14_rxusrclk_i;
      GT14_RXUSRCLK2_OUT <= gt14_rxusrclk2_i;
 
      GT15_TXUSRCLK_OUT <= gt15_txusrclk_i; 
      GT15_TXUSRCLK2_OUT <= gt15_txusrclk2_i;
      GT15_RXUSRCLK_OUT <= gt15_rxusrclk_i;
      GT15_RXUSRCLK2_OUT <= gt15_rxusrclk2_i;
 
      GT16_TXUSRCLK_OUT <= gt16_txusrclk_i; 
      GT16_TXUSRCLK2_OUT <= gt16_txusrclk2_i;
      GT16_RXUSRCLK_OUT <= gt16_rxusrclk_i;
      GT16_RXUSRCLK2_OUT <= gt16_rxusrclk2_i;
 
      GT17_TXUSRCLK_OUT <= gt17_txusrclk_i; 
      GT17_TXUSRCLK2_OUT <= gt17_txusrclk2_i;
      GT17_RXUSRCLK_OUT <= gt17_rxusrclk_i;
      GT17_RXUSRCLK2_OUT <= gt17_rxusrclk2_i;
 
      GT18_TXUSRCLK_OUT <= gt18_txusrclk_i; 
      GT18_TXUSRCLK2_OUT <= gt18_txusrclk2_i;
      GT18_RXUSRCLK_OUT <= gt18_rxusrclk_i;
      GT18_RXUSRCLK2_OUT <= gt18_rxusrclk2_i;
 
      GT19_TXUSRCLK_OUT <= gt19_txusrclk_i; 
      GT19_TXUSRCLK2_OUT <= gt19_txusrclk2_i;
      GT19_RXUSRCLK_OUT <= gt19_rxusrclk_i;
      GT19_RXUSRCLK2_OUT <= gt19_rxusrclk2_i;
 
      GT20_TXUSRCLK_OUT <= gt20_txusrclk_i; 
      GT20_TXUSRCLK2_OUT <= gt20_txusrclk2_i;
      GT20_RXUSRCLK_OUT <= gt20_rxusrclk_i;
      GT20_RXUSRCLK2_OUT <= gt20_rxusrclk2_i;
 
      GT21_TXUSRCLK_OUT <= gt21_txusrclk_i; 
      GT21_TXUSRCLK2_OUT <= gt21_txusrclk2_i;
      GT21_RXUSRCLK_OUT <= gt21_rxusrclk_i;
      GT21_RXUSRCLK2_OUT <= gt21_rxusrclk2_i;
 
      GT22_TXUSRCLK_OUT <= gt22_txusrclk_i; 
      GT22_TXUSRCLK2_OUT <= gt22_txusrclk2_i;
      GT22_RXUSRCLK_OUT <= gt22_rxusrclk_i;
      GT22_RXUSRCLK2_OUT <= gt22_rxusrclk2_i;
 
      GT23_TXUSRCLK_OUT <= gt23_txusrclk_i; 
      GT23_TXUSRCLK2_OUT <= gt23_txusrclk2_i;
      GT23_RXUSRCLK_OUT <= gt23_rxusrclk_i;
      GT23_RXUSRCLK2_OUT <= gt23_rxusrclk2_i;
 
      GT24_TXUSRCLK_OUT <= gt24_txusrclk_i; 
      GT24_TXUSRCLK2_OUT <= gt24_txusrclk2_i;
      GT24_RXUSRCLK_OUT <= gt24_rxusrclk_i;
      GT24_RXUSRCLK2_OUT <= gt24_rxusrclk2_i;
 
      GT25_TXUSRCLK_OUT <= gt25_txusrclk_i; 
      GT25_TXUSRCLK2_OUT <= gt25_txusrclk2_i;
      GT25_RXUSRCLK_OUT <= gt25_rxusrclk_i;
      GT25_RXUSRCLK2_OUT <= gt25_rxusrclk2_i;
 
      GT26_TXUSRCLK_OUT <= gt26_txusrclk_i; 
      GT26_TXUSRCLK2_OUT <= gt26_txusrclk2_i;
      GT26_RXUSRCLK_OUT <= gt26_rxusrclk_i;
      GT26_RXUSRCLK2_OUT <= gt26_rxusrclk2_i;
 
      GT27_TXUSRCLK_OUT <= gt27_txusrclk_i; 
      GT27_TXUSRCLK2_OUT <= gt27_txusrclk2_i;
      GT27_RXUSRCLK_OUT <= gt27_rxusrclk_i;
      GT27_RXUSRCLK2_OUT <= gt27_rxusrclk2_i;
 
      GT28_TXUSRCLK_OUT <= gt28_txusrclk_i; 
      GT28_TXUSRCLK2_OUT <= gt28_txusrclk2_i;
      GT28_RXUSRCLK_OUT <= gt28_rxusrclk_i;
      GT28_RXUSRCLK2_OUT <= gt28_rxusrclk2_i;
 
      GT29_TXUSRCLK_OUT <= gt29_txusrclk_i; 
      GT29_TXUSRCLK2_OUT <= gt29_txusrclk2_i;
      GT29_RXUSRCLK_OUT <= gt29_rxusrclk_i;
      GT29_RXUSRCLK2_OUT <= gt29_rxusrclk2_i;
 
      GT30_TXUSRCLK_OUT <= gt30_txusrclk_i; 
      GT30_TXUSRCLK2_OUT <= gt30_txusrclk2_i;
      GT30_RXUSRCLK_OUT <= gt30_rxusrclk_i;
      GT30_RXUSRCLK2_OUT <= gt30_rxusrclk2_i;
 
      GT31_TXUSRCLK_OUT <= gt31_txusrclk_i; 
      GT31_TXUSRCLK2_OUT <= gt31_txusrclk2_i;
      GT31_RXUSRCLK_OUT <= gt31_rxusrclk_i;
      GT31_RXUSRCLK2_OUT <= gt31_rxusrclk2_i;


    
  
    
  
    
  
    
  
    
  
    
  
    
  
    
  
    
  
    
  
    
  
    
  
    
  
    
  
    
  
    
  
    
  
    
  
    
  
    
  
    
  
    
  
    
  
    
  
    
  
    
  
    
  
    
  
    
  
    
  
    
  
    
  
    gt_usrclk_source : gtwizard_0_GT_USRCLK_SOURCE
    port map
   (
    txusrclk2_in => txusrclk2_in,
    txusrclk_in => txusrclk_in,
        GT0_TXUSRCLK_OUT                =>      gt0_txusrclk_i,
        GT0_TXUSRCLK2_OUT               =>      gt0_txusrclk2_i,
        GT0_TXOUTCLK_IN                 =>      gt0_txoutclk_i,
        GT0_TXCLK_LOCK_OUT              =>      gt0_txmmcm_lock_i,
        GT0_TX_MMCM_RESET_IN            =>      gt0_txmmcm_reset_i,
        GT0_RXUSRCLK_OUT                =>      gt0_rxusrclk_i,
        GT0_RXUSRCLK2_OUT               =>      gt0_rxusrclk2_i,
        GT0_RXOUTCLK_IN                 =>      gt0_rxoutclk_i,
        GT0_RXCLK_LOCK_OUT              =>      gt0_rxmmcm_lock_i,
        GT0_RX_MMCM_RESET_IN            =>      gt0_rxmmcm_reset_i,
 
        GT1_TXUSRCLK_OUT                =>      gt1_txusrclk_i,
        GT1_TXUSRCLK2_OUT               =>      gt1_txusrclk2_i,
        GT1_TXOUTCLK_IN                 =>      gt1_txoutclk_i,
        GT1_TXCLK_LOCK_OUT              =>      gt1_txmmcm_lock_i,
        GT1_TX_MMCM_RESET_IN            =>      gt1_txmmcm_reset_i,
        GT1_RXUSRCLK_OUT                =>      gt1_rxusrclk_i,
        GT1_RXUSRCLK2_OUT               =>      gt1_rxusrclk2_i,
        GT1_RXOUTCLK_IN                 =>      gt1_rxoutclk_i,
        GT1_RXCLK_LOCK_OUT              =>      gt1_rxmmcm_lock_i,
        GT1_RX_MMCM_RESET_IN            =>      gt1_rxmmcm_reset_i,
 
        GT2_TXUSRCLK_OUT                =>      gt2_txusrclk_i,
        GT2_TXUSRCLK2_OUT               =>      gt2_txusrclk2_i,
        GT2_TXOUTCLK_IN                 =>      gt2_txoutclk_i,
        GT2_TXCLK_LOCK_OUT              =>      gt2_txmmcm_lock_i,
        GT2_TX_MMCM_RESET_IN            =>      gt2_txmmcm_reset_i,
        GT2_RXUSRCLK_OUT                =>      gt2_rxusrclk_i,
        GT2_RXUSRCLK2_OUT               =>      gt2_rxusrclk2_i,
        GT2_RXOUTCLK_IN                 =>      gt2_rxoutclk_i,
        GT2_RXCLK_LOCK_OUT              =>      gt2_rxmmcm_lock_i,
        GT2_RX_MMCM_RESET_IN            =>      gt2_rxmmcm_reset_i,
 
        GT3_TXUSRCLK_OUT                =>      gt3_txusrclk_i,
        GT3_TXUSRCLK2_OUT               =>      gt3_txusrclk2_i,
        GT3_TXOUTCLK_IN                 =>      gt3_txoutclk_i,
        GT3_TXCLK_LOCK_OUT              =>      gt3_txmmcm_lock_i,
        GT3_TX_MMCM_RESET_IN            =>      gt3_txmmcm_reset_i,
        GT3_RXUSRCLK_OUT                =>      gt3_rxusrclk_i,
        GT3_RXUSRCLK2_OUT               =>      gt3_rxusrclk2_i,
        GT3_RXOUTCLK_IN                 =>      gt3_rxoutclk_i,
        GT3_RXCLK_LOCK_OUT              =>      gt3_rxmmcm_lock_i,
        GT3_RX_MMCM_RESET_IN            =>      gt3_rxmmcm_reset_i,
 
        GT4_TXUSRCLK_OUT                =>      gt4_txusrclk_i,
        GT4_TXUSRCLK2_OUT               =>      gt4_txusrclk2_i,
        GT4_TXOUTCLK_IN                 =>      gt4_txoutclk_i,
        GT4_TXCLK_LOCK_OUT              =>      gt4_txmmcm_lock_i,
        GT4_TX_MMCM_RESET_IN            =>      gt4_txmmcm_reset_i,
        GT4_RXUSRCLK_OUT                =>      gt4_rxusrclk_i,
        GT4_RXUSRCLK2_OUT               =>      gt4_rxusrclk2_i,
        GT4_RXOUTCLK_IN                 =>      gt4_rxoutclk_i,
        GT4_RXCLK_LOCK_OUT              =>      gt4_rxmmcm_lock_i,
        GT4_RX_MMCM_RESET_IN            =>      gt4_rxmmcm_reset_i,
 
        GT5_TXUSRCLK_OUT                =>      gt5_txusrclk_i,
        GT5_TXUSRCLK2_OUT               =>      gt5_txusrclk2_i,
        GT5_TXOUTCLK_IN                 =>      gt5_txoutclk_i,
        GT5_TXCLK_LOCK_OUT              =>      gt5_txmmcm_lock_i,
        GT5_TX_MMCM_RESET_IN            =>      gt5_txmmcm_reset_i,
        GT5_RXUSRCLK_OUT                =>      gt5_rxusrclk_i,
        GT5_RXUSRCLK2_OUT               =>      gt5_rxusrclk2_i,
        GT5_RXOUTCLK_IN                 =>      gt5_rxoutclk_i,
        GT5_RXCLK_LOCK_OUT              =>      gt5_rxmmcm_lock_i,
        GT5_RX_MMCM_RESET_IN            =>      gt5_rxmmcm_reset_i,
 
        GT6_TXUSRCLK_OUT                =>      gt6_txusrclk_i,
        GT6_TXUSRCLK2_OUT               =>      gt6_txusrclk2_i,
        GT6_TXOUTCLK_IN                 =>      gt6_txoutclk_i,
        GT6_TXCLK_LOCK_OUT              =>      gt6_txmmcm_lock_i,
        GT6_TX_MMCM_RESET_IN            =>      gt6_txmmcm_reset_i,
        GT6_RXUSRCLK_OUT                =>      gt6_rxusrclk_i,
        GT6_RXUSRCLK2_OUT               =>      gt6_rxusrclk2_i,
        GT6_RXOUTCLK_IN                 =>      gt6_rxoutclk_i,
        GT6_RXCLK_LOCK_OUT              =>      gt6_rxmmcm_lock_i,
        GT6_RX_MMCM_RESET_IN            =>      gt6_rxmmcm_reset_i,
 
        GT7_TXUSRCLK_OUT                =>      gt7_txusrclk_i,
        GT7_TXUSRCLK2_OUT               =>      gt7_txusrclk2_i,
        GT7_TXOUTCLK_IN                 =>      gt7_txoutclk_i,
        GT7_TXCLK_LOCK_OUT              =>      gt7_txmmcm_lock_i,
        GT7_TX_MMCM_RESET_IN            =>      gt7_txmmcm_reset_i,
        GT7_RXUSRCLK_OUT                =>      gt7_rxusrclk_i,
        GT7_RXUSRCLK2_OUT               =>      gt7_rxusrclk2_i,
        GT7_RXOUTCLK_IN                 =>      gt7_rxoutclk_i,
        GT7_RXCLK_LOCK_OUT              =>      gt7_rxmmcm_lock_i,
        GT7_RX_MMCM_RESET_IN            =>      gt7_rxmmcm_reset_i,
 
        GT8_TXUSRCLK_OUT                =>      gt8_txusrclk_i,
        GT8_TXUSRCLK2_OUT               =>      gt8_txusrclk2_i,
        GT8_TXOUTCLK_IN                 =>      gt8_txoutclk_i,
        GT8_TXCLK_LOCK_OUT              =>      gt8_txmmcm_lock_i,
        GT8_TX_MMCM_RESET_IN            =>      gt8_txmmcm_reset_i,
        GT8_RXUSRCLK_OUT                =>      gt8_rxusrclk_i,
        GT8_RXUSRCLK2_OUT               =>      gt8_rxusrclk2_i,
        GT8_RXOUTCLK_IN                 =>      gt8_rxoutclk_i,
        GT8_RXCLK_LOCK_OUT              =>      gt8_rxmmcm_lock_i,
        GT8_RX_MMCM_RESET_IN            =>      gt8_rxmmcm_reset_i,
 
        GT9_TXUSRCLK_OUT                =>      gt9_txusrclk_i,
        GT9_TXUSRCLK2_OUT               =>      gt9_txusrclk2_i,
        GT9_TXOUTCLK_IN                 =>      gt9_txoutclk_i,
        GT9_TXCLK_LOCK_OUT              =>      gt9_txmmcm_lock_i,
        GT9_TX_MMCM_RESET_IN            =>      gt9_txmmcm_reset_i,
        GT9_RXUSRCLK_OUT                =>      gt9_rxusrclk_i,
        GT9_RXUSRCLK2_OUT               =>      gt9_rxusrclk2_i,
        GT9_RXOUTCLK_IN                 =>      gt9_rxoutclk_i,
        GT9_RXCLK_LOCK_OUT              =>      gt9_rxmmcm_lock_i,
        GT9_RX_MMCM_RESET_IN            =>      gt9_rxmmcm_reset_i,
 
        GT10_TXUSRCLK_OUT               =>      gt10_txusrclk_i,
        GT10_TXUSRCLK2_OUT              =>      gt10_txusrclk2_i,
        GT10_TXOUTCLK_IN                =>      gt10_txoutclk_i,
        GT10_TXCLK_LOCK_OUT             =>      gt10_txmmcm_lock_i,
        GT10_TX_MMCM_RESET_IN           =>      gt10_txmmcm_reset_i,
        GT10_RXUSRCLK_OUT               =>      gt10_rxusrclk_i,
        GT10_RXUSRCLK2_OUT              =>      gt10_rxusrclk2_i,
        GT10_RXOUTCLK_IN                =>      gt10_rxoutclk_i,
        GT10_RXCLK_LOCK_OUT             =>      gt10_rxmmcm_lock_i,
        GT10_RX_MMCM_RESET_IN           =>      gt10_rxmmcm_reset_i,
 
        GT11_TXUSRCLK_OUT               =>      gt11_txusrclk_i,
        GT11_TXUSRCLK2_OUT              =>      gt11_txusrclk2_i,
        GT11_TXOUTCLK_IN                =>      gt11_txoutclk_i,
        GT11_TXCLK_LOCK_OUT             =>      gt11_txmmcm_lock_i,
        GT11_TX_MMCM_RESET_IN           =>      gt11_txmmcm_reset_i,
        GT11_RXUSRCLK_OUT               =>      gt11_rxusrclk_i,
        GT11_RXUSRCLK2_OUT              =>      gt11_rxusrclk2_i,
        GT11_RXOUTCLK_IN                =>      gt11_rxoutclk_i,
        GT11_RXCLK_LOCK_OUT             =>      gt11_rxmmcm_lock_i,
        GT11_RX_MMCM_RESET_IN           =>      gt11_rxmmcm_reset_i,
 
        GT12_TXUSRCLK_OUT               =>      gt12_txusrclk_i,
        GT12_TXUSRCLK2_OUT              =>      gt12_txusrclk2_i,
        GT12_TXOUTCLK_IN                =>      gt12_txoutclk_i,
        GT12_TXCLK_LOCK_OUT             =>      gt12_txmmcm_lock_i,
        GT12_TX_MMCM_RESET_IN           =>      gt12_txmmcm_reset_i,
        GT12_RXUSRCLK_OUT               =>      gt12_rxusrclk_i,
        GT12_RXUSRCLK2_OUT              =>      gt12_rxusrclk2_i,
        GT12_RXOUTCLK_IN                =>      gt12_rxoutclk_i,
        GT12_RXCLK_LOCK_OUT             =>      gt12_rxmmcm_lock_i,
        GT12_RX_MMCM_RESET_IN           =>      gt12_rxmmcm_reset_i,
 
        GT13_TXUSRCLK_OUT               =>      gt13_txusrclk_i,
        GT13_TXUSRCLK2_OUT              =>      gt13_txusrclk2_i,
        GT13_TXOUTCLK_IN                =>      gt13_txoutclk_i,
        GT13_TXCLK_LOCK_OUT             =>      gt13_txmmcm_lock_i,
        GT13_TX_MMCM_RESET_IN           =>      gt13_txmmcm_reset_i,
        GT13_RXUSRCLK_OUT               =>      gt13_rxusrclk_i,
        GT13_RXUSRCLK2_OUT              =>      gt13_rxusrclk2_i,
        GT13_RXOUTCLK_IN                =>      gt13_rxoutclk_i,
        GT13_RXCLK_LOCK_OUT             =>      gt13_rxmmcm_lock_i,
        GT13_RX_MMCM_RESET_IN           =>      gt13_rxmmcm_reset_i,
 
        GT14_TXUSRCLK_OUT               =>      gt14_txusrclk_i,
        GT14_TXUSRCLK2_OUT              =>      gt14_txusrclk2_i,
        GT14_TXOUTCLK_IN                =>      gt14_txoutclk_i,
        GT14_TXCLK_LOCK_OUT             =>      gt14_txmmcm_lock_i,
        GT14_TX_MMCM_RESET_IN           =>      gt14_txmmcm_reset_i,
        GT14_RXUSRCLK_OUT               =>      gt14_rxusrclk_i,
        GT14_RXUSRCLK2_OUT              =>      gt14_rxusrclk2_i,
        GT14_RXOUTCLK_IN                =>      gt14_rxoutclk_i,
        GT14_RXCLK_LOCK_OUT             =>      gt14_rxmmcm_lock_i,
        GT14_RX_MMCM_RESET_IN           =>      gt14_rxmmcm_reset_i,
 
        GT15_TXUSRCLK_OUT               =>      gt15_txusrclk_i,
        GT15_TXUSRCLK2_OUT              =>      gt15_txusrclk2_i,
        GT15_TXOUTCLK_IN                =>      gt15_txoutclk_i,
        GT15_TXCLK_LOCK_OUT             =>      gt15_txmmcm_lock_i,
        GT15_TX_MMCM_RESET_IN           =>      gt15_txmmcm_reset_i,
        GT15_RXUSRCLK_OUT               =>      gt15_rxusrclk_i,
        GT15_RXUSRCLK2_OUT              =>      gt15_rxusrclk2_i,
        GT15_RXOUTCLK_IN                =>      gt15_rxoutclk_i,
        GT15_RXCLK_LOCK_OUT             =>      gt15_rxmmcm_lock_i,
        GT15_RX_MMCM_RESET_IN           =>      gt15_rxmmcm_reset_i,
 
        GT16_TXUSRCLK_OUT               =>      gt16_txusrclk_i,
        GT16_TXUSRCLK2_OUT              =>      gt16_txusrclk2_i,
        GT16_TXOUTCLK_IN                =>      gt16_txoutclk_i,
        GT16_TXCLK_LOCK_OUT             =>      gt16_txmmcm_lock_i,
        GT16_TX_MMCM_RESET_IN           =>      gt16_txmmcm_reset_i,
        GT16_RXUSRCLK_OUT               =>      gt16_rxusrclk_i,
        GT16_RXUSRCLK2_OUT              =>      gt16_rxusrclk2_i,
        GT16_RXOUTCLK_IN                =>      gt16_rxoutclk_i,
        GT16_RXCLK_LOCK_OUT             =>      gt16_rxmmcm_lock_i,
        GT16_RX_MMCM_RESET_IN           =>      gt16_rxmmcm_reset_i,
 
        GT17_TXUSRCLK_OUT               =>      gt17_txusrclk_i,
        GT17_TXUSRCLK2_OUT              =>      gt17_txusrclk2_i,
        GT17_TXOUTCLK_IN                =>      gt17_txoutclk_i,
        GT17_TXCLK_LOCK_OUT             =>      gt17_txmmcm_lock_i,
        GT17_TX_MMCM_RESET_IN           =>      gt17_txmmcm_reset_i,
        GT17_RXUSRCLK_OUT               =>      gt17_rxusrclk_i,
        GT17_RXUSRCLK2_OUT              =>      gt17_rxusrclk2_i,
        GT17_RXOUTCLK_IN                =>      gt17_rxoutclk_i,
        GT17_RXCLK_LOCK_OUT             =>      gt17_rxmmcm_lock_i,
        GT17_RX_MMCM_RESET_IN           =>      gt17_rxmmcm_reset_i,
 
        GT18_TXUSRCLK_OUT               =>      gt18_txusrclk_i,
        GT18_TXUSRCLK2_OUT              =>      gt18_txusrclk2_i,
        GT18_TXOUTCLK_IN                =>      gt18_txoutclk_i,
        GT18_TXCLK_LOCK_OUT             =>      gt18_txmmcm_lock_i,
        GT18_TX_MMCM_RESET_IN           =>      gt18_txmmcm_reset_i,
        GT18_RXUSRCLK_OUT               =>      gt18_rxusrclk_i,
        GT18_RXUSRCLK2_OUT              =>      gt18_rxusrclk2_i,
        GT18_RXOUTCLK_IN                =>      gt18_rxoutclk_i,
        GT18_RXCLK_LOCK_OUT             =>      gt18_rxmmcm_lock_i,
        GT18_RX_MMCM_RESET_IN           =>      gt18_rxmmcm_reset_i,
 
        GT19_TXUSRCLK_OUT               =>      gt19_txusrclk_i,
        GT19_TXUSRCLK2_OUT              =>      gt19_txusrclk2_i,
        GT19_TXOUTCLK_IN                =>      gt19_txoutclk_i,
        GT19_TXCLK_LOCK_OUT             =>      gt19_txmmcm_lock_i,
        GT19_TX_MMCM_RESET_IN           =>      gt19_txmmcm_reset_i,
        GT19_RXUSRCLK_OUT               =>      gt19_rxusrclk_i,
        GT19_RXUSRCLK2_OUT              =>      gt19_rxusrclk2_i,
        GT19_RXOUTCLK_IN                =>      gt19_rxoutclk_i,
        GT19_RXCLK_LOCK_OUT             =>      gt19_rxmmcm_lock_i,
        GT19_RX_MMCM_RESET_IN           =>      gt19_rxmmcm_reset_i,
 
        GT20_TXUSRCLK_OUT               =>      gt20_txusrclk_i,
        GT20_TXUSRCLK2_OUT              =>      gt20_txusrclk2_i,
        GT20_TXOUTCLK_IN                =>      gt20_txoutclk_i,
        GT20_TXCLK_LOCK_OUT             =>      gt20_txmmcm_lock_i,
        GT20_TX_MMCM_RESET_IN           =>      gt20_txmmcm_reset_i,
        GT20_RXUSRCLK_OUT               =>      gt20_rxusrclk_i,
        GT20_RXUSRCLK2_OUT              =>      gt20_rxusrclk2_i,
        GT20_RXOUTCLK_IN                =>      gt20_rxoutclk_i,
        GT20_RXCLK_LOCK_OUT             =>      gt20_rxmmcm_lock_i,
        GT20_RX_MMCM_RESET_IN           =>      gt20_rxmmcm_reset_i,
 
        GT21_TXUSRCLK_OUT               =>      gt21_txusrclk_i,
        GT21_TXUSRCLK2_OUT              =>      gt21_txusrclk2_i,
        GT21_TXOUTCLK_IN                =>      gt21_txoutclk_i,
        GT21_TXCLK_LOCK_OUT             =>      gt21_txmmcm_lock_i,
        GT21_TX_MMCM_RESET_IN           =>      gt21_txmmcm_reset_i,
        GT21_RXUSRCLK_OUT               =>      gt21_rxusrclk_i,
        GT21_RXUSRCLK2_OUT              =>      gt21_rxusrclk2_i,
        GT21_RXOUTCLK_IN                =>      gt21_rxoutclk_i,
        GT21_RXCLK_LOCK_OUT             =>      gt21_rxmmcm_lock_i,
        GT21_RX_MMCM_RESET_IN           =>      gt21_rxmmcm_reset_i,
 
        GT22_TXUSRCLK_OUT               =>      gt22_txusrclk_i,
        GT22_TXUSRCLK2_OUT              =>      gt22_txusrclk2_i,
        GT22_TXOUTCLK_IN                =>      gt22_txoutclk_i,
        GT22_TXCLK_LOCK_OUT             =>      gt22_txmmcm_lock_i,
        GT22_TX_MMCM_RESET_IN           =>      gt22_txmmcm_reset_i,
        GT22_RXUSRCLK_OUT               =>      gt22_rxusrclk_i,
        GT22_RXUSRCLK2_OUT              =>      gt22_rxusrclk2_i,
        GT22_RXOUTCLK_IN                =>      gt22_rxoutclk_i,
        GT22_RXCLK_LOCK_OUT             =>      gt22_rxmmcm_lock_i,
        GT22_RX_MMCM_RESET_IN           =>      gt22_rxmmcm_reset_i,
 
        GT23_TXUSRCLK_OUT               =>      gt23_txusrclk_i,
        GT23_TXUSRCLK2_OUT              =>      gt23_txusrclk2_i,
        GT23_TXOUTCLK_IN                =>      gt23_txoutclk_i,
        GT23_TXCLK_LOCK_OUT             =>      gt23_txmmcm_lock_i,
        GT23_TX_MMCM_RESET_IN           =>      gt23_txmmcm_reset_i,
        GT23_RXUSRCLK_OUT               =>      gt23_rxusrclk_i,
        GT23_RXUSRCLK2_OUT              =>      gt23_rxusrclk2_i,
        GT23_RXOUTCLK_IN                =>      gt23_rxoutclk_i,
        GT23_RXCLK_LOCK_OUT             =>      gt23_rxmmcm_lock_i,
        GT23_RX_MMCM_RESET_IN           =>      gt23_rxmmcm_reset_i,
 
        GT24_TXUSRCLK_OUT               =>      gt24_txusrclk_i,
        GT24_TXUSRCLK2_OUT              =>      gt24_txusrclk2_i,
        GT24_TXOUTCLK_IN                =>      gt24_txoutclk_i,
        GT24_TXCLK_LOCK_OUT             =>      gt24_txmmcm_lock_i,
        GT24_TX_MMCM_RESET_IN           =>      gt24_txmmcm_reset_i,
        GT24_RXUSRCLK_OUT               =>      gt24_rxusrclk_i,
        GT24_RXUSRCLK2_OUT              =>      gt24_rxusrclk2_i,
        GT24_RXOUTCLK_IN                =>      gt24_rxoutclk_i,
        GT24_RXCLK_LOCK_OUT             =>      gt24_rxmmcm_lock_i,
        GT24_RX_MMCM_RESET_IN           =>      gt24_rxmmcm_reset_i,
 
        GT25_TXUSRCLK_OUT               =>      gt25_txusrclk_i,
        GT25_TXUSRCLK2_OUT              =>      gt25_txusrclk2_i,
        GT25_TXOUTCLK_IN                =>      gt25_txoutclk_i,
        GT25_TXCLK_LOCK_OUT             =>      gt25_txmmcm_lock_i,
        GT25_TX_MMCM_RESET_IN           =>      gt25_txmmcm_reset_i,
        GT25_RXUSRCLK_OUT               =>      gt25_rxusrclk_i,
        GT25_RXUSRCLK2_OUT              =>      gt25_rxusrclk2_i,
        GT25_RXOUTCLK_IN                =>      gt25_rxoutclk_i,
        GT25_RXCLK_LOCK_OUT             =>      gt25_rxmmcm_lock_i,
        GT25_RX_MMCM_RESET_IN           =>      gt25_rxmmcm_reset_i,
 
        GT26_TXUSRCLK_OUT               =>      gt26_txusrclk_i,
        GT26_TXUSRCLK2_OUT              =>      gt26_txusrclk2_i,
        GT26_TXOUTCLK_IN                =>      gt26_txoutclk_i,
        GT26_TXCLK_LOCK_OUT             =>      gt26_txmmcm_lock_i,
        GT26_TX_MMCM_RESET_IN           =>      gt26_txmmcm_reset_i,
        GT26_RXUSRCLK_OUT               =>      gt26_rxusrclk_i,
        GT26_RXUSRCLK2_OUT              =>      gt26_rxusrclk2_i,
        GT26_RXOUTCLK_IN                =>      gt26_rxoutclk_i,
        GT26_RXCLK_LOCK_OUT             =>      gt26_rxmmcm_lock_i,
        GT26_RX_MMCM_RESET_IN           =>      gt26_rxmmcm_reset_i,
 
        GT27_TXUSRCLK_OUT               =>      gt27_txusrclk_i,
        GT27_TXUSRCLK2_OUT              =>      gt27_txusrclk2_i,
        GT27_TXOUTCLK_IN                =>      gt27_txoutclk_i,
        GT27_TXCLK_LOCK_OUT             =>      gt27_txmmcm_lock_i,
        GT27_TX_MMCM_RESET_IN           =>      gt27_txmmcm_reset_i,
        GT27_RXUSRCLK_OUT               =>      gt27_rxusrclk_i,
        GT27_RXUSRCLK2_OUT              =>      gt27_rxusrclk2_i,
        GT27_RXOUTCLK_IN                =>      gt27_rxoutclk_i,
        GT27_RXCLK_LOCK_OUT             =>      gt27_rxmmcm_lock_i,
        GT27_RX_MMCM_RESET_IN           =>      gt27_rxmmcm_reset_i,
 
        GT28_TXUSRCLK_OUT               =>      gt28_txusrclk_i,
        GT28_TXUSRCLK2_OUT              =>      gt28_txusrclk2_i,
        GT28_TXOUTCLK_IN                =>      gt28_txoutclk_i,
        GT28_TXCLK_LOCK_OUT             =>      gt28_txmmcm_lock_i,
        GT28_TX_MMCM_RESET_IN           =>      gt28_txmmcm_reset_i,
        GT28_RXUSRCLK_OUT               =>      gt28_rxusrclk_i,
        GT28_RXUSRCLK2_OUT              =>      gt28_rxusrclk2_i,
        GT28_RXOUTCLK_IN                =>      gt28_rxoutclk_i,
        GT28_RXCLK_LOCK_OUT             =>      gt28_rxmmcm_lock_i,
        GT28_RX_MMCM_RESET_IN           =>      gt28_rxmmcm_reset_i,
 
        GT29_TXUSRCLK_OUT               =>      gt29_txusrclk_i,
        GT29_TXUSRCLK2_OUT              =>      gt29_txusrclk2_i,
        GT29_TXOUTCLK_IN                =>      gt29_txoutclk_i,
        GT29_TXCLK_LOCK_OUT             =>      gt29_txmmcm_lock_i,
        GT29_TX_MMCM_RESET_IN           =>      gt29_txmmcm_reset_i,
        GT29_RXUSRCLK_OUT               =>      gt29_rxusrclk_i,
        GT29_RXUSRCLK2_OUT              =>      gt29_rxusrclk2_i,
        GT29_RXOUTCLK_IN                =>      gt29_rxoutclk_i,
        GT29_RXCLK_LOCK_OUT             =>      gt29_rxmmcm_lock_i,
        GT29_RX_MMCM_RESET_IN           =>      gt29_rxmmcm_reset_i,
 
        GT30_TXUSRCLK_OUT               =>      gt30_txusrclk_i,
        GT30_TXUSRCLK2_OUT              =>      gt30_txusrclk2_i,
        GT30_TXOUTCLK_IN                =>      gt30_txoutclk_i,
        GT30_TXCLK_LOCK_OUT             =>      gt30_txmmcm_lock_i,
        GT30_TX_MMCM_RESET_IN           =>      gt30_txmmcm_reset_i,
        GT30_RXUSRCLK_OUT               =>      gt30_rxusrclk_i,
        GT30_RXUSRCLK2_OUT              =>      gt30_rxusrclk2_i,
        GT30_RXOUTCLK_IN                =>      gt30_rxoutclk_i,
        GT30_RXCLK_LOCK_OUT             =>      gt30_rxmmcm_lock_i,
        GT30_RX_MMCM_RESET_IN           =>      gt30_rxmmcm_reset_i,
 
        GT31_TXUSRCLK_OUT               =>      gt31_txusrclk_i,
        GT31_TXUSRCLK2_OUT              =>      gt31_txusrclk2_i,
        GT31_TXOUTCLK_IN                =>      gt31_txoutclk_i,
        GT31_TXCLK_LOCK_OUT             =>      gt31_txmmcm_lock_i,
        GT31_TX_MMCM_RESET_IN           =>      gt31_txmmcm_reset_i,
        GT31_RXUSRCLK_OUT               =>      gt31_rxusrclk_i,
        GT31_RXUSRCLK2_OUT              =>      gt31_rxusrclk2_i,
        GT31_RXOUTCLK_IN                =>      gt31_rxoutclk_i,
        GT31_RXCLK_LOCK_OUT             =>      gt31_rxmmcm_lock_i,
        GT31_RX_MMCM_RESET_IN           =>      gt31_rxmmcm_reset_i,
        Q2_CLK0_GTREFCLK_PAD_N_IN       =>      Q2_CLK0_GTREFCLK_PAD_N_IN,
        Q2_CLK0_GTREFCLK_PAD_P_IN       =>      Q2_CLK0_GTREFCLK_PAD_P_IN,
        Q2_CLK0_GTREFCLK_OUT            =>      q2_clk0_refclk_i,
        Q5_CLK0_GTREFCLK_PAD_N_IN       =>      Q5_CLK0_GTREFCLK_PAD_N_IN,
        Q5_CLK0_GTREFCLK_PAD_P_IN       =>      Q5_CLK0_GTREFCLK_PAD_P_IN,
        Q5_CLK0_GTREFCLK_OUT            =>      q5_clk0_refclk_i,
        Q7_CLK0_GTREFCLK_PAD_N_IN       =>      Q7_CLK0_GTREFCLK_PAD_N_IN,
        Q7_CLK0_GTREFCLK_PAD_P_IN       =>      Q7_CLK0_GTREFCLK_PAD_P_IN,
        Q7_CLK0_GTREFCLK_OUT            =>      q7_clk0_refclk_i

    );

sysclk_in_i <= sysclk_in;

    common0_i:gtwizard_0_common 
  generic map
  (
   WRAPPER_SIM_GTRESET_SPEEDUP => EXAMPLE_SIM_GTRESET_SPEEDUP,
   SIM_QPLLREFCLK_SEL => "001"
  )
 port map
   (
    QPLLREFCLKSEL_IN    => "001",
    GTREFCLK0_IN      => q2_clk0_refclk_i,
    GTREFCLK1_IN      => tied_to_ground_i,
    QPLLLOCK_OUT => gt0_qplllock_i,
    QPLLLOCKDETCLK_IN => sysclk_in_i,
    QPLLOUTCLK_OUT => gt0_qplloutclk_i,
    QPLLOUTREFCLK_OUT => gt0_qplloutrefclk_i,
    QPLLREFCLKLOST_OUT => gt0_qpllrefclklost_i,    
    QPLLRESET_IN => gt0_qpllreset_t

);

    common1_i:gtwizard_0_common 
  generic map
  (
   WRAPPER_SIM_GTRESET_SPEEDUP => EXAMPLE_SIM_GTRESET_SPEEDUP,
   SIM_QPLLREFCLK_SEL => "001"
  )
 port map
   (
    QPLLREFCLKSEL_IN    => "001",
    GTREFCLK0_IN      => q2_clk0_refclk_i,
    GTREFCLK1_IN      => tied_to_ground_i,
    QPLLLOCK_OUT => gt1_qplllock_i,
    QPLLLOCKDETCLK_IN => sysclk_in_i,
    QPLLOUTCLK_OUT => gt1_qplloutclk_i,
    QPLLOUTREFCLK_OUT => gt1_qplloutrefclk_i,
    QPLLREFCLKLOST_OUT => gt1_qpllrefclklost_i,    
    QPLLRESET_IN => gt1_qpllreset_t

);

    common2_i:gtwizard_0_common 
  generic map
  (
   WRAPPER_SIM_GTRESET_SPEEDUP => EXAMPLE_SIM_GTRESET_SPEEDUP,
   SIM_QPLLREFCLK_SEL => "001"
  )
 port map
   (
    QPLLREFCLKSEL_IN    => "001",
    GTREFCLK0_IN      => q2_clk0_refclk_i,
    GTREFCLK1_IN      => tied_to_ground_i,
    QPLLLOCK_OUT => gt2_qplllock_i,
    QPLLLOCKDETCLK_IN => sysclk_in_i,
    QPLLOUTCLK_OUT => gt2_qplloutclk_i,
    QPLLOUTREFCLK_OUT => gt2_qplloutrefclk_i,
    QPLLREFCLKLOST_OUT => gt2_qpllrefclklost_i,    
    QPLLRESET_IN => gt2_qpllreset_t

);

    common3_i:gtwizard_0_common 
  generic map
  (
   WRAPPER_SIM_GTRESET_SPEEDUP => EXAMPLE_SIM_GTRESET_SPEEDUP,
   SIM_QPLLREFCLK_SEL => "001"
  )
 port map
   (
    QPLLREFCLKSEL_IN    => "001",
    GTREFCLK0_IN      => q5_clk0_refclk_i,
    GTREFCLK1_IN      => tied_to_ground_i,
    QPLLLOCK_OUT => gt3_qplllock_i,
    QPLLLOCKDETCLK_IN => sysclk_in_i,
    QPLLOUTCLK_OUT => gt3_qplloutclk_i,
    QPLLOUTREFCLK_OUT => gt3_qplloutrefclk_i,
    QPLLREFCLKLOST_OUT => gt3_qpllrefclklost_i,    
    QPLLRESET_IN => gt3_qpllreset_t

);

    common4_i:gtwizard_0_common 
  generic map
  (
   WRAPPER_SIM_GTRESET_SPEEDUP => EXAMPLE_SIM_GTRESET_SPEEDUP,
   SIM_QPLLREFCLK_SEL => "001"
  )
 port map
   (
    QPLLREFCLKSEL_IN    => "001",
    GTREFCLK0_IN      => q5_clk0_refclk_i,
    GTREFCLK1_IN      => tied_to_ground_i,
    QPLLLOCK_OUT => gt4_qplllock_i,
    QPLLLOCKDETCLK_IN => sysclk_in_i,
    QPLLOUTCLK_OUT => gt4_qplloutclk_i,
    QPLLOUTREFCLK_OUT => gt4_qplloutrefclk_i,
    QPLLREFCLKLOST_OUT => gt4_qpllrefclklost_i,    
    QPLLRESET_IN => gt4_qpllreset_t

);

    common5_i:gtwizard_0_common 
  generic map
  (
   WRAPPER_SIM_GTRESET_SPEEDUP => EXAMPLE_SIM_GTRESET_SPEEDUP,
   SIM_QPLLREFCLK_SEL => "001"
  )
 port map
   (
    QPLLREFCLKSEL_IN    => "001",
    GTREFCLK0_IN      => q5_clk0_refclk_i,
    GTREFCLK1_IN      => tied_to_ground_i,
    QPLLLOCK_OUT => gt5_qplllock_i,
    QPLLLOCKDETCLK_IN => sysclk_in_i,
    QPLLOUTCLK_OUT => gt5_qplloutclk_i,
    QPLLOUTREFCLK_OUT => gt5_qplloutrefclk_i,
    QPLLREFCLKLOST_OUT => gt5_qpllrefclklost_i,    
    QPLLRESET_IN => gt5_qpllreset_t

);

    common6_i:gtwizard_0_common 
  generic map
  (
   WRAPPER_SIM_GTRESET_SPEEDUP => EXAMPLE_SIM_GTRESET_SPEEDUP,
   SIM_QPLLREFCLK_SEL => "001"
  )
 port map
   (
    QPLLREFCLKSEL_IN    => "001",
    GTREFCLK0_IN      => q7_clk0_refclk_i,
    GTREFCLK1_IN      => tied_to_ground_i,
    QPLLLOCK_OUT => gt6_qplllock_i,
    QPLLLOCKDETCLK_IN => sysclk_in_i,
    QPLLOUTCLK_OUT => gt6_qplloutclk_i,
    QPLLOUTREFCLK_OUT => gt6_qplloutrefclk_i,
    QPLLREFCLKLOST_OUT => gt6_qpllrefclklost_i,    
    QPLLRESET_IN => gt6_qpllreset_t

);

    common7_i:gtwizard_0_common 
  generic map
  (
   WRAPPER_SIM_GTRESET_SPEEDUP => EXAMPLE_SIM_GTRESET_SPEEDUP,
   SIM_QPLLREFCLK_SEL => "001"
  )
 port map
   (
    QPLLREFCLKSEL_IN    => "001",
    GTREFCLK0_IN      => q7_clk0_refclk_i,
    GTREFCLK1_IN      => tied_to_ground_i,
    QPLLLOCK_OUT => gt7_qplllock_i,
    QPLLLOCKDETCLK_IN => sysclk_in_i,
    QPLLOUTCLK_OUT => gt7_qplloutclk_i,
    QPLLOUTREFCLK_OUT => gt7_qplloutrefclk_i,
    QPLLREFCLKLOST_OUT => gt7_qpllrefclklost_i,    
    QPLLRESET_IN => gt7_qpllreset_t

);

    common_reset_i:gtwizard_0_common_reset 
   generic map 
   (
      STABLE_CLOCK_PERIOD =>STABLE_CLOCK_PERIOD        -- Period of the stable clock driving this state-machine, unit is [ns]
   )
   port map
   (    
      STABLE_CLOCK => sysclk_in_i,             --Stable Clock, either a stable clock from the PCB
     
      SOFT_RESET => soft_reset_tx_in,               --User Reset, can be pulled any time
      COMMON_RESET => commonreset_i              --Reset QPLL
   );


    gtwizard_0_init_i : gtwizard_0_init
    port map
    (
        sysclk_in                       =>      sysclk_in_i,
        soft_reset_tx_in                =>      SOFT_RESET_TX_IN,
        soft_reset_rx_in                =>      SOFT_RESET_RX_IN,
        dont_reset_on_data_error_in     =>      DONT_RESET_ON_DATA_ERROR_IN,
        gt0_tx_mmcm_lock_in             =>      gt0_txmmcm_lock_i,
        gt0_tx_mmcm_reset_out           =>      gt0_txmmcm_reset_i,
        gt0_rx_mmcm_lock_in             =>      gt0_rxmmcm_lock_i,
        gt0_rx_mmcm_reset_out           =>      gt0_rxmmcm_reset_i,
        gt0_drp_busy_out                =>      open,
        gt0_tx_fsm_reset_done_out       =>      gt0_tx_fsm_reset_done_out,
        gt0_rx_fsm_reset_done_out       =>      gt0_rx_fsm_reset_done_out,
        gt0_data_valid_in               =>      gt0_data_valid_in,
        gt1_tx_mmcm_lock_in             =>      gt1_txmmcm_lock_i,
        gt1_tx_mmcm_reset_out           =>      gt1_txmmcm_reset_i,
        gt1_rx_mmcm_lock_in             =>      gt1_rxmmcm_lock_i,
        gt1_rx_mmcm_reset_out           =>      gt1_rxmmcm_reset_i,
        gt1_drp_busy_out                =>      open,
        gt1_tx_fsm_reset_done_out       =>      gt1_tx_fsm_reset_done_out,
        gt1_rx_fsm_reset_done_out       =>      gt1_rx_fsm_reset_done_out,
        gt1_data_valid_in               =>      gt1_data_valid_in,
        gt2_tx_mmcm_lock_in             =>      gt2_txmmcm_lock_i,
        gt2_tx_mmcm_reset_out           =>      gt2_txmmcm_reset_i,
        gt2_rx_mmcm_lock_in             =>      gt2_rxmmcm_lock_i,
        gt2_rx_mmcm_reset_out           =>      gt2_rxmmcm_reset_i,
        gt2_drp_busy_out                =>      open,
        gt2_tx_fsm_reset_done_out       =>      gt2_tx_fsm_reset_done_out,
        gt2_rx_fsm_reset_done_out       =>      gt2_rx_fsm_reset_done_out,
        gt2_data_valid_in               =>      gt2_data_valid_in,
        gt3_tx_mmcm_lock_in             =>      gt3_txmmcm_lock_i,
        gt3_tx_mmcm_reset_out           =>      gt3_txmmcm_reset_i,
        gt3_rx_mmcm_lock_in             =>      gt3_rxmmcm_lock_i,
        gt3_rx_mmcm_reset_out           =>      gt3_rxmmcm_reset_i,
        gt3_drp_busy_out                =>      open,
        gt3_tx_fsm_reset_done_out       =>      gt3_tx_fsm_reset_done_out,
        gt3_rx_fsm_reset_done_out       =>      gt3_rx_fsm_reset_done_out,
        gt3_data_valid_in               =>      gt3_data_valid_in,
        gt4_tx_mmcm_lock_in             =>      gt4_txmmcm_lock_i,
        gt4_tx_mmcm_reset_out           =>      gt4_txmmcm_reset_i,
        gt4_rx_mmcm_lock_in             =>      gt4_rxmmcm_lock_i,
        gt4_rx_mmcm_reset_out           =>      gt4_rxmmcm_reset_i,
        gt4_drp_busy_out                =>      open,
        gt4_tx_fsm_reset_done_out       =>      gt4_tx_fsm_reset_done_out,
        gt4_rx_fsm_reset_done_out       =>      gt4_rx_fsm_reset_done_out,
        gt4_data_valid_in               =>      gt4_data_valid_in,
        gt5_tx_mmcm_lock_in             =>      gt5_txmmcm_lock_i,
        gt5_tx_mmcm_reset_out           =>      gt5_txmmcm_reset_i,
        gt5_rx_mmcm_lock_in             =>      gt5_rxmmcm_lock_i,
        gt5_rx_mmcm_reset_out           =>      gt5_rxmmcm_reset_i,
        gt5_drp_busy_out                =>      open,
        gt5_tx_fsm_reset_done_out       =>      gt5_tx_fsm_reset_done_out,
        gt5_rx_fsm_reset_done_out       =>      gt5_rx_fsm_reset_done_out,
        gt5_data_valid_in               =>      gt5_data_valid_in,
        gt6_tx_mmcm_lock_in             =>      gt6_txmmcm_lock_i,
        gt6_tx_mmcm_reset_out           =>      gt6_txmmcm_reset_i,
        gt6_rx_mmcm_lock_in             =>      gt6_rxmmcm_lock_i,
        gt6_rx_mmcm_reset_out           =>      gt6_rxmmcm_reset_i,
        gt6_drp_busy_out                =>      open,
        gt6_tx_fsm_reset_done_out       =>      gt6_tx_fsm_reset_done_out,
        gt6_rx_fsm_reset_done_out       =>      gt6_rx_fsm_reset_done_out,
        gt6_data_valid_in               =>      gt6_data_valid_in,
        gt7_tx_mmcm_lock_in             =>      gt7_txmmcm_lock_i,
        gt7_tx_mmcm_reset_out           =>      gt7_txmmcm_reset_i,
        gt7_rx_mmcm_lock_in             =>      gt7_rxmmcm_lock_i,
        gt7_rx_mmcm_reset_out           =>      gt7_rxmmcm_reset_i,
        gt7_drp_busy_out                =>      open,
        gt7_tx_fsm_reset_done_out       =>      gt7_tx_fsm_reset_done_out,
        gt7_rx_fsm_reset_done_out       =>      gt7_rx_fsm_reset_done_out,
        gt7_data_valid_in               =>      gt7_data_valid_in,
        gt8_tx_mmcm_lock_in             =>      gt8_txmmcm_lock_i,
        gt8_tx_mmcm_reset_out           =>      gt8_txmmcm_reset_i,
        gt8_rx_mmcm_lock_in             =>      gt8_rxmmcm_lock_i,
        gt8_rx_mmcm_reset_out           =>      gt8_rxmmcm_reset_i,
        gt8_drp_busy_out                =>      open,
        gt8_tx_fsm_reset_done_out       =>      gt8_tx_fsm_reset_done_out,
        gt8_rx_fsm_reset_done_out       =>      gt8_rx_fsm_reset_done_out,
        gt8_data_valid_in               =>      gt8_data_valid_in,
        gt9_tx_mmcm_lock_in             =>      gt9_txmmcm_lock_i,
        gt9_tx_mmcm_reset_out           =>      gt9_txmmcm_reset_i,
        gt9_rx_mmcm_lock_in             =>      gt9_rxmmcm_lock_i,
        gt9_rx_mmcm_reset_out           =>      gt9_rxmmcm_reset_i,
        gt9_drp_busy_out                =>      open,
        gt9_tx_fsm_reset_done_out       =>      gt9_tx_fsm_reset_done_out,
        gt9_rx_fsm_reset_done_out       =>      gt9_rx_fsm_reset_done_out,
        gt9_data_valid_in               =>      gt9_data_valid_in,
        gt10_tx_mmcm_lock_in            =>      gt10_txmmcm_lock_i,
        gt10_tx_mmcm_reset_out          =>      gt10_txmmcm_reset_i,
        gt10_rx_mmcm_lock_in            =>      gt10_rxmmcm_lock_i,
        gt10_rx_mmcm_reset_out          =>      gt10_rxmmcm_reset_i,
        gt10_drp_busy_out               =>      open,
        gt10_tx_fsm_reset_done_out      =>      gt10_tx_fsm_reset_done_out,
        gt10_rx_fsm_reset_done_out      =>      gt10_rx_fsm_reset_done_out,
        gt10_data_valid_in              =>      gt10_data_valid_in,
        gt11_tx_mmcm_lock_in            =>      gt11_txmmcm_lock_i,
        gt11_tx_mmcm_reset_out          =>      gt11_txmmcm_reset_i,
        gt11_rx_mmcm_lock_in            =>      gt11_rxmmcm_lock_i,
        gt11_rx_mmcm_reset_out          =>      gt11_rxmmcm_reset_i,
        gt11_drp_busy_out               =>      open,
        gt11_tx_fsm_reset_done_out      =>      gt11_tx_fsm_reset_done_out,
        gt11_rx_fsm_reset_done_out      =>      gt11_rx_fsm_reset_done_out,
        gt11_data_valid_in              =>      gt11_data_valid_in,
        gt12_tx_mmcm_lock_in            =>      gt12_txmmcm_lock_i,
        gt12_tx_mmcm_reset_out          =>      gt12_txmmcm_reset_i,
        gt12_rx_mmcm_lock_in            =>      gt12_rxmmcm_lock_i,
        gt12_rx_mmcm_reset_out          =>      gt12_rxmmcm_reset_i,
        gt12_drp_busy_out               =>      open,
        gt12_tx_fsm_reset_done_out      =>      gt12_tx_fsm_reset_done_out,
        gt12_rx_fsm_reset_done_out      =>      gt12_rx_fsm_reset_done_out,
        gt12_data_valid_in              =>      gt12_data_valid_in,
        gt13_tx_mmcm_lock_in            =>      gt13_txmmcm_lock_i,
        gt13_tx_mmcm_reset_out          =>      gt13_txmmcm_reset_i,
        gt13_rx_mmcm_lock_in            =>      gt13_rxmmcm_lock_i,
        gt13_rx_mmcm_reset_out          =>      gt13_rxmmcm_reset_i,
        gt13_drp_busy_out               =>      open,
        gt13_tx_fsm_reset_done_out      =>      gt13_tx_fsm_reset_done_out,
        gt13_rx_fsm_reset_done_out      =>      gt13_rx_fsm_reset_done_out,
        gt13_data_valid_in              =>      gt13_data_valid_in,
        gt14_tx_mmcm_lock_in            =>      gt14_txmmcm_lock_i,
        gt14_tx_mmcm_reset_out          =>      gt14_txmmcm_reset_i,
        gt14_rx_mmcm_lock_in            =>      gt14_rxmmcm_lock_i,
        gt14_rx_mmcm_reset_out          =>      gt14_rxmmcm_reset_i,
        gt14_drp_busy_out               =>      open,
        gt14_tx_fsm_reset_done_out      =>      gt14_tx_fsm_reset_done_out,
        gt14_rx_fsm_reset_done_out      =>      gt14_rx_fsm_reset_done_out,
        gt14_data_valid_in              =>      gt14_data_valid_in,
        gt15_tx_mmcm_lock_in            =>      gt15_txmmcm_lock_i,
        gt15_tx_mmcm_reset_out          =>      gt15_txmmcm_reset_i,
        gt15_rx_mmcm_lock_in            =>      gt15_rxmmcm_lock_i,
        gt15_rx_mmcm_reset_out          =>      gt15_rxmmcm_reset_i,
        gt15_drp_busy_out               =>      open,
        gt15_tx_fsm_reset_done_out      =>      gt15_tx_fsm_reset_done_out,
        gt15_rx_fsm_reset_done_out      =>      gt15_rx_fsm_reset_done_out,
        gt15_data_valid_in              =>      gt15_data_valid_in,
        gt16_tx_mmcm_lock_in            =>      gt16_txmmcm_lock_i,
        gt16_tx_mmcm_reset_out          =>      gt16_txmmcm_reset_i,
        gt16_rx_mmcm_lock_in            =>      gt16_rxmmcm_lock_i,
        gt16_rx_mmcm_reset_out          =>      gt16_rxmmcm_reset_i,
        gt16_drp_busy_out               =>      open,
        gt16_tx_fsm_reset_done_out      =>      gt16_tx_fsm_reset_done_out,
        gt16_rx_fsm_reset_done_out      =>      gt16_rx_fsm_reset_done_out,
        gt16_data_valid_in              =>      gt16_data_valid_in,
        gt17_tx_mmcm_lock_in            =>      gt17_txmmcm_lock_i,
        gt17_tx_mmcm_reset_out          =>      gt17_txmmcm_reset_i,
        gt17_rx_mmcm_lock_in            =>      gt17_rxmmcm_lock_i,
        gt17_rx_mmcm_reset_out          =>      gt17_rxmmcm_reset_i,
        gt17_drp_busy_out               =>      open,
        gt17_tx_fsm_reset_done_out      =>      gt17_tx_fsm_reset_done_out,
        gt17_rx_fsm_reset_done_out      =>      gt17_rx_fsm_reset_done_out,
        gt17_data_valid_in              =>      gt17_data_valid_in,
        gt18_tx_mmcm_lock_in            =>      gt18_txmmcm_lock_i,
        gt18_tx_mmcm_reset_out          =>      gt18_txmmcm_reset_i,
        gt18_rx_mmcm_lock_in            =>      gt18_rxmmcm_lock_i,
        gt18_rx_mmcm_reset_out          =>      gt18_rxmmcm_reset_i,
        gt18_drp_busy_out               =>      open,
        gt18_tx_fsm_reset_done_out      =>      gt18_tx_fsm_reset_done_out,
        gt18_rx_fsm_reset_done_out      =>      gt18_rx_fsm_reset_done_out,
        gt18_data_valid_in              =>      gt18_data_valid_in,
        gt19_tx_mmcm_lock_in            =>      gt19_txmmcm_lock_i,
        gt19_tx_mmcm_reset_out          =>      gt19_txmmcm_reset_i,
        gt19_rx_mmcm_lock_in            =>      gt19_rxmmcm_lock_i,
        gt19_rx_mmcm_reset_out          =>      gt19_rxmmcm_reset_i,
        gt19_drp_busy_out               =>      open,
        gt19_tx_fsm_reset_done_out      =>      gt19_tx_fsm_reset_done_out,
        gt19_rx_fsm_reset_done_out      =>      gt19_rx_fsm_reset_done_out,
        gt19_data_valid_in              =>      gt19_data_valid_in,
        gt20_tx_mmcm_lock_in            =>      gt20_txmmcm_lock_i,
        gt20_tx_mmcm_reset_out          =>      gt20_txmmcm_reset_i,
        gt20_rx_mmcm_lock_in            =>      gt20_rxmmcm_lock_i,
        gt20_rx_mmcm_reset_out          =>      gt20_rxmmcm_reset_i,
        gt20_drp_busy_out               =>      open,
        gt20_tx_fsm_reset_done_out      =>      gt20_tx_fsm_reset_done_out,
        gt20_rx_fsm_reset_done_out      =>      gt20_rx_fsm_reset_done_out,
        gt20_data_valid_in              =>      gt20_data_valid_in,
        gt21_tx_mmcm_lock_in            =>      gt21_txmmcm_lock_i,
        gt21_tx_mmcm_reset_out          =>      gt21_txmmcm_reset_i,
        gt21_rx_mmcm_lock_in            =>      gt21_rxmmcm_lock_i,
        gt21_rx_mmcm_reset_out          =>      gt21_rxmmcm_reset_i,
        gt21_drp_busy_out               =>      open,
        gt21_tx_fsm_reset_done_out      =>      gt21_tx_fsm_reset_done_out,
        gt21_rx_fsm_reset_done_out      =>      gt21_rx_fsm_reset_done_out,
        gt21_data_valid_in              =>      gt21_data_valid_in,
        gt22_tx_mmcm_lock_in            =>      gt22_txmmcm_lock_i,
        gt22_tx_mmcm_reset_out          =>      gt22_txmmcm_reset_i,
        gt22_rx_mmcm_lock_in            =>      gt22_rxmmcm_lock_i,
        gt22_rx_mmcm_reset_out          =>      gt22_rxmmcm_reset_i,
        gt22_drp_busy_out               =>      open,
        gt22_tx_fsm_reset_done_out      =>      gt22_tx_fsm_reset_done_out,
        gt22_rx_fsm_reset_done_out      =>      gt22_rx_fsm_reset_done_out,
        gt22_data_valid_in              =>      gt22_data_valid_in,
        gt23_tx_mmcm_lock_in            =>      gt23_txmmcm_lock_i,
        gt23_tx_mmcm_reset_out          =>      gt23_txmmcm_reset_i,
        gt23_rx_mmcm_lock_in            =>      gt23_rxmmcm_lock_i,
        gt23_rx_mmcm_reset_out          =>      gt23_rxmmcm_reset_i,
        gt23_drp_busy_out               =>      open,
        gt23_tx_fsm_reset_done_out      =>      gt23_tx_fsm_reset_done_out,
        gt23_rx_fsm_reset_done_out      =>      gt23_rx_fsm_reset_done_out,
        gt23_data_valid_in              =>      gt23_data_valid_in,
        gt24_tx_mmcm_lock_in            =>      gt24_txmmcm_lock_i,
        gt24_tx_mmcm_reset_out          =>      gt24_txmmcm_reset_i,
        gt24_rx_mmcm_lock_in            =>      gt24_rxmmcm_lock_i,
        gt24_rx_mmcm_reset_out          =>      gt24_rxmmcm_reset_i,
        gt24_drp_busy_out               =>      open,
        gt24_tx_fsm_reset_done_out      =>      gt24_tx_fsm_reset_done_out,
        gt24_rx_fsm_reset_done_out      =>      gt24_rx_fsm_reset_done_out,
        gt24_data_valid_in              =>      gt24_data_valid_in,
        gt25_tx_mmcm_lock_in            =>      gt25_txmmcm_lock_i,
        gt25_tx_mmcm_reset_out          =>      gt25_txmmcm_reset_i,
        gt25_rx_mmcm_lock_in            =>      gt25_rxmmcm_lock_i,
        gt25_rx_mmcm_reset_out          =>      gt25_rxmmcm_reset_i,
        gt25_drp_busy_out               =>      open,
        gt25_tx_fsm_reset_done_out      =>      gt25_tx_fsm_reset_done_out,
        gt25_rx_fsm_reset_done_out      =>      gt25_rx_fsm_reset_done_out,
        gt25_data_valid_in              =>      gt25_data_valid_in,
        gt26_tx_mmcm_lock_in            =>      gt26_txmmcm_lock_i,
        gt26_tx_mmcm_reset_out          =>      gt26_txmmcm_reset_i,
        gt26_rx_mmcm_lock_in            =>      gt26_rxmmcm_lock_i,
        gt26_rx_mmcm_reset_out          =>      gt26_rxmmcm_reset_i,
        gt26_drp_busy_out               =>      open,
        gt26_tx_fsm_reset_done_out      =>      gt26_tx_fsm_reset_done_out,
        gt26_rx_fsm_reset_done_out      =>      gt26_rx_fsm_reset_done_out,
        gt26_data_valid_in              =>      gt26_data_valid_in,
        gt27_tx_mmcm_lock_in            =>      gt27_txmmcm_lock_i,
        gt27_tx_mmcm_reset_out          =>      gt27_txmmcm_reset_i,
        gt27_rx_mmcm_lock_in            =>      gt27_rxmmcm_lock_i,
        gt27_rx_mmcm_reset_out          =>      gt27_rxmmcm_reset_i,
        gt27_drp_busy_out               =>      open,
        gt27_tx_fsm_reset_done_out      =>      gt27_tx_fsm_reset_done_out,
        gt27_rx_fsm_reset_done_out      =>      gt27_rx_fsm_reset_done_out,
        gt27_data_valid_in              =>      gt27_data_valid_in,
        gt28_tx_mmcm_lock_in            =>      gt28_txmmcm_lock_i,
        gt28_tx_mmcm_reset_out          =>      gt28_txmmcm_reset_i,
        gt28_rx_mmcm_lock_in            =>      gt28_rxmmcm_lock_i,
        gt28_rx_mmcm_reset_out          =>      gt28_rxmmcm_reset_i,
        gt28_drp_busy_out               =>      open,
        gt28_tx_fsm_reset_done_out      =>      gt28_tx_fsm_reset_done_out,
        gt28_rx_fsm_reset_done_out      =>      gt28_rx_fsm_reset_done_out,
        gt28_data_valid_in              =>      gt28_data_valid_in,
        gt29_tx_mmcm_lock_in            =>      gt29_txmmcm_lock_i,
        gt29_tx_mmcm_reset_out          =>      gt29_txmmcm_reset_i,
        gt29_rx_mmcm_lock_in            =>      gt29_rxmmcm_lock_i,
        gt29_rx_mmcm_reset_out          =>      gt29_rxmmcm_reset_i,
        gt29_drp_busy_out               =>      open,
        gt29_tx_fsm_reset_done_out      =>      gt29_tx_fsm_reset_done_out,
        gt29_rx_fsm_reset_done_out      =>      gt29_rx_fsm_reset_done_out,
        gt29_data_valid_in              =>      gt29_data_valid_in,
        gt30_tx_mmcm_lock_in            =>      gt30_txmmcm_lock_i,
        gt30_tx_mmcm_reset_out          =>      gt30_txmmcm_reset_i,
        gt30_rx_mmcm_lock_in            =>      gt30_rxmmcm_lock_i,
        gt30_rx_mmcm_reset_out          =>      gt30_rxmmcm_reset_i,
        gt30_drp_busy_out               =>      open,
        gt30_tx_fsm_reset_done_out      =>      gt30_tx_fsm_reset_done_out,
        gt30_rx_fsm_reset_done_out      =>      gt30_rx_fsm_reset_done_out,
        gt30_data_valid_in              =>      gt30_data_valid_in,
        gt31_tx_mmcm_lock_in            =>      gt31_txmmcm_lock_i,
        gt31_tx_mmcm_reset_out          =>      gt31_txmmcm_reset_i,
        gt31_rx_mmcm_lock_in            =>      gt31_rxmmcm_lock_i,
        gt31_rx_mmcm_reset_out          =>      gt31_rxmmcm_reset_i,
        gt31_drp_busy_out               =>      open,
        gt31_tx_fsm_reset_done_out      =>      gt31_tx_fsm_reset_done_out,
        gt31_rx_fsm_reset_done_out      =>      gt31_rx_fsm_reset_done_out,
        gt31_data_valid_in              =>      gt31_data_valid_in,

        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT0  (X1Y4)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt0_drpaddr_in                  =>      gt0_drpaddr_in,
        gt0_drpclk_in                   =>      sysclk_in_i,
        gt0_drpdi_in                    =>      gt0_drpdi_in,
        gt0_drpdo_out                   =>      gt0_drpdo_out,
        gt0_drpen_in                    =>      gt0_drpen_in,
        gt0_drprdy_out                  =>      gt0_drprdy_out,
        gt0_drpwe_in                    =>      gt0_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt0_eyescanreset_in             =>      gt0_eyescanreset_in,
        gt0_rxuserrdy_in                =>      gt0_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt0_eyescandataerror_out        =>      gt0_eyescandataerror_out,
        gt0_eyescantrigger_in           =>      gt0_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt0_rxslide_in                  =>      gt0_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt0_dmonitorout_out             =>      gt0_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt0_rxusrclk_in                 =>      gt0_rxusrclk_i,
        gt0_rxusrclk2_in                =>      gt0_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt0_rxdata_out                  =>      gt0_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt0_rxdisperr_out               =>      gt0_rxdisperr_out,
        gt0_rxnotintable_out            =>      gt0_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt0_gthrxn_in                   =>      gt0_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt0_rxphmonitor_out             =>      gt0_rxphmonitor_out,
        gt0_rxphslipmonitor_out         =>      gt0_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt0_rxbyteisaligned_out         =>      gt0_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt0_rxmonitorout_out            =>      gt0_rxmonitorout_out,
        gt0_rxmonitorsel_in             =>      gt0_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt0_rxoutclk_out                =>      gt0_rxoutclk_i,
        gt0_rxoutclkfabric_out          =>      gt0_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt0_gtrxreset_in                =>      gt0_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt0_rxcharisk_out               =>      gt0_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt0_gthrxp_in                   =>      gt0_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt0_rxresetdone_out             =>      gt0_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt0_gttxreset_in                =>      gt0_gttxreset_in,
        gt0_txuserrdy_in                =>      gt0_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt0_txusrclk_in                 =>      gt0_txusrclk_i,
        gt0_txusrclk2_in                =>      gt0_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt0_txdata_in                   =>      gt0_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt0_gthtxn_out                  =>      gt0_gthtxn_out,
        gt0_gthtxp_out                  =>      gt0_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt0_txoutclk_out                =>      gt0_txoutclk_i,
        gt0_txoutclkfabric_out          =>      gt0_txoutclkfabric_out,
        gt0_txoutclkpcs_out             =>      gt0_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt0_txresetdone_out             =>      gt0_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt0_txcharisk_in                =>      gt0_txcharisk_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT1  (X1Y5)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt1_drpaddr_in                  =>      gt1_drpaddr_in,
        gt1_drpclk_in                   =>      sysclk_in_i,
        gt1_drpdi_in                    =>      gt1_drpdi_in,
        gt1_drpdo_out                   =>      gt1_drpdo_out,
        gt1_drpen_in                    =>      gt1_drpen_in,
        gt1_drprdy_out                  =>      gt1_drprdy_out,
        gt1_drpwe_in                    =>      gt1_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt1_eyescanreset_in             =>      gt1_eyescanreset_in,
        gt1_rxuserrdy_in                =>      gt1_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt1_eyescandataerror_out        =>      gt1_eyescandataerror_out,
        gt1_eyescantrigger_in           =>      gt1_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt1_rxslide_in                  =>      gt1_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt1_dmonitorout_out             =>      gt1_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt1_rxusrclk_in                 =>      gt1_rxusrclk_i,
        gt1_rxusrclk2_in                =>      gt1_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt1_rxdata_out                  =>      gt1_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt1_rxdisperr_out               =>      gt1_rxdisperr_out,
        gt1_rxnotintable_out            =>      gt1_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt1_gthrxn_in                   =>      gt1_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt1_rxphmonitor_out             =>      gt1_rxphmonitor_out,
        gt1_rxphslipmonitor_out         =>      gt1_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt1_rxbyteisaligned_out         =>      gt1_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt1_rxmonitorout_out            =>      gt1_rxmonitorout_out,
        gt1_rxmonitorsel_in             =>      gt1_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt1_rxoutclk_out                =>      gt1_rxoutclk_i,
        gt1_rxoutclkfabric_out          =>      gt1_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt1_gtrxreset_in                =>      gt1_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt1_rxcharisk_out               =>      gt1_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt1_gthrxp_in                   =>      gt1_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt1_rxresetdone_out             =>      gt1_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt1_gttxreset_in                =>      gt1_gttxreset_in,
        gt1_txuserrdy_in                =>      gt1_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt1_txusrclk_in                 =>      gt1_txusrclk_i,
        gt1_txusrclk2_in                =>      gt1_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt1_txdata_in                   =>      gt1_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt1_gthtxn_out                  =>      gt1_gthtxn_out,
        gt1_gthtxp_out                  =>      gt1_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt1_txoutclk_out                =>      gt1_txoutclk_i,
        gt1_txoutclkfabric_out          =>      gt1_txoutclkfabric_out,
        gt1_txoutclkpcs_out             =>      gt1_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt1_txresetdone_out             =>      gt1_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt1_txcharisk_in                =>      gt1_txcharisk_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT2  (X1Y6)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt2_drpaddr_in                  =>      gt2_drpaddr_in,
        gt2_drpclk_in                   =>      sysclk_in_i,
        gt2_drpdi_in                    =>      gt2_drpdi_in,
        gt2_drpdo_out                   =>      gt2_drpdo_out,
        gt2_drpen_in                    =>      gt2_drpen_in,
        gt2_drprdy_out                  =>      gt2_drprdy_out,
        gt2_drpwe_in                    =>      gt2_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt2_eyescanreset_in             =>      gt2_eyescanreset_in,
        gt2_rxuserrdy_in                =>      gt2_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt2_eyescandataerror_out        =>      gt2_eyescandataerror_out,
        gt2_eyescantrigger_in           =>      gt2_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt2_rxslide_in                  =>      gt2_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt2_dmonitorout_out             =>      gt2_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt2_rxusrclk_in                 =>      gt2_rxusrclk_i,
        gt2_rxusrclk2_in                =>      gt2_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt2_rxdata_out                  =>      gt2_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt2_rxdisperr_out               =>      gt2_rxdisperr_out,
        gt2_rxnotintable_out            =>      gt2_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt2_gthrxn_in                   =>      gt2_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt2_rxphmonitor_out             =>      gt2_rxphmonitor_out,
        gt2_rxphslipmonitor_out         =>      gt2_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt2_rxbyteisaligned_out         =>      gt2_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt2_rxmonitorout_out            =>      gt2_rxmonitorout_out,
        gt2_rxmonitorsel_in             =>      gt2_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt2_rxoutclk_out                =>      gt2_rxoutclk_i,
        gt2_rxoutclkfabric_out          =>      gt2_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt2_gtrxreset_in                =>      gt2_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt2_rxcharisk_out               =>      gt2_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt2_gthrxp_in                   =>      gt2_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt2_rxresetdone_out             =>      gt2_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt2_gttxreset_in                =>      gt2_gttxreset_in,
        gt2_txuserrdy_in                =>      gt2_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt2_txusrclk_in                 =>      gt2_txusrclk_i,
        gt2_txusrclk2_in                =>      gt2_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt2_txdata_in                   =>      gt2_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt2_gthtxn_out                  =>      gt2_gthtxn_out,
        gt2_gthtxp_out                  =>      gt2_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt2_txoutclk_out                =>      gt2_txoutclk_i,
        gt2_txoutclkfabric_out          =>      gt2_txoutclkfabric_out,
        gt2_txoutclkpcs_out             =>      gt2_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt2_txresetdone_out             =>      gt2_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt2_txcharisk_in                =>      gt2_txcharisk_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT3  (X1Y7)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt3_drpaddr_in                  =>      gt3_drpaddr_in,
        gt3_drpclk_in                   =>      sysclk_in_i,
        gt3_drpdi_in                    =>      gt3_drpdi_in,
        gt3_drpdo_out                   =>      gt3_drpdo_out,
        gt3_drpen_in                    =>      gt3_drpen_in,
        gt3_drprdy_out                  =>      gt3_drprdy_out,
        gt3_drpwe_in                    =>      gt3_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt3_eyescanreset_in             =>      gt3_eyescanreset_in,
        gt3_rxuserrdy_in                =>      gt3_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt3_eyescandataerror_out        =>      gt3_eyescandataerror_out,
        gt3_eyescantrigger_in           =>      gt3_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt3_rxslide_in                  =>      gt3_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt3_dmonitorout_out             =>      gt3_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt3_rxusrclk_in                 =>      gt3_rxusrclk_i,
        gt3_rxusrclk2_in                =>      gt3_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt3_rxdata_out                  =>      gt3_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt3_rxdisperr_out               =>      gt3_rxdisperr_out,
        gt3_rxnotintable_out            =>      gt3_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt3_gthrxn_in                   =>      gt3_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt3_rxphmonitor_out             =>      gt3_rxphmonitor_out,
        gt3_rxphslipmonitor_out         =>      gt3_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt3_rxbyteisaligned_out         =>      gt3_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt3_rxmonitorout_out            =>      gt3_rxmonitorout_out,
        gt3_rxmonitorsel_in             =>      gt3_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt3_rxoutclk_out                =>      gt3_rxoutclk_i,
        gt3_rxoutclkfabric_out          =>      gt3_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt3_gtrxreset_in                =>      gt3_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt3_rxcharisk_out               =>      gt3_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt3_gthrxp_in                   =>      gt3_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt3_rxresetdone_out             =>      gt3_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt3_gttxreset_in                =>      gt3_gttxreset_in,
        gt3_txuserrdy_in                =>      gt3_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt3_txusrclk_in                 =>      gt3_txusrclk_i,
        gt3_txusrclk2_in                =>      gt3_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt3_txdata_in                   =>      gt3_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt3_gthtxn_out                  =>      gt3_gthtxn_out,
        gt3_gthtxp_out                  =>      gt3_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt3_txoutclk_out                =>      gt3_txoutclk_i,
        gt3_txoutclkfabric_out          =>      gt3_txoutclkfabric_out,
        gt3_txoutclkpcs_out             =>      gt3_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt3_txresetdone_out             =>      gt3_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt3_txcharisk_in                =>      gt3_txcharisk_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT4  (X1Y8)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt4_drpaddr_in                  =>      gt4_drpaddr_in,
        gt4_drpclk_in                   =>      sysclk_in_i,
        gt4_drpdi_in                    =>      gt4_drpdi_in,
        gt4_drpdo_out                   =>      gt4_drpdo_out,
        gt4_drpen_in                    =>      gt4_drpen_in,
        gt4_drprdy_out                  =>      gt4_drprdy_out,
        gt4_drpwe_in                    =>      gt4_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt4_eyescanreset_in             =>      gt4_eyescanreset_in,
        gt4_rxuserrdy_in                =>      gt4_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt4_eyescandataerror_out        =>      gt4_eyescandataerror_out,
        gt4_eyescantrigger_in           =>      gt4_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt4_rxslide_in                  =>      gt4_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt4_dmonitorout_out             =>      gt4_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt4_rxusrclk_in                 =>      gt4_rxusrclk_i,
        gt4_rxusrclk2_in                =>      gt4_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt4_rxdata_out                  =>      gt4_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt4_rxdisperr_out               =>      gt4_rxdisperr_out,
        gt4_rxnotintable_out            =>      gt4_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt4_gthrxn_in                   =>      gt4_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt4_rxphmonitor_out             =>      gt4_rxphmonitor_out,
        gt4_rxphslipmonitor_out         =>      gt4_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt4_rxbyteisaligned_out         =>      gt4_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt4_rxmonitorout_out            =>      gt4_rxmonitorout_out,
        gt4_rxmonitorsel_in             =>      gt4_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt4_rxoutclk_out                =>      gt4_rxoutclk_i,
        gt4_rxoutclkfabric_out          =>      gt4_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt4_gtrxreset_in                =>      gt4_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt4_rxcharisk_out               =>      gt4_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt4_gthrxp_in                   =>      gt4_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt4_rxresetdone_out             =>      gt4_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt4_gttxreset_in                =>      gt4_gttxreset_in,
        gt4_txuserrdy_in                =>      gt4_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt4_txusrclk_in                 =>      gt4_txusrclk_i,
        gt4_txusrclk2_in                =>      gt4_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt4_txdata_in                   =>      gt4_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt4_gthtxn_out                  =>      gt4_gthtxn_out,
        gt4_gthtxp_out                  =>      gt4_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt4_txoutclk_out                =>      gt4_txoutclk_i,
        gt4_txoutclkfabric_out          =>      gt4_txoutclkfabric_out,
        gt4_txoutclkpcs_out             =>      gt4_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt4_txresetdone_out             =>      gt4_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt4_txcharisk_in                =>      gt4_txcharisk_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT5  (X1Y9)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt5_drpaddr_in                  =>      gt5_drpaddr_in,
        gt5_drpclk_in                   =>      sysclk_in_i,
        gt5_drpdi_in                    =>      gt5_drpdi_in,
        gt5_drpdo_out                   =>      gt5_drpdo_out,
        gt5_drpen_in                    =>      gt5_drpen_in,
        gt5_drprdy_out                  =>      gt5_drprdy_out,
        gt5_drpwe_in                    =>      gt5_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt5_eyescanreset_in             =>      gt5_eyescanreset_in,
        gt5_rxuserrdy_in                =>      gt5_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt5_eyescandataerror_out        =>      gt5_eyescandataerror_out,
        gt5_eyescantrigger_in           =>      gt5_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt5_rxslide_in                  =>      gt5_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt5_dmonitorout_out             =>      gt5_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt5_rxusrclk_in                 =>      gt5_rxusrclk_i,
        gt5_rxusrclk2_in                =>      gt5_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt5_rxdata_out                  =>      gt5_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt5_rxdisperr_out               =>      gt5_rxdisperr_out,
        gt5_rxnotintable_out            =>      gt5_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt5_gthrxn_in                   =>      gt5_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt5_rxphmonitor_out             =>      gt5_rxphmonitor_out,
        gt5_rxphslipmonitor_out         =>      gt5_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt5_rxbyteisaligned_out         =>      gt5_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt5_rxmonitorout_out            =>      gt5_rxmonitorout_out,
        gt5_rxmonitorsel_in             =>      gt5_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt5_rxoutclk_out                =>      gt5_rxoutclk_i,
        gt5_rxoutclkfabric_out          =>      gt5_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt5_gtrxreset_in                =>      gt5_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt5_rxcharisk_out               =>      gt5_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt5_gthrxp_in                   =>      gt5_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt5_rxresetdone_out             =>      gt5_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt5_gttxreset_in                =>      gt5_gttxreset_in,
        gt5_txuserrdy_in                =>      gt5_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt5_txusrclk_in                 =>      gt5_txusrclk_i,
        gt5_txusrclk2_in                =>      gt5_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt5_txdata_in                   =>      gt5_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt5_gthtxn_out                  =>      gt5_gthtxn_out,
        gt5_gthtxp_out                  =>      gt5_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt5_txoutclk_out                =>      gt5_txoutclk_i,
        gt5_txoutclkfabric_out          =>      gt5_txoutclkfabric_out,
        gt5_txoutclkpcs_out             =>      gt5_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt5_txresetdone_out             =>      gt5_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt5_txcharisk_in                =>      gt5_txcharisk_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT6  (X1Y10)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt6_drpaddr_in                  =>      gt6_drpaddr_in,
        gt6_drpclk_in                   =>      sysclk_in_i,
        gt6_drpdi_in                    =>      gt6_drpdi_in,
        gt6_drpdo_out                   =>      gt6_drpdo_out,
        gt6_drpen_in                    =>      gt6_drpen_in,
        gt6_drprdy_out                  =>      gt6_drprdy_out,
        gt6_drpwe_in                    =>      gt6_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt6_eyescanreset_in             =>      gt6_eyescanreset_in,
        gt6_rxuserrdy_in                =>      gt6_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt6_eyescandataerror_out        =>      gt6_eyescandataerror_out,
        gt6_eyescantrigger_in           =>      gt6_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt6_rxslide_in                  =>      gt6_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt6_dmonitorout_out             =>      gt6_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt6_rxusrclk_in                 =>      gt6_rxusrclk_i,
        gt6_rxusrclk2_in                =>      gt6_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt6_rxdata_out                  =>      gt6_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt6_rxdisperr_out               =>      gt6_rxdisperr_out,
        gt6_rxnotintable_out            =>      gt6_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt6_gthrxn_in                   =>      gt6_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt6_rxphmonitor_out             =>      gt6_rxphmonitor_out,
        gt6_rxphslipmonitor_out         =>      gt6_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt6_rxbyteisaligned_out         =>      gt6_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt6_rxmonitorout_out            =>      gt6_rxmonitorout_out,
        gt6_rxmonitorsel_in             =>      gt6_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt6_rxoutclk_out                =>      gt6_rxoutclk_i,
        gt6_rxoutclkfabric_out          =>      gt6_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt6_gtrxreset_in                =>      gt6_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt6_rxcharisk_out               =>      gt6_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt6_gthrxp_in                   =>      gt6_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt6_rxresetdone_out             =>      gt6_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt6_gttxreset_in                =>      gt6_gttxreset_in,
        gt6_txuserrdy_in                =>      gt6_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt6_txusrclk_in                 =>      gt6_txusrclk_i,
        gt6_txusrclk2_in                =>      gt6_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt6_txdata_in                   =>      gt6_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt6_gthtxn_out                  =>      gt6_gthtxn_out,
        gt6_gthtxp_out                  =>      gt6_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt6_txoutclk_out                =>      gt6_txoutclk_i,
        gt6_txoutclkfabric_out          =>      gt6_txoutclkfabric_out,
        gt6_txoutclkpcs_out             =>      gt6_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt6_txresetdone_out             =>      gt6_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt6_txcharisk_in                =>      gt6_txcharisk_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT7  (X1Y11)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt7_drpaddr_in                  =>      gt7_drpaddr_in,
        gt7_drpclk_in                   =>      sysclk_in_i,
        gt7_drpdi_in                    =>      gt7_drpdi_in,
        gt7_drpdo_out                   =>      gt7_drpdo_out,
        gt7_drpen_in                    =>      gt7_drpen_in,
        gt7_drprdy_out                  =>      gt7_drprdy_out,
        gt7_drpwe_in                    =>      gt7_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt7_eyescanreset_in             =>      gt7_eyescanreset_in,
        gt7_rxuserrdy_in                =>      gt7_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt7_eyescandataerror_out        =>      gt7_eyescandataerror_out,
        gt7_eyescantrigger_in           =>      gt7_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt7_rxslide_in                  =>      gt7_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt7_dmonitorout_out             =>      gt7_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt7_rxusrclk_in                 =>      gt7_rxusrclk_i,
        gt7_rxusrclk2_in                =>      gt7_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt7_rxdata_out                  =>      gt7_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt7_rxdisperr_out               =>      gt7_rxdisperr_out,
        gt7_rxnotintable_out            =>      gt7_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt7_gthrxn_in                   =>      gt7_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt7_rxphmonitor_out             =>      gt7_rxphmonitor_out,
        gt7_rxphslipmonitor_out         =>      gt7_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt7_rxbyteisaligned_out         =>      gt7_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt7_rxmonitorout_out            =>      gt7_rxmonitorout_out,
        gt7_rxmonitorsel_in             =>      gt7_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt7_rxoutclk_out                =>      gt7_rxoutclk_i,
        gt7_rxoutclkfabric_out          =>      gt7_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt7_gtrxreset_in                =>      gt7_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt7_rxcharisk_out               =>      gt7_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt7_gthrxp_in                   =>      gt7_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt7_rxresetdone_out             =>      gt7_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt7_gttxreset_in                =>      gt7_gttxreset_in,
        gt7_txuserrdy_in                =>      gt7_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt7_txusrclk_in                 =>      gt7_txusrclk_i,
        gt7_txusrclk2_in                =>      gt7_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt7_txdata_in                   =>      gt7_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt7_gthtxn_out                  =>      gt7_gthtxn_out,
        gt7_gthtxp_out                  =>      gt7_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt7_txoutclk_out                =>      gt7_txoutclk_i,
        gt7_txoutclkfabric_out          =>      gt7_txoutclkfabric_out,
        gt7_txoutclkpcs_out             =>      gt7_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt7_txresetdone_out             =>      gt7_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt7_txcharisk_in                =>      gt7_txcharisk_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT8  (X1Y12)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt8_drpaddr_in                  =>      gt8_drpaddr_in,
        gt8_drpclk_in                   =>      sysclk_in_i,
        gt8_drpdi_in                    =>      gt8_drpdi_in,
        gt8_drpdo_out                   =>      gt8_drpdo_out,
        gt8_drpen_in                    =>      gt8_drpen_in,
        gt8_drprdy_out                  =>      gt8_drprdy_out,
        gt8_drpwe_in                    =>      gt8_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt8_eyescanreset_in             =>      gt8_eyescanreset_in,
        gt8_rxuserrdy_in                =>      gt8_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt8_eyescandataerror_out        =>      gt8_eyescandataerror_out,
        gt8_eyescantrigger_in           =>      gt8_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt8_rxslide_in                  =>      gt8_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt8_dmonitorout_out             =>      gt8_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt8_rxusrclk_in                 =>      gt8_rxusrclk_i,
        gt8_rxusrclk2_in                =>      gt8_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt8_rxdata_out                  =>      gt8_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt8_rxdisperr_out               =>      gt8_rxdisperr_out,
        gt8_rxnotintable_out            =>      gt8_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt8_gthrxn_in                   =>      gt8_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt8_rxphmonitor_out             =>      gt8_rxphmonitor_out,
        gt8_rxphslipmonitor_out         =>      gt8_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt8_rxbyteisaligned_out         =>      gt8_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt8_rxmonitorout_out            =>      gt8_rxmonitorout_out,
        gt8_rxmonitorsel_in             =>      gt8_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt8_rxoutclk_out                =>      gt8_rxoutclk_i,
        gt8_rxoutclkfabric_out          =>      gt8_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt8_gtrxreset_in                =>      gt8_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt8_rxcharisk_out               =>      gt8_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt8_gthrxp_in                   =>      gt8_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt8_rxresetdone_out             =>      gt8_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt8_gttxreset_in                =>      gt8_gttxreset_in,
        gt8_txuserrdy_in                =>      gt8_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt8_txusrclk_in                 =>      gt8_txusrclk_i,
        gt8_txusrclk2_in                =>      gt8_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt8_txdata_in                   =>      gt8_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt8_gthtxn_out                  =>      gt8_gthtxn_out,
        gt8_gthtxp_out                  =>      gt8_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt8_txoutclk_out                =>      gt8_txoutclk_i,
        gt8_txoutclkfabric_out          =>      gt8_txoutclkfabric_out,
        gt8_txoutclkpcs_out             =>      gt8_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt8_txresetdone_out             =>      gt8_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt8_txcharisk_in                =>      gt8_txcharisk_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT9  (X1Y13)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt9_drpaddr_in                  =>      gt9_drpaddr_in,
        gt9_drpclk_in                   =>      sysclk_in_i,
        gt9_drpdi_in                    =>      gt9_drpdi_in,
        gt9_drpdo_out                   =>      gt9_drpdo_out,
        gt9_drpen_in                    =>      gt9_drpen_in,
        gt9_drprdy_out                  =>      gt9_drprdy_out,
        gt9_drpwe_in                    =>      gt9_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt9_eyescanreset_in             =>      gt9_eyescanreset_in,
        gt9_rxuserrdy_in                =>      gt9_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt9_eyescandataerror_out        =>      gt9_eyescandataerror_out,
        gt9_eyescantrigger_in           =>      gt9_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt9_rxslide_in                  =>      gt9_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt9_dmonitorout_out             =>      gt9_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt9_rxusrclk_in                 =>      gt9_rxusrclk_i,
        gt9_rxusrclk2_in                =>      gt9_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt9_rxdata_out                  =>      gt9_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt9_rxdisperr_out               =>      gt9_rxdisperr_out,
        gt9_rxnotintable_out            =>      gt9_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt9_gthrxn_in                   =>      gt9_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt9_rxphmonitor_out             =>      gt9_rxphmonitor_out,
        gt9_rxphslipmonitor_out         =>      gt9_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt9_rxbyteisaligned_out         =>      gt9_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt9_rxmonitorout_out            =>      gt9_rxmonitorout_out,
        gt9_rxmonitorsel_in             =>      gt9_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt9_rxoutclk_out                =>      gt9_rxoutclk_i,
        gt9_rxoutclkfabric_out          =>      gt9_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt9_gtrxreset_in                =>      gt9_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt9_rxcharisk_out               =>      gt9_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt9_gthrxp_in                   =>      gt9_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt9_rxresetdone_out             =>      gt9_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt9_gttxreset_in                =>      gt9_gttxreset_in,
        gt9_txuserrdy_in                =>      gt9_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt9_txusrclk_in                 =>      gt9_txusrclk_i,
        gt9_txusrclk2_in                =>      gt9_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt9_txdata_in                   =>      gt9_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt9_gthtxn_out                  =>      gt9_gthtxn_out,
        gt9_gthtxp_out                  =>      gt9_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt9_txoutclk_out                =>      gt9_txoutclk_i,
        gt9_txoutclkfabric_out          =>      gt9_txoutclkfabric_out,
        gt9_txoutclkpcs_out             =>      gt9_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt9_txresetdone_out             =>      gt9_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt9_txcharisk_in                =>      gt9_txcharisk_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT10  (X1Y14)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt10_drpaddr_in                 =>      gt10_drpaddr_in,
        gt10_drpclk_in                  =>      sysclk_in_i,
        gt10_drpdi_in                   =>      gt10_drpdi_in,
        gt10_drpdo_out                  =>      gt10_drpdo_out,
        gt10_drpen_in                   =>      gt10_drpen_in,
        gt10_drprdy_out                 =>      gt10_drprdy_out,
        gt10_drpwe_in                   =>      gt10_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt10_eyescanreset_in            =>      gt10_eyescanreset_in,
        gt10_rxuserrdy_in               =>      gt10_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt10_eyescandataerror_out       =>      gt10_eyescandataerror_out,
        gt10_eyescantrigger_in          =>      gt10_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt10_rxslide_in                 =>      gt10_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt10_dmonitorout_out            =>      gt10_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt10_rxusrclk_in                =>      gt10_rxusrclk_i,
        gt10_rxusrclk2_in               =>      gt10_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt10_rxdata_out                 =>      gt10_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt10_rxdisperr_out              =>      gt10_rxdisperr_out,
        gt10_rxnotintable_out           =>      gt10_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt10_gthrxn_in                  =>      gt10_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt10_rxphmonitor_out            =>      gt10_rxphmonitor_out,
        gt10_rxphslipmonitor_out        =>      gt10_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt10_rxbyteisaligned_out        =>      gt10_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt10_rxmonitorout_out           =>      gt10_rxmonitorout_out,
        gt10_rxmonitorsel_in            =>      gt10_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt10_rxoutclk_out               =>      gt10_rxoutclk_i,
        gt10_rxoutclkfabric_out         =>      gt10_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt10_gtrxreset_in               =>      gt10_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt10_rxcharisk_out              =>      gt10_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt10_gthrxp_in                  =>      gt10_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt10_rxresetdone_out            =>      gt10_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt10_gttxreset_in               =>      gt10_gttxreset_in,
        gt10_txuserrdy_in               =>      gt10_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt10_txusrclk_in                =>      gt10_txusrclk_i,
        gt10_txusrclk2_in               =>      gt10_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt10_txdata_in                  =>      gt10_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt10_gthtxn_out                 =>      gt10_gthtxn_out,
        gt10_gthtxp_out                 =>      gt10_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt10_txoutclk_out               =>      gt10_txoutclk_i,
        gt10_txoutclkfabric_out         =>      gt10_txoutclkfabric_out,
        gt10_txoutclkpcs_out            =>      gt10_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt10_txresetdone_out            =>      gt10_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt10_txcharisk_in               =>      gt10_txcharisk_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT11  (X1Y15)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt11_drpaddr_in                 =>      gt11_drpaddr_in,
        gt11_drpclk_in                  =>      sysclk_in_i,
        gt11_drpdi_in                   =>      gt11_drpdi_in,
        gt11_drpdo_out                  =>      gt11_drpdo_out,
        gt11_drpen_in                   =>      gt11_drpen_in,
        gt11_drprdy_out                 =>      gt11_drprdy_out,
        gt11_drpwe_in                   =>      gt11_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt11_eyescanreset_in            =>      gt11_eyescanreset_in,
        gt11_rxuserrdy_in               =>      gt11_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt11_eyescandataerror_out       =>      gt11_eyescandataerror_out,
        gt11_eyescantrigger_in          =>      gt11_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt11_rxslide_in                 =>      gt11_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt11_dmonitorout_out            =>      gt11_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt11_rxusrclk_in                =>      gt11_rxusrclk_i,
        gt11_rxusrclk2_in               =>      gt11_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt11_rxdata_out                 =>      gt11_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt11_rxdisperr_out              =>      gt11_rxdisperr_out,
        gt11_rxnotintable_out           =>      gt11_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt11_gthrxn_in                  =>      gt11_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt11_rxphmonitor_out            =>      gt11_rxphmonitor_out,
        gt11_rxphslipmonitor_out        =>      gt11_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt11_rxbyteisaligned_out        =>      gt11_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt11_rxmonitorout_out           =>      gt11_rxmonitorout_out,
        gt11_rxmonitorsel_in            =>      gt11_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt11_rxoutclk_out               =>      gt11_rxoutclk_i,
        gt11_rxoutclkfabric_out         =>      gt11_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt11_gtrxreset_in               =>      gt11_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt11_rxcharisk_out              =>      gt11_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt11_gthrxp_in                  =>      gt11_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt11_rxresetdone_out            =>      gt11_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt11_gttxreset_in               =>      gt11_gttxreset_in,
        gt11_txuserrdy_in               =>      gt11_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt11_txusrclk_in                =>      gt11_txusrclk_i,
        gt11_txusrclk2_in               =>      gt11_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt11_txdata_in                  =>      gt11_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt11_gthtxn_out                 =>      gt11_gthtxn_out,
        gt11_gthtxp_out                 =>      gt11_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt11_txoutclk_out               =>      gt11_txoutclk_i,
        gt11_txoutclkfabric_out         =>      gt11_txoutclkfabric_out,
        gt11_txoutclkpcs_out            =>      gt11_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt11_txresetdone_out            =>      gt11_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt11_txcharisk_in               =>      gt11_txcharisk_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT12  (X1Y16)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt12_drpaddr_in                 =>      gt12_drpaddr_in,
        gt12_drpclk_in                  =>      sysclk_in_i,
        gt12_drpdi_in                   =>      gt12_drpdi_in,
        gt12_drpdo_out                  =>      gt12_drpdo_out,
        gt12_drpen_in                   =>      gt12_drpen_in,
        gt12_drprdy_out                 =>      gt12_drprdy_out,
        gt12_drpwe_in                   =>      gt12_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt12_eyescanreset_in            =>      gt12_eyescanreset_in,
        gt12_rxuserrdy_in               =>      gt12_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt12_eyescandataerror_out       =>      gt12_eyescandataerror_out,
        gt12_eyescantrigger_in          =>      gt12_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt12_rxslide_in                 =>      gt12_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt12_dmonitorout_out            =>      gt12_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt12_rxusrclk_in                =>      gt12_rxusrclk_i,
        gt12_rxusrclk2_in               =>      gt12_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt12_rxdata_out                 =>      gt12_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt12_rxdisperr_out              =>      gt12_rxdisperr_out,
        gt12_rxnotintable_out           =>      gt12_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt12_gthrxn_in                  =>      gt12_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt12_rxphmonitor_out            =>      gt12_rxphmonitor_out,
        gt12_rxphslipmonitor_out        =>      gt12_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt12_rxbyteisaligned_out        =>      gt12_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt12_rxmonitorout_out           =>      gt12_rxmonitorout_out,
        gt12_rxmonitorsel_in            =>      gt12_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt12_rxoutclk_out               =>      gt12_rxoutclk_i,
        gt12_rxoutclkfabric_out         =>      gt12_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt12_gtrxreset_in               =>      gt12_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt12_rxcharisk_out              =>      gt12_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt12_gthrxp_in                  =>      gt12_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt12_rxresetdone_out            =>      gt12_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt12_gttxreset_in               =>      gt12_gttxreset_in,
        gt12_txuserrdy_in               =>      gt12_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt12_txusrclk_in                =>      gt12_txusrclk_i,
        gt12_txusrclk2_in               =>      gt12_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt12_txdata_in                  =>      gt12_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt12_gthtxn_out                 =>      gt12_gthtxn_out,
        gt12_gthtxp_out                 =>      gt12_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt12_txoutclk_out               =>      gt12_txoutclk_i,
        gt12_txoutclkfabric_out         =>      gt12_txoutclkfabric_out,
        gt12_txoutclkpcs_out            =>      gt12_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt12_txresetdone_out            =>      gt12_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt12_txcharisk_in               =>      gt12_txcharisk_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT13  (X1Y17)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt13_drpaddr_in                 =>      gt13_drpaddr_in,
        gt13_drpclk_in                  =>      sysclk_in_i,
        gt13_drpdi_in                   =>      gt13_drpdi_in,
        gt13_drpdo_out                  =>      gt13_drpdo_out,
        gt13_drpen_in                   =>      gt13_drpen_in,
        gt13_drprdy_out                 =>      gt13_drprdy_out,
        gt13_drpwe_in                   =>      gt13_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt13_eyescanreset_in            =>      gt13_eyescanreset_in,
        gt13_rxuserrdy_in               =>      gt13_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt13_eyescandataerror_out       =>      gt13_eyescandataerror_out,
        gt13_eyescantrigger_in          =>      gt13_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt13_rxslide_in                 =>      gt13_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt13_dmonitorout_out            =>      gt13_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt13_rxusrclk_in                =>      gt13_rxusrclk_i,
        gt13_rxusrclk2_in               =>      gt13_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt13_rxdata_out                 =>      gt13_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt13_rxdisperr_out              =>      gt13_rxdisperr_out,
        gt13_rxnotintable_out           =>      gt13_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt13_gthrxn_in                  =>      gt13_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt13_rxphmonitor_out            =>      gt13_rxphmonitor_out,
        gt13_rxphslipmonitor_out        =>      gt13_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt13_rxbyteisaligned_out        =>      gt13_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt13_rxmonitorout_out           =>      gt13_rxmonitorout_out,
        gt13_rxmonitorsel_in            =>      gt13_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt13_rxoutclk_out               =>      gt13_rxoutclk_i,
        gt13_rxoutclkfabric_out         =>      gt13_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt13_gtrxreset_in               =>      gt13_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt13_rxcharisk_out              =>      gt13_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt13_gthrxp_in                  =>      gt13_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt13_rxresetdone_out            =>      gt13_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt13_gttxreset_in               =>      gt13_gttxreset_in,
        gt13_txuserrdy_in               =>      gt13_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt13_txusrclk_in                =>      gt13_txusrclk_i,
        gt13_txusrclk2_in               =>      gt13_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt13_txdata_in                  =>      gt13_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt13_gthtxn_out                 =>      gt13_gthtxn_out,
        gt13_gthtxp_out                 =>      gt13_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt13_txoutclk_out               =>      gt13_txoutclk_i,
        gt13_txoutclkfabric_out         =>      gt13_txoutclkfabric_out,
        gt13_txoutclkpcs_out            =>      gt13_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt13_txresetdone_out            =>      gt13_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt13_txcharisk_in               =>      gt13_txcharisk_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT14  (X1Y18)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt14_drpaddr_in                 =>      gt14_drpaddr_in,
        gt14_drpclk_in                  =>      sysclk_in_i,
        gt14_drpdi_in                   =>      gt14_drpdi_in,
        gt14_drpdo_out                  =>      gt14_drpdo_out,
        gt14_drpen_in                   =>      gt14_drpen_in,
        gt14_drprdy_out                 =>      gt14_drprdy_out,
        gt14_drpwe_in                   =>      gt14_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt14_eyescanreset_in            =>      gt14_eyescanreset_in,
        gt14_rxuserrdy_in               =>      gt14_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt14_eyescandataerror_out       =>      gt14_eyescandataerror_out,
        gt14_eyescantrigger_in          =>      gt14_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt14_rxslide_in                 =>      gt14_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt14_dmonitorout_out            =>      gt14_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt14_rxusrclk_in                =>      gt14_rxusrclk_i,
        gt14_rxusrclk2_in               =>      gt14_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt14_rxdata_out                 =>      gt14_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt14_rxdisperr_out              =>      gt14_rxdisperr_out,
        gt14_rxnotintable_out           =>      gt14_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt14_gthrxn_in                  =>      gt14_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt14_rxphmonitor_out            =>      gt14_rxphmonitor_out,
        gt14_rxphslipmonitor_out        =>      gt14_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt14_rxbyteisaligned_out        =>      gt14_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt14_rxmonitorout_out           =>      gt14_rxmonitorout_out,
        gt14_rxmonitorsel_in            =>      gt14_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt14_rxoutclk_out               =>      gt14_rxoutclk_i,
        gt14_rxoutclkfabric_out         =>      gt14_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt14_gtrxreset_in               =>      gt14_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt14_rxcharisk_out              =>      gt14_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt14_gthrxp_in                  =>      gt14_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt14_rxresetdone_out            =>      gt14_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt14_gttxreset_in               =>      gt14_gttxreset_in,
        gt14_txuserrdy_in               =>      gt14_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt14_txusrclk_in                =>      gt14_txusrclk_i,
        gt14_txusrclk2_in               =>      gt14_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt14_txdata_in                  =>      gt14_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt14_gthtxn_out                 =>      gt14_gthtxn_out,
        gt14_gthtxp_out                 =>      gt14_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt14_txoutclk_out               =>      gt14_txoutclk_i,
        gt14_txoutclkfabric_out         =>      gt14_txoutclkfabric_out,
        gt14_txoutclkpcs_out            =>      gt14_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt14_txresetdone_out            =>      gt14_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt14_txcharisk_in               =>      gt14_txcharisk_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT15  (X1Y19)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt15_drpaddr_in                 =>      gt15_drpaddr_in,
        gt15_drpclk_in                  =>      sysclk_in_i,
        gt15_drpdi_in                   =>      gt15_drpdi_in,
        gt15_drpdo_out                  =>      gt15_drpdo_out,
        gt15_drpen_in                   =>      gt15_drpen_in,
        gt15_drprdy_out                 =>      gt15_drprdy_out,
        gt15_drpwe_in                   =>      gt15_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt15_eyescanreset_in            =>      gt15_eyescanreset_in,
        gt15_rxuserrdy_in               =>      gt15_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt15_eyescandataerror_out       =>      gt15_eyescandataerror_out,
        gt15_eyescantrigger_in          =>      gt15_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt15_rxslide_in                 =>      gt15_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt15_dmonitorout_out            =>      gt15_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt15_rxusrclk_in                =>      gt15_rxusrclk_i,
        gt15_rxusrclk2_in               =>      gt15_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt15_rxdata_out                 =>      gt15_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt15_rxdisperr_out              =>      gt15_rxdisperr_out,
        gt15_rxnotintable_out           =>      gt15_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt15_gthrxn_in                  =>      gt15_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt15_rxphmonitor_out            =>      gt15_rxphmonitor_out,
        gt15_rxphslipmonitor_out        =>      gt15_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt15_rxbyteisaligned_out        =>      gt15_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt15_rxmonitorout_out           =>      gt15_rxmonitorout_out,
        gt15_rxmonitorsel_in            =>      gt15_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt15_rxoutclk_out               =>      gt15_rxoutclk_i,
        gt15_rxoutclkfabric_out         =>      gt15_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt15_gtrxreset_in               =>      gt15_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt15_rxcharisk_out              =>      gt15_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt15_gthrxp_in                  =>      gt15_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt15_rxresetdone_out            =>      gt15_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt15_gttxreset_in               =>      gt15_gttxreset_in,
        gt15_txuserrdy_in               =>      gt15_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt15_txusrclk_in                =>      gt15_txusrclk_i,
        gt15_txusrclk2_in               =>      gt15_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt15_txdata_in                  =>      gt15_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt15_gthtxn_out                 =>      gt15_gthtxn_out,
        gt15_gthtxp_out                 =>      gt15_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt15_txoutclk_out               =>      gt15_txoutclk_i,
        gt15_txoutclkfabric_out         =>      gt15_txoutclkfabric_out,
        gt15_txoutclkpcs_out            =>      gt15_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt15_txresetdone_out            =>      gt15_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt15_txcharisk_in               =>      gt15_txcharisk_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT16  (X1Y20)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt16_drpaddr_in                 =>      gt16_drpaddr_in,
        gt16_drpclk_in                  =>      sysclk_in_i,
        gt16_drpdi_in                   =>      gt16_drpdi_in,
        gt16_drpdo_out                  =>      gt16_drpdo_out,
        gt16_drpen_in                   =>      gt16_drpen_in,
        gt16_drprdy_out                 =>      gt16_drprdy_out,
        gt16_drpwe_in                   =>      gt16_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt16_eyescanreset_in            =>      gt16_eyescanreset_in,
        gt16_rxuserrdy_in               =>      gt16_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt16_eyescandataerror_out       =>      gt16_eyescandataerror_out,
        gt16_eyescantrigger_in          =>      gt16_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt16_rxslide_in                 =>      gt16_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt16_dmonitorout_out            =>      gt16_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt16_rxusrclk_in                =>      gt16_rxusrclk_i,
        gt16_rxusrclk2_in               =>      gt16_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt16_rxdata_out                 =>      gt16_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt16_rxdisperr_out              =>      gt16_rxdisperr_out,
        gt16_rxnotintable_out           =>      gt16_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt16_gthrxn_in                  =>      gt16_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt16_rxphmonitor_out            =>      gt16_rxphmonitor_out,
        gt16_rxphslipmonitor_out        =>      gt16_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt16_rxbyteisaligned_out        =>      gt16_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt16_rxmonitorout_out           =>      gt16_rxmonitorout_out,
        gt16_rxmonitorsel_in            =>      gt16_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt16_rxoutclk_out               =>      gt16_rxoutclk_i,
        gt16_rxoutclkfabric_out         =>      gt16_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt16_gtrxreset_in               =>      gt16_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt16_rxcharisk_out              =>      gt16_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt16_gthrxp_in                  =>      gt16_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt16_rxresetdone_out            =>      gt16_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt16_gttxreset_in               =>      gt16_gttxreset_in,
        gt16_txuserrdy_in               =>      gt16_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt16_txusrclk_in                =>      gt16_txusrclk_i,
        gt16_txusrclk2_in               =>      gt16_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt16_txdata_in                  =>      gt16_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt16_gthtxn_out                 =>      gt16_gthtxn_out,
        gt16_gthtxp_out                 =>      gt16_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt16_txoutclk_out               =>      gt16_txoutclk_i,
        gt16_txoutclkfabric_out         =>      gt16_txoutclkfabric_out,
        gt16_txoutclkpcs_out            =>      gt16_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt16_txresetdone_out            =>      gt16_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt16_txcharisk_in               =>      gt16_txcharisk_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT17  (X1Y21)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt17_drpaddr_in                 =>      gt17_drpaddr_in,
        gt17_drpclk_in                  =>      sysclk_in_i,
        gt17_drpdi_in                   =>      gt17_drpdi_in,
        gt17_drpdo_out                  =>      gt17_drpdo_out,
        gt17_drpen_in                   =>      gt17_drpen_in,
        gt17_drprdy_out                 =>      gt17_drprdy_out,
        gt17_drpwe_in                   =>      gt17_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt17_eyescanreset_in            =>      gt17_eyescanreset_in,
        gt17_rxuserrdy_in               =>      gt17_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt17_eyescandataerror_out       =>      gt17_eyescandataerror_out,
        gt17_eyescantrigger_in          =>      gt17_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt17_rxslide_in                 =>      gt17_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt17_dmonitorout_out            =>      gt17_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt17_rxusrclk_in                =>      gt17_rxusrclk_i,
        gt17_rxusrclk2_in               =>      gt17_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt17_rxdata_out                 =>      gt17_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt17_rxdisperr_out              =>      gt17_rxdisperr_out,
        gt17_rxnotintable_out           =>      gt17_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt17_gthrxn_in                  =>      gt17_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt17_rxphmonitor_out            =>      gt17_rxphmonitor_out,
        gt17_rxphslipmonitor_out        =>      gt17_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt17_rxbyteisaligned_out        =>      gt17_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt17_rxmonitorout_out           =>      gt17_rxmonitorout_out,
        gt17_rxmonitorsel_in            =>      gt17_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt17_rxoutclk_out               =>      gt17_rxoutclk_i,
        gt17_rxoutclkfabric_out         =>      gt17_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt17_gtrxreset_in               =>      gt17_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt17_rxcharisk_out              =>      gt17_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt17_gthrxp_in                  =>      gt17_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt17_rxresetdone_out            =>      gt17_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt17_gttxreset_in               =>      gt17_gttxreset_in,
        gt17_txuserrdy_in               =>      gt17_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt17_txusrclk_in                =>      gt17_txusrclk_i,
        gt17_txusrclk2_in               =>      gt17_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt17_txdata_in                  =>      gt17_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt17_gthtxn_out                 =>      gt17_gthtxn_out,
        gt17_gthtxp_out                 =>      gt17_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt17_txoutclk_out               =>      gt17_txoutclk_i,
        gt17_txoutclkfabric_out         =>      gt17_txoutclkfabric_out,
        gt17_txoutclkpcs_out            =>      gt17_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt17_txresetdone_out            =>      gt17_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt17_txcharisk_in               =>      gt17_txcharisk_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT18  (X1Y22)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt18_drpaddr_in                 =>      gt18_drpaddr_in,
        gt18_drpclk_in                  =>      sysclk_in_i,
        gt18_drpdi_in                   =>      gt18_drpdi_in,
        gt18_drpdo_out                  =>      gt18_drpdo_out,
        gt18_drpen_in                   =>      gt18_drpen_in,
        gt18_drprdy_out                 =>      gt18_drprdy_out,
        gt18_drpwe_in                   =>      gt18_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt18_eyescanreset_in            =>      gt18_eyescanreset_in,
        gt18_rxuserrdy_in               =>      gt18_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt18_eyescandataerror_out       =>      gt18_eyescandataerror_out,
        gt18_eyescantrigger_in          =>      gt18_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt18_rxslide_in                 =>      gt18_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt18_dmonitorout_out            =>      gt18_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt18_rxusrclk_in                =>      gt18_rxusrclk_i,
        gt18_rxusrclk2_in               =>      gt18_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt18_rxdata_out                 =>      gt18_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt18_rxdisperr_out              =>      gt18_rxdisperr_out,
        gt18_rxnotintable_out           =>      gt18_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt18_gthrxn_in                  =>      gt18_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt18_rxphmonitor_out            =>      gt18_rxphmonitor_out,
        gt18_rxphslipmonitor_out        =>      gt18_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt18_rxbyteisaligned_out        =>      gt18_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt18_rxmonitorout_out           =>      gt18_rxmonitorout_out,
        gt18_rxmonitorsel_in            =>      gt18_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt18_rxoutclk_out               =>      gt18_rxoutclk_i,
        gt18_rxoutclkfabric_out         =>      gt18_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt18_gtrxreset_in               =>      gt18_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt18_rxcharisk_out              =>      gt18_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt18_gthrxp_in                  =>      gt18_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt18_rxresetdone_out            =>      gt18_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt18_gttxreset_in               =>      gt18_gttxreset_in,
        gt18_txuserrdy_in               =>      gt18_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt18_txusrclk_in                =>      gt18_txusrclk_i,
        gt18_txusrclk2_in               =>      gt18_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt18_txdata_in                  =>      gt18_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt18_gthtxn_out                 =>      gt18_gthtxn_out,
        gt18_gthtxp_out                 =>      gt18_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt18_txoutclk_out               =>      gt18_txoutclk_i,
        gt18_txoutclkfabric_out         =>      gt18_txoutclkfabric_out,
        gt18_txoutclkpcs_out            =>      gt18_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt18_txresetdone_out            =>      gt18_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt18_txcharisk_in               =>      gt18_txcharisk_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT19  (X1Y23)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt19_drpaddr_in                 =>      gt19_drpaddr_in,
        gt19_drpclk_in                  =>      sysclk_in_i,
        gt19_drpdi_in                   =>      gt19_drpdi_in,
        gt19_drpdo_out                  =>      gt19_drpdo_out,
        gt19_drpen_in                   =>      gt19_drpen_in,
        gt19_drprdy_out                 =>      gt19_drprdy_out,
        gt19_drpwe_in                   =>      gt19_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt19_eyescanreset_in            =>      gt19_eyescanreset_in,
        gt19_rxuserrdy_in               =>      gt19_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt19_eyescandataerror_out       =>      gt19_eyescandataerror_out,
        gt19_eyescantrigger_in          =>      gt19_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt19_rxslide_in                 =>      gt19_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt19_dmonitorout_out            =>      gt19_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt19_rxusrclk_in                =>      gt19_rxusrclk_i,
        gt19_rxusrclk2_in               =>      gt19_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt19_rxdata_out                 =>      gt19_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt19_rxdisperr_out              =>      gt19_rxdisperr_out,
        gt19_rxnotintable_out           =>      gt19_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt19_gthrxn_in                  =>      gt19_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt19_rxphmonitor_out            =>      gt19_rxphmonitor_out,
        gt19_rxphslipmonitor_out        =>      gt19_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt19_rxbyteisaligned_out        =>      gt19_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt19_rxmonitorout_out           =>      gt19_rxmonitorout_out,
        gt19_rxmonitorsel_in            =>      gt19_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt19_rxoutclk_out               =>      gt19_rxoutclk_i,
        gt19_rxoutclkfabric_out         =>      gt19_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt19_gtrxreset_in               =>      gt19_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt19_rxcharisk_out              =>      gt19_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt19_gthrxp_in                  =>      gt19_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt19_rxresetdone_out            =>      gt19_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt19_gttxreset_in               =>      gt19_gttxreset_in,
        gt19_txuserrdy_in               =>      gt19_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt19_txusrclk_in                =>      gt19_txusrclk_i,
        gt19_txusrclk2_in               =>      gt19_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt19_txdata_in                  =>      gt19_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt19_gthtxn_out                 =>      gt19_gthtxn_out,
        gt19_gthtxp_out                 =>      gt19_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt19_txoutclk_out               =>      gt19_txoutclk_i,
        gt19_txoutclkfabric_out         =>      gt19_txoutclkfabric_out,
        gt19_txoutclkpcs_out            =>      gt19_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt19_txresetdone_out            =>      gt19_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt19_txcharisk_in               =>      gt19_txcharisk_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT20  (X1Y24)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt20_drpaddr_in                 =>      gt20_drpaddr_in,
        gt20_drpclk_in                  =>      sysclk_in_i,
        gt20_drpdi_in                   =>      gt20_drpdi_in,
        gt20_drpdo_out                  =>      gt20_drpdo_out,
        gt20_drpen_in                   =>      gt20_drpen_in,
        gt20_drprdy_out                 =>      gt20_drprdy_out,
        gt20_drpwe_in                   =>      gt20_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt20_eyescanreset_in            =>      gt20_eyescanreset_in,
        gt20_rxuserrdy_in               =>      gt20_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt20_eyescandataerror_out       =>      gt20_eyescandataerror_out,
        gt20_eyescantrigger_in          =>      gt20_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt20_rxslide_in                 =>      gt20_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt20_dmonitorout_out            =>      gt20_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt20_rxusrclk_in                =>      gt20_rxusrclk_i,
        gt20_rxusrclk2_in               =>      gt20_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt20_rxdata_out                 =>      gt20_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt20_rxdisperr_out              =>      gt20_rxdisperr_out,
        gt20_rxnotintable_out           =>      gt20_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt20_gthrxn_in                  =>      gt20_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt20_rxphmonitor_out            =>      gt20_rxphmonitor_out,
        gt20_rxphslipmonitor_out        =>      gt20_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt20_rxbyteisaligned_out        =>      gt20_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt20_rxmonitorout_out           =>      gt20_rxmonitorout_out,
        gt20_rxmonitorsel_in            =>      gt20_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt20_rxoutclk_out               =>      gt20_rxoutclk_i,
        gt20_rxoutclkfabric_out         =>      gt20_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt20_gtrxreset_in               =>      gt20_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt20_rxcharisk_out              =>      gt20_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt20_gthrxp_in                  =>      gt20_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt20_rxresetdone_out            =>      gt20_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt20_gttxreset_in               =>      gt20_gttxreset_in,
        gt20_txuserrdy_in               =>      gt20_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt20_txusrclk_in                =>      gt20_txusrclk_i,
        gt20_txusrclk2_in               =>      gt20_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt20_txdata_in                  =>      gt20_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt20_gthtxn_out                 =>      gt20_gthtxn_out,
        gt20_gthtxp_out                 =>      gt20_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt20_txoutclk_out               =>      gt20_txoutclk_i,
        gt20_txoutclkfabric_out         =>      gt20_txoutclkfabric_out,
        gt20_txoutclkpcs_out            =>      gt20_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt20_txresetdone_out            =>      gt20_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt20_txcharisk_in               =>      gt20_txcharisk_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT21  (X1Y25)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt21_drpaddr_in                 =>      gt21_drpaddr_in,
        gt21_drpclk_in                  =>      sysclk_in_i,
        gt21_drpdi_in                   =>      gt21_drpdi_in,
        gt21_drpdo_out                  =>      gt21_drpdo_out,
        gt21_drpen_in                   =>      gt21_drpen_in,
        gt21_drprdy_out                 =>      gt21_drprdy_out,
        gt21_drpwe_in                   =>      gt21_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt21_eyescanreset_in            =>      gt21_eyescanreset_in,
        gt21_rxuserrdy_in               =>      gt21_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt21_eyescandataerror_out       =>      gt21_eyescandataerror_out,
        gt21_eyescantrigger_in          =>      gt21_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt21_rxslide_in                 =>      gt21_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt21_dmonitorout_out            =>      gt21_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt21_rxusrclk_in                =>      gt21_rxusrclk_i,
        gt21_rxusrclk2_in               =>      gt21_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt21_rxdata_out                 =>      gt21_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt21_rxdisperr_out              =>      gt21_rxdisperr_out,
        gt21_rxnotintable_out           =>      gt21_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt21_gthrxn_in                  =>      gt21_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt21_rxphmonitor_out            =>      gt21_rxphmonitor_out,
        gt21_rxphslipmonitor_out        =>      gt21_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt21_rxbyteisaligned_out        =>      gt21_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt21_rxmonitorout_out           =>      gt21_rxmonitorout_out,
        gt21_rxmonitorsel_in            =>      gt21_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt21_rxoutclk_out               =>      gt21_rxoutclk_i,
        gt21_rxoutclkfabric_out         =>      gt21_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt21_gtrxreset_in               =>      gt21_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt21_rxcharisk_out              =>      gt21_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt21_gthrxp_in                  =>      gt21_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt21_rxresetdone_out            =>      gt21_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt21_gttxreset_in               =>      gt21_gttxreset_in,
        gt21_txuserrdy_in               =>      gt21_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt21_txusrclk_in                =>      gt21_txusrclk_i,
        gt21_txusrclk2_in               =>      gt21_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt21_txdata_in                  =>      gt21_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt21_gthtxn_out                 =>      gt21_gthtxn_out,
        gt21_gthtxp_out                 =>      gt21_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt21_txoutclk_out               =>      gt21_txoutclk_i,
        gt21_txoutclkfabric_out         =>      gt21_txoutclkfabric_out,
        gt21_txoutclkpcs_out            =>      gt21_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt21_txresetdone_out            =>      gt21_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt21_txcharisk_in               =>      gt21_txcharisk_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT22  (X1Y26)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt22_drpaddr_in                 =>      gt22_drpaddr_in,
        gt22_drpclk_in                  =>      sysclk_in_i,
        gt22_drpdi_in                   =>      gt22_drpdi_in,
        gt22_drpdo_out                  =>      gt22_drpdo_out,
        gt22_drpen_in                   =>      gt22_drpen_in,
        gt22_drprdy_out                 =>      gt22_drprdy_out,
        gt22_drpwe_in                   =>      gt22_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt22_eyescanreset_in            =>      gt22_eyescanreset_in,
        gt22_rxuserrdy_in               =>      gt22_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt22_eyescandataerror_out       =>      gt22_eyescandataerror_out,
        gt22_eyescantrigger_in          =>      gt22_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt22_rxslide_in                 =>      gt22_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt22_dmonitorout_out            =>      gt22_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt22_rxusrclk_in                =>      gt22_rxusrclk_i,
        gt22_rxusrclk2_in               =>      gt22_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt22_rxdata_out                 =>      gt22_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt22_rxdisperr_out              =>      gt22_rxdisperr_out,
        gt22_rxnotintable_out           =>      gt22_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt22_gthrxn_in                  =>      gt22_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt22_rxphmonitor_out            =>      gt22_rxphmonitor_out,
        gt22_rxphslipmonitor_out        =>      gt22_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt22_rxbyteisaligned_out        =>      gt22_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt22_rxmonitorout_out           =>      gt22_rxmonitorout_out,
        gt22_rxmonitorsel_in            =>      gt22_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt22_rxoutclk_out               =>      gt22_rxoutclk_i,
        gt22_rxoutclkfabric_out         =>      gt22_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt22_gtrxreset_in               =>      gt22_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt22_rxcharisk_out              =>      gt22_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt22_gthrxp_in                  =>      gt22_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt22_rxresetdone_out            =>      gt22_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt22_gttxreset_in               =>      gt22_gttxreset_in,
        gt22_txuserrdy_in               =>      gt22_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt22_txusrclk_in                =>      gt22_txusrclk_i,
        gt22_txusrclk2_in               =>      gt22_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt22_txdata_in                  =>      gt22_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt22_gthtxn_out                 =>      gt22_gthtxn_out,
        gt22_gthtxp_out                 =>      gt22_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt22_txoutclk_out               =>      gt22_txoutclk_i,
        gt22_txoutclkfabric_out         =>      gt22_txoutclkfabric_out,
        gt22_txoutclkpcs_out            =>      gt22_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt22_txresetdone_out            =>      gt22_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt22_txcharisk_in               =>      gt22_txcharisk_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT23  (X1Y27)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt23_drpaddr_in                 =>      gt23_drpaddr_in,
        gt23_drpclk_in                  =>      sysclk_in_i,
        gt23_drpdi_in                   =>      gt23_drpdi_in,
        gt23_drpdo_out                  =>      gt23_drpdo_out,
        gt23_drpen_in                   =>      gt23_drpen_in,
        gt23_drprdy_out                 =>      gt23_drprdy_out,
        gt23_drpwe_in                   =>      gt23_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt23_eyescanreset_in            =>      gt23_eyescanreset_in,
        gt23_rxuserrdy_in               =>      gt23_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt23_eyescandataerror_out       =>      gt23_eyescandataerror_out,
        gt23_eyescantrigger_in          =>      gt23_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt23_rxslide_in                 =>      gt23_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt23_dmonitorout_out            =>      gt23_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt23_rxusrclk_in                =>      gt23_rxusrclk_i,
        gt23_rxusrclk2_in               =>      gt23_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt23_rxdata_out                 =>      gt23_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt23_rxdisperr_out              =>      gt23_rxdisperr_out,
        gt23_rxnotintable_out           =>      gt23_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt23_gthrxn_in                  =>      gt23_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt23_rxphmonitor_out            =>      gt23_rxphmonitor_out,
        gt23_rxphslipmonitor_out        =>      gt23_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt23_rxbyteisaligned_out        =>      gt23_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt23_rxmonitorout_out           =>      gt23_rxmonitorout_out,
        gt23_rxmonitorsel_in            =>      gt23_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt23_rxoutclk_out               =>      gt23_rxoutclk_i,
        gt23_rxoutclkfabric_out         =>      gt23_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt23_gtrxreset_in               =>      gt23_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt23_rxcharisk_out              =>      gt23_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt23_gthrxp_in                  =>      gt23_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt23_rxresetdone_out            =>      gt23_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt23_gttxreset_in               =>      gt23_gttxreset_in,
        gt23_txuserrdy_in               =>      gt23_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt23_txusrclk_in                =>      gt23_txusrclk_i,
        gt23_txusrclk2_in               =>      gt23_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt23_txdata_in                  =>      gt23_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt23_gthtxn_out                 =>      gt23_gthtxn_out,
        gt23_gthtxp_out                 =>      gt23_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt23_txoutclk_out               =>      gt23_txoutclk_i,
        gt23_txoutclkfabric_out         =>      gt23_txoutclkfabric_out,
        gt23_txoutclkpcs_out            =>      gt23_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt23_txresetdone_out            =>      gt23_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt23_txcharisk_in               =>      gt23_txcharisk_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT24  (X1Y28)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt24_drpaddr_in                 =>      gt24_drpaddr_in,
        gt24_drpclk_in                  =>      sysclk_in_i,
        gt24_drpdi_in                   =>      gt24_drpdi_in,
        gt24_drpdo_out                  =>      gt24_drpdo_out,
        gt24_drpen_in                   =>      gt24_drpen_in,
        gt24_drprdy_out                 =>      gt24_drprdy_out,
        gt24_drpwe_in                   =>      gt24_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt24_eyescanreset_in            =>      gt24_eyescanreset_in,
        gt24_rxuserrdy_in               =>      gt24_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt24_eyescandataerror_out       =>      gt24_eyescandataerror_out,
        gt24_eyescantrigger_in          =>      gt24_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt24_rxslide_in                 =>      gt24_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt24_dmonitorout_out            =>      gt24_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt24_rxusrclk_in                =>      gt24_rxusrclk_i,
        gt24_rxusrclk2_in               =>      gt24_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt24_rxdata_out                 =>      gt24_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt24_rxdisperr_out              =>      gt24_rxdisperr_out,
        gt24_rxnotintable_out           =>      gt24_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt24_gthrxn_in                  =>      gt24_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt24_rxphmonitor_out            =>      gt24_rxphmonitor_out,
        gt24_rxphslipmonitor_out        =>      gt24_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt24_rxbyteisaligned_out        =>      gt24_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt24_rxmonitorout_out           =>      gt24_rxmonitorout_out,
        gt24_rxmonitorsel_in            =>      gt24_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt24_rxoutclk_out               =>      gt24_rxoutclk_i,
        gt24_rxoutclkfabric_out         =>      gt24_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt24_gtrxreset_in               =>      gt24_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt24_rxcharisk_out              =>      gt24_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt24_gthrxp_in                  =>      gt24_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt24_rxresetdone_out            =>      gt24_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt24_gttxreset_in               =>      gt24_gttxreset_in,
        gt24_txuserrdy_in               =>      gt24_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt24_txusrclk_in                =>      gt24_txusrclk_i,
        gt24_txusrclk2_in               =>      gt24_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt24_txdata_in                  =>      gt24_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt24_gthtxn_out                 =>      gt24_gthtxn_out,
        gt24_gthtxp_out                 =>      gt24_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt24_txoutclk_out               =>      gt24_txoutclk_i,
        gt24_txoutclkfabric_out         =>      gt24_txoutclkfabric_out,
        gt24_txoutclkpcs_out            =>      gt24_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt24_txresetdone_out            =>      gt24_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt24_txcharisk_in               =>      gt24_txcharisk_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT25  (X1Y29)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt25_drpaddr_in                 =>      gt25_drpaddr_in,
        gt25_drpclk_in                  =>      sysclk_in_i,
        gt25_drpdi_in                   =>      gt25_drpdi_in,
        gt25_drpdo_out                  =>      gt25_drpdo_out,
        gt25_drpen_in                   =>      gt25_drpen_in,
        gt25_drprdy_out                 =>      gt25_drprdy_out,
        gt25_drpwe_in                   =>      gt25_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt25_eyescanreset_in            =>      gt25_eyescanreset_in,
        gt25_rxuserrdy_in               =>      gt25_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt25_eyescandataerror_out       =>      gt25_eyescandataerror_out,
        gt25_eyescantrigger_in          =>      gt25_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt25_rxslide_in                 =>      gt25_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt25_dmonitorout_out            =>      gt25_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt25_rxusrclk_in                =>      gt25_rxusrclk_i,
        gt25_rxusrclk2_in               =>      gt25_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt25_rxdata_out                 =>      gt25_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt25_rxdisperr_out              =>      gt25_rxdisperr_out,
        gt25_rxnotintable_out           =>      gt25_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt25_gthrxn_in                  =>      gt25_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt25_rxphmonitor_out            =>      gt25_rxphmonitor_out,
        gt25_rxphslipmonitor_out        =>      gt25_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt25_rxbyteisaligned_out        =>      gt25_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt25_rxmonitorout_out           =>      gt25_rxmonitorout_out,
        gt25_rxmonitorsel_in            =>      gt25_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt25_rxoutclk_out               =>      gt25_rxoutclk_i,
        gt25_rxoutclkfabric_out         =>      gt25_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt25_gtrxreset_in               =>      gt25_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt25_rxcharisk_out              =>      gt25_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt25_gthrxp_in                  =>      gt25_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt25_rxresetdone_out            =>      gt25_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt25_gttxreset_in               =>      gt25_gttxreset_in,
        gt25_txuserrdy_in               =>      gt25_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt25_txusrclk_in                =>      gt25_txusrclk_i,
        gt25_txusrclk2_in               =>      gt25_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt25_txdata_in                  =>      gt25_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt25_gthtxn_out                 =>      gt25_gthtxn_out,
        gt25_gthtxp_out                 =>      gt25_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt25_txoutclk_out               =>      gt25_txoutclk_i,
        gt25_txoutclkfabric_out         =>      gt25_txoutclkfabric_out,
        gt25_txoutclkpcs_out            =>      gt25_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt25_txresetdone_out            =>      gt25_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt25_txcharisk_in               =>      gt25_txcharisk_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT26  (X1Y30)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt26_drpaddr_in                 =>      gt26_drpaddr_in,
        gt26_drpclk_in                  =>      sysclk_in_i,
        gt26_drpdi_in                   =>      gt26_drpdi_in,
        gt26_drpdo_out                  =>      gt26_drpdo_out,
        gt26_drpen_in                   =>      gt26_drpen_in,
        gt26_drprdy_out                 =>      gt26_drprdy_out,
        gt26_drpwe_in                   =>      gt26_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt26_eyescanreset_in            =>      gt26_eyescanreset_in,
        gt26_rxuserrdy_in               =>      gt26_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt26_eyescandataerror_out       =>      gt26_eyescandataerror_out,
        gt26_eyescantrigger_in          =>      gt26_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt26_rxslide_in                 =>      gt26_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt26_dmonitorout_out            =>      gt26_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt26_rxusrclk_in                =>      gt26_rxusrclk_i,
        gt26_rxusrclk2_in               =>      gt26_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt26_rxdata_out                 =>      gt26_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt26_rxdisperr_out              =>      gt26_rxdisperr_out,
        gt26_rxnotintable_out           =>      gt26_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt26_gthrxn_in                  =>      gt26_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt26_rxphmonitor_out            =>      gt26_rxphmonitor_out,
        gt26_rxphslipmonitor_out        =>      gt26_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt26_rxbyteisaligned_out        =>      gt26_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt26_rxmonitorout_out           =>      gt26_rxmonitorout_out,
        gt26_rxmonitorsel_in            =>      gt26_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt26_rxoutclk_out               =>      gt26_rxoutclk_i,
        gt26_rxoutclkfabric_out         =>      gt26_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt26_gtrxreset_in               =>      gt26_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt26_rxcharisk_out              =>      gt26_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt26_gthrxp_in                  =>      gt26_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt26_rxresetdone_out            =>      gt26_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt26_gttxreset_in               =>      gt26_gttxreset_in,
        gt26_txuserrdy_in               =>      gt26_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt26_txusrclk_in                =>      gt26_txusrclk_i,
        gt26_txusrclk2_in               =>      gt26_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt26_txdata_in                  =>      gt26_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt26_gthtxn_out                 =>      gt26_gthtxn_out,
        gt26_gthtxp_out                 =>      gt26_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt26_txoutclk_out               =>      gt26_txoutclk_i,
        gt26_txoutclkfabric_out         =>      gt26_txoutclkfabric_out,
        gt26_txoutclkpcs_out            =>      gt26_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt26_txresetdone_out            =>      gt26_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt26_txcharisk_in               =>      gt26_txcharisk_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT27  (X1Y31)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt27_drpaddr_in                 =>      gt27_drpaddr_in,
        gt27_drpclk_in                  =>      sysclk_in_i,
        gt27_drpdi_in                   =>      gt27_drpdi_in,
        gt27_drpdo_out                  =>      gt27_drpdo_out,
        gt27_drpen_in                   =>      gt27_drpen_in,
        gt27_drprdy_out                 =>      gt27_drprdy_out,
        gt27_drpwe_in                   =>      gt27_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt27_eyescanreset_in            =>      gt27_eyescanreset_in,
        gt27_rxuserrdy_in               =>      gt27_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt27_eyescandataerror_out       =>      gt27_eyescandataerror_out,
        gt27_eyescantrigger_in          =>      gt27_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt27_rxslide_in                 =>      gt27_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt27_dmonitorout_out            =>      gt27_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt27_rxusrclk_in                =>      gt27_rxusrclk_i,
        gt27_rxusrclk2_in               =>      gt27_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt27_rxdata_out                 =>      gt27_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt27_rxdisperr_out              =>      gt27_rxdisperr_out,
        gt27_rxnotintable_out           =>      gt27_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt27_gthrxn_in                  =>      gt27_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt27_rxphmonitor_out            =>      gt27_rxphmonitor_out,
        gt27_rxphslipmonitor_out        =>      gt27_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt27_rxbyteisaligned_out        =>      gt27_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt27_rxmonitorout_out           =>      gt27_rxmonitorout_out,
        gt27_rxmonitorsel_in            =>      gt27_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt27_rxoutclk_out               =>      gt27_rxoutclk_i,
        gt27_rxoutclkfabric_out         =>      gt27_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt27_gtrxreset_in               =>      gt27_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt27_rxcharisk_out              =>      gt27_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt27_gthrxp_in                  =>      gt27_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt27_rxresetdone_out            =>      gt27_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt27_gttxreset_in               =>      gt27_gttxreset_in,
        gt27_txuserrdy_in               =>      gt27_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt27_txusrclk_in                =>      gt27_txusrclk_i,
        gt27_txusrclk2_in               =>      gt27_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt27_txdata_in                  =>      gt27_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt27_gthtxn_out                 =>      gt27_gthtxn_out,
        gt27_gthtxp_out                 =>      gt27_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt27_txoutclk_out               =>      gt27_txoutclk_i,
        gt27_txoutclkfabric_out         =>      gt27_txoutclkfabric_out,
        gt27_txoutclkpcs_out            =>      gt27_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt27_txresetdone_out            =>      gt27_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt27_txcharisk_in               =>      gt27_txcharisk_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT28  (X1Y32)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt28_drpaddr_in                 =>      gt28_drpaddr_in,
        gt28_drpclk_in                  =>      sysclk_in_i,
        gt28_drpdi_in                   =>      gt28_drpdi_in,
        gt28_drpdo_out                  =>      gt28_drpdo_out,
        gt28_drpen_in                   =>      gt28_drpen_in,
        gt28_drprdy_out                 =>      gt28_drprdy_out,
        gt28_drpwe_in                   =>      gt28_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt28_eyescanreset_in            =>      gt28_eyescanreset_in,
        gt28_rxuserrdy_in               =>      gt28_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt28_eyescandataerror_out       =>      gt28_eyescandataerror_out,
        gt28_eyescantrigger_in          =>      gt28_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt28_rxslide_in                 =>      gt28_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt28_dmonitorout_out            =>      gt28_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt28_rxusrclk_in                =>      gt28_rxusrclk_i,
        gt28_rxusrclk2_in               =>      gt28_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt28_rxdata_out                 =>      gt28_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt28_rxdisperr_out              =>      gt28_rxdisperr_out,
        gt28_rxnotintable_out           =>      gt28_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt28_gthrxn_in                  =>      gt28_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt28_rxphmonitor_out            =>      gt28_rxphmonitor_out,
        gt28_rxphslipmonitor_out        =>      gt28_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt28_rxbyteisaligned_out        =>      gt28_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt28_rxmonitorout_out           =>      gt28_rxmonitorout_out,
        gt28_rxmonitorsel_in            =>      gt28_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt28_rxoutclk_out               =>      gt28_rxoutclk_i,
        gt28_rxoutclkfabric_out         =>      gt28_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt28_gtrxreset_in               =>      gt28_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt28_rxcharisk_out              =>      gt28_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt28_gthrxp_in                  =>      gt28_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt28_rxresetdone_out            =>      gt28_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt28_gttxreset_in               =>      gt28_gttxreset_in,
        gt28_txuserrdy_in               =>      gt28_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt28_txusrclk_in                =>      gt28_txusrclk_i,
        gt28_txusrclk2_in               =>      gt28_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt28_txdata_in                  =>      gt28_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt28_gthtxn_out                 =>      gt28_gthtxn_out,
        gt28_gthtxp_out                 =>      gt28_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt28_txoutclk_out               =>      gt28_txoutclk_i,
        gt28_txoutclkfabric_out         =>      gt28_txoutclkfabric_out,
        gt28_txoutclkpcs_out            =>      gt28_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt28_txresetdone_out            =>      gt28_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt28_txcharisk_in               =>      gt28_txcharisk_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT29  (X1Y33)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt29_drpaddr_in                 =>      gt29_drpaddr_in,
        gt29_drpclk_in                  =>      sysclk_in_i,
        gt29_drpdi_in                   =>      gt29_drpdi_in,
        gt29_drpdo_out                  =>      gt29_drpdo_out,
        gt29_drpen_in                   =>      gt29_drpen_in,
        gt29_drprdy_out                 =>      gt29_drprdy_out,
        gt29_drpwe_in                   =>      gt29_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt29_eyescanreset_in            =>      gt29_eyescanreset_in,
        gt29_rxuserrdy_in               =>      gt29_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt29_eyescandataerror_out       =>      gt29_eyescandataerror_out,
        gt29_eyescantrigger_in          =>      gt29_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt29_rxslide_in                 =>      gt29_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt29_dmonitorout_out            =>      gt29_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt29_rxusrclk_in                =>      gt29_rxusrclk_i,
        gt29_rxusrclk2_in               =>      gt29_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt29_rxdata_out                 =>      gt29_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt29_rxdisperr_out              =>      gt29_rxdisperr_out,
        gt29_rxnotintable_out           =>      gt29_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt29_gthrxn_in                  =>      gt29_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt29_rxphmonitor_out            =>      gt29_rxphmonitor_out,
        gt29_rxphslipmonitor_out        =>      gt29_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt29_rxbyteisaligned_out        =>      gt29_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt29_rxmonitorout_out           =>      gt29_rxmonitorout_out,
        gt29_rxmonitorsel_in            =>      gt29_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt29_rxoutclk_out               =>      gt29_rxoutclk_i,
        gt29_rxoutclkfabric_out         =>      gt29_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt29_gtrxreset_in               =>      gt29_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt29_rxcharisk_out              =>      gt29_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt29_gthrxp_in                  =>      gt29_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt29_rxresetdone_out            =>      gt29_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt29_gttxreset_in               =>      gt29_gttxreset_in,
        gt29_txuserrdy_in               =>      gt29_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt29_txusrclk_in                =>      gt29_txusrclk_i,
        gt29_txusrclk2_in               =>      gt29_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt29_txdata_in                  =>      gt29_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt29_gthtxn_out                 =>      gt29_gthtxn_out,
        gt29_gthtxp_out                 =>      gt29_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt29_txoutclk_out               =>      gt29_txoutclk_i,
        gt29_txoutclkfabric_out         =>      gt29_txoutclkfabric_out,
        gt29_txoutclkpcs_out            =>      gt29_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt29_txresetdone_out            =>      gt29_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt29_txcharisk_in               =>      gt29_txcharisk_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT30  (X1Y34)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt30_drpaddr_in                 =>      gt30_drpaddr_in,
        gt30_drpclk_in                  =>      sysclk_in_i,
        gt30_drpdi_in                   =>      gt30_drpdi_in,
        gt30_drpdo_out                  =>      gt30_drpdo_out,
        gt30_drpen_in                   =>      gt30_drpen_in,
        gt30_drprdy_out                 =>      gt30_drprdy_out,
        gt30_drpwe_in                   =>      gt30_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt30_eyescanreset_in            =>      gt30_eyescanreset_in,
        gt30_rxuserrdy_in               =>      gt30_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt30_eyescandataerror_out       =>      gt30_eyescandataerror_out,
        gt30_eyescantrigger_in          =>      gt30_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt30_rxslide_in                 =>      gt30_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt30_dmonitorout_out            =>      gt30_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt30_rxusrclk_in                =>      gt30_rxusrclk_i,
        gt30_rxusrclk2_in               =>      gt30_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt30_rxdata_out                 =>      gt30_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt30_rxdisperr_out              =>      gt30_rxdisperr_out,
        gt30_rxnotintable_out           =>      gt30_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt30_gthrxn_in                  =>      gt30_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt30_rxphmonitor_out            =>      gt30_rxphmonitor_out,
        gt30_rxphslipmonitor_out        =>      gt30_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt30_rxbyteisaligned_out        =>      gt30_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt30_rxmonitorout_out           =>      gt30_rxmonitorout_out,
        gt30_rxmonitorsel_in            =>      gt30_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt30_rxoutclk_out               =>      gt30_rxoutclk_i,
        gt30_rxoutclkfabric_out         =>      gt30_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt30_gtrxreset_in               =>      gt30_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt30_rxcharisk_out              =>      gt30_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt30_gthrxp_in                  =>      gt30_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt30_rxresetdone_out            =>      gt30_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt30_gttxreset_in               =>      gt30_gttxreset_in,
        gt30_txuserrdy_in               =>      gt30_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt30_txusrclk_in                =>      gt30_txusrclk_i,
        gt30_txusrclk2_in               =>      gt30_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt30_txdata_in                  =>      gt30_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt30_gthtxn_out                 =>      gt30_gthtxn_out,
        gt30_gthtxp_out                 =>      gt30_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt30_txoutclk_out               =>      gt30_txoutclk_i,
        gt30_txoutclkfabric_out         =>      gt30_txoutclkfabric_out,
        gt30_txoutclkpcs_out            =>      gt30_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt30_txresetdone_out            =>      gt30_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt30_txcharisk_in               =>      gt30_txcharisk_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT31  (X1Y35)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt31_drpaddr_in                 =>      gt31_drpaddr_in,
        gt31_drpclk_in                  =>      sysclk_in_i,
        gt31_drpdi_in                   =>      gt31_drpdi_in,
        gt31_drpdo_out                  =>      gt31_drpdo_out,
        gt31_drpen_in                   =>      gt31_drpen_in,
        gt31_drprdy_out                 =>      gt31_drprdy_out,
        gt31_drpwe_in                   =>      gt31_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt31_eyescanreset_in            =>      gt31_eyescanreset_in,
        gt31_rxuserrdy_in               =>      gt31_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt31_eyescandataerror_out       =>      gt31_eyescandataerror_out,
        gt31_eyescantrigger_in          =>      gt31_eyescantrigger_in,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        gt31_rxslide_in                 =>      gt31_rxslide_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt31_dmonitorout_out            =>      gt31_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt31_rxusrclk_in                =>      gt31_rxusrclk_i,
        gt31_rxusrclk2_in               =>      gt31_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt31_rxdata_out                 =>      gt31_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt31_rxdisperr_out              =>      gt31_rxdisperr_out,
        gt31_rxnotintable_out           =>      gt31_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt31_gthrxn_in                  =>      gt31_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt31_rxphmonitor_out            =>      gt31_rxphmonitor_out,
        gt31_rxphslipmonitor_out        =>      gt31_rxphslipmonitor_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt31_rxbyteisaligned_out        =>      gt31_rxbyteisaligned_out,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt31_rxmonitorout_out           =>      gt31_rxmonitorout_out,
        gt31_rxmonitorsel_in            =>      gt31_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt31_rxoutclk_out               =>      gt31_rxoutclk_i,
        gt31_rxoutclkfabric_out         =>      gt31_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt31_gtrxreset_in               =>      gt31_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt31_rxcharisk_out              =>      gt31_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt31_gthrxp_in                  =>      gt31_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt31_rxresetdone_out            =>      gt31_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt31_gttxreset_in               =>      gt31_gttxreset_in,
        gt31_txuserrdy_in               =>      gt31_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt31_txusrclk_in                =>      gt31_txusrclk_i,
        gt31_txusrclk2_in               =>      gt31_txusrclk2_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt31_txdata_in                  =>      gt31_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt31_gthtxn_out                 =>      gt31_gthtxn_out,
        gt31_gthtxp_out                 =>      gt31_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt31_txoutclk_out               =>      gt31_txoutclk_i,
        gt31_txoutclkfabric_out         =>      gt31_txoutclkfabric_out,
        gt31_txoutclkpcs_out            =>      gt31_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt31_txresetdone_out            =>      gt31_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt31_txcharisk_in               =>      gt31_txcharisk_in,



    gt0_qplllock_in => gt0_qplllock_i,
    gt0_qpllrefclklost_in => gt0_qpllrefclklost_i,
    gt0_qpllreset_out => gt0_qpllreset_i,
    gt0_qplloutclk_in => gt0_qplloutclk_i,
    gt0_qplloutrefclk_in => gt0_qplloutrefclk_i,
    gt1_qplllock_in => gt1_qplllock_i,
    gt1_qpllrefclklost_in => gt1_qpllrefclklost_i,
    gt1_qpllreset_out => gt1_qpllreset_i,
    gt1_qplloutclk_in => gt1_qplloutclk_i,
    gt1_qplloutrefclk_in => gt1_qplloutrefclk_i,
    gt2_qplllock_in => gt2_qplllock_i,
    gt2_qpllrefclklost_in => gt2_qpllrefclklost_i,
    gt2_qpllreset_out => gt2_qpllreset_i,
    gt2_qplloutclk_in => gt2_qplloutclk_i,
    gt2_qplloutrefclk_in => gt2_qplloutrefclk_i,
    gt3_qplllock_in => gt3_qplllock_i,
    gt3_qpllrefclklost_in => gt3_qpllrefclklost_i,
    gt3_qpllreset_out => gt3_qpllreset_i,
    gt3_qplloutclk_in => gt3_qplloutclk_i,
    gt3_qplloutrefclk_in => gt3_qplloutrefclk_i,
    gt4_qplllock_in => gt4_qplllock_i,
    gt4_qpllrefclklost_in => gt4_qpllrefclklost_i,
    gt4_qpllreset_out => gt4_qpllreset_i,
    gt4_qplloutclk_in => gt4_qplloutclk_i,
    gt4_qplloutrefclk_in => gt4_qplloutrefclk_i,
    gt5_qplllock_in => gt5_qplllock_i,
    gt5_qpllrefclklost_in => gt5_qpllrefclklost_i,
    gt5_qpllreset_out => gt5_qpllreset_i,
    gt5_qplloutclk_in => gt5_qplloutclk_i,
    gt5_qplloutrefclk_in => gt5_qplloutrefclk_i,
    gt6_qplllock_in => gt6_qplllock_i,
    gt6_qpllrefclklost_in => gt6_qpllrefclklost_i,
    gt6_qpllreset_out => gt6_qpllreset_i,
    gt6_qplloutclk_in => gt6_qplloutclk_i,
    gt6_qplloutrefclk_in => gt6_qplloutrefclk_i,
    gt7_qplllock_in => gt7_qplllock_i,
    gt7_qpllrefclklost_in => gt7_qpllrefclklost_i,
    gt7_qpllreset_out => gt7_qpllreset_i,
    gt7_qplloutclk_in => gt7_qplloutclk_i,
    gt7_qplloutrefclk_in => gt7_qplloutrefclk_i
    );



end RTL;
