

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EeIOalsB9A7gyFzgjBZExeIPJuRpFELHlfpU3L/uqPMoO6TuIez2KobOfgsxw4FitpHwSA97/lIN
csNqzUP09g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hwzf6tFLlGdH/LlAouRRMzleWlGs8Tvfr64AeA2s2z4reQzhfo3uL+7NKshrdnE3tMEN66HYuwVd
9xQlnCboKstjE9oTcxVT1Q9+i6ynCWa3yDpjnUvWm0p5bbxLnANX37Tx0FTTAfpo8DSKKm9W9UkH
5GCk1+VjPB9HCpd9nRE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bL2EnncrNSLn2ffq1uLRkntupOO+jbrSmLJY+5LxOcioiLBdds86PhRnmpvnUOMHuvC456xH0laA
GUJu8mYWsLkeJ/gjFzllQcWIPJ8fmH+TDnW5/yyAde/a0JpR0BbhVMzIYr60Z0Rs9B0t212q0Gi5
cfOdS9LTaW5pBjCKt0jNfdZ8Lr4AQUDsXpboqkvDmK3/+QJqqF7qvFtia5MvW70KQywr5vkgRws1
BASbR4GzizLUz3PzW0ZpTpLs/v+rps64Cwqc+09rCJXCFOqMTOnvf26vB8oglq7BMh6zBeWRxEuP
co0bzIox5OWgSFlu3oTH0cogMWKub8qQURYsWA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cIw/9EXCGVcaeoMMOWuYgFWlA9RUYNad2DCpvqx230raBxPvQNhdOwE34j858OOUuWrDVHLj1nWJ
y5EJbcyT1Tah86TN1vYqo8sqn5YXS+1zRWIej0AYDEi19T5qjqQjxcf11goih0I+aTjhgw55UIbx
DOlEcwyPrQQ1bBWTza7LH/J9VH+m0Nj/ooSJpuXCu3H7BNulUXfTKVRWBHnUEaUIRnumtCzfbcC9
ERqZzs4FrgS6flY1m9XbUdMT4p1Eo893HLMAHq10sTH6EHY/8n0KLkE0TdZ534HUCGr6KkB4RIDF
99mj7IvY4KQjySVBm3SLkgpins9y6UuDnCijkQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IcyVbDfeKPQ4Wv8Ubt7+Je8EyB4He+T9m7hctmPOEOS01haLEIPmxZJ+0X54mZvQdvPqdj7E23u1
R3OAzZqlLWLW+d0PIGnEownI+S9ocJwuizHj1sJuwEI4jfxmJNZjE4H7mK9ZjmgjaH4o48SdhJi2
yTDL4y4yJ9WH40IPNyPODb7zhqRTxClMXzjuJVpcO9fl61K8ntq/eG0XNZEJOUgYAk+JXVhPJ/R8
LP1drMB6yJI5AgR28Irm3VsSjJoMYUTX0eURD1i60OoVxl2DyucunlM5CIRZ9EHKoz5SjCNfLkmU
FtKjFd9bGHkZXD09XWdopli+1qzB7QvkJwZtJA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ApmmzO+E6sydVLZl1/2U7QnosCNZyxTsKqLSJRPek46QkWcHHZkNFVIHCIci4gSId93OhQssVzwz
WXxP3kwkA1nXIZbFYCJMBa9u+RSxeQycrHAglmUYWkuVydXtuVb2yoM2k+rwZmSZ4EL9o6DJBzpF
8rAtNuDZO+/14GwY/z8=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mLieXakPF5k1udgyxKQoGQOFSmNMp9LBLBSpMy1hh3mZegEUQzRC/x5AREnUXKCJVi2A45mQS+/v
sWYfEz/mEcmJNfzQRumZAzzIhT6OZ1BKHYHb35ddARKqGfi1VsbWUgVRiujIoWzcq/UVTRYREjX4
QTMnCGRVa9CTZ5zSpFRgcb6v/R9mln69hqjdTg41euhxw8cfIA1i23jDHJi3nWhqoyUvQDcLM9/8
Dyyt1tIBHV0Mj2Wh0eMPypOfqhIduKFcpK/XdxKtvUexe1DxPTzpolzVZLafUNx2epnjraWTb5kB
0Z5dogCBc3Gek9KtkaoCoZYrz7kpzUy4L2reXA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 129920)
`protect data_block
Yjp1IVfLVXlaXo6Hd49QAB4mjfoxzwNbMnhC6uCqZn7gZcEMyx5qoriI+zcQm29pCbhlArHaXGu1
oYReK4QAxMlMnr4h1M8A5awp9sI/gdopPXe6yxC4KndjHFdWme2ncNM0BT1AMvy1XQrlB0etn83j
e28ZYbAYgXneQx8TlN7FWHOD7qp7RvX0BYointNVHtBn1Q4tE4euHz8HB77zW8/hA+dKFOxaual5
/6DPYzNcy7XOa30noUnR+A/Eo3c9DCX/u3ZkefCUrJAeN/nqD01iPfJlBncSzBsmsOizaFiHZh85
XfoCVPCELbZcaYueckbdEdb6GW/lr8HWRlx0UnbweS0NaqJLYHrmzx407TNPnmcQr5m0WEy0khQI
6aws8q+p/RmsmLfHZh/hxI/tKvKtd2CZ8vUyvCaSspXsnUF0bUtVYh4nRLATt05ibjujqqN2pdeT
hbt+d8jOoepRvStISrFM6dqHDuLuKWfHq1Iz036GqZInKPzBl3gzaP9xMv9zaXlXbXWNzmpa5lhO
gKpjrUyt9UQ660BjVPEh1LKWUpBChSabRV5R92ionM3X39sWJB7SKDkK0Ybo4Fwu+p8LV44YD8WK
rgzdvznJvZWKQ3+/skbouw/XrU4ZH/kiQxOS7MC+pY+kAipgRn7egJFXBq3K5Xyp299wPG3Vde1L
zKQ/XPdxvVe11OJcpOLBbspjNmowuFe3qQeJaRulJscb1Vb9rDLxsLjiiag41th6Tpc7t37Ti3N/
EqZ1xx+Sa0ZhZnRnF9pFtg85F1bTbTgugGQJFD0MsY7lkrd2Avh3L+p56NEVj6r9V5gNaOHVa1nb
8fr1LnWKSQ7reMiT6PKL1703DVetmYD3gyhgxg3OrKWVvvxwRyfHh0CQYWj6pmE3njUQoIgklHII
TNx4o+BMJO1PmPsEkIMCB5XEg+FWRlb2n5YMywm7nXg0mPcIonwFBPsepeAGnTvOeLh4qVsXMa9U
7kurDF94Ce8Vlii6qzv/WtI1zYNu8nOgGE0wMoDNMef/DSeOGQEP5dFz1Comlki8Zs9glha2dAr2
REcch+xcmO5Z4RlVAxAjSgpdXZYNuRc6mrJZn039JeuzOn+Kyn5LGJtskM/FUnVIHPquqH9vN0WP
qJ7W8zYQuZjefGQHsq6m3OkB28nLZf16W1a24/Jw0GQgZ/8AQe309ti4lNn+DOGm41dHH2S74+dD
3+eEZnmOaTXiiy6cviyfoqIBRkkPjRrT5LjWUSahLjzeHCDpiIThwUPCPTI4UhCACos5pncsdqn9
lWg46U1niEJvm0/jLRbKa6fZ5OwLRt9imQTd/4ebLjjwVFC3vSLkWJyLDSOumKmqeCwRbimqxTH/
nmS2cbEu2/NSczL5CxtnlLam0F9hb73yeW2TqLobKjgKIuHkaP6PNR5JWr8zlnqSYY6wZpkOnL88
onocXdewafM/DGXPwi4sldTg3zGpRmDtGsl79ZsNjmqypZm6xVZl9CvSwRj9irQc2avleAiAPyqp
9EV5kh/ubIoJkprTPHglDnHWvm8ADPkvvXce6IjBN8Gy3Qe8HwN+h0hsK06Bg5YXepvxFK2Cthnb
OIJk3cqXi2piNj54DOsmuLW30N+bjN3XkhsX2ST5uIkEGkCAPpo0Zb0UL0Z/BbVpcgkFMTZ0trUW
SBGM4/zRV54o+6tblcba3LWdp1kOiSrktNzudbl1OHwOeTqudNa1sKpEBhUCMnjj8ObXwH9SKZ7w
eREGP514zeGVRKzc+Il5Jpp7llS8r4eg6Xd8k0VnNUKND8XBOX2IiHV8W4BDJw9iM52eRNOv63c2
nVD88X3+OnTx6Om0WTLwtOFRBaTFNFgVYWTaSNxKWI17ZwtCIEDheya6eendTHemFyS+5MAX8Jvc
3VGk4x4znimWlx/9SDpRXKA9qJoK2nDWsixQn5VnRj6Gx3qN5whqkEjNpxLJvjiPSDxRe1BdMOzF
nILJbuN0jPeectklYqGvg25iFCTk9cSRoaoiJagTAiuPalyf3/A7A9N5kioGzSQ5wuzRTCveMqk1
QOZCwuQJGK5dIvN/XSQSJd2F4C6wOy9nznNkSc+JgAIFIEHfrSZEzhvj0ycEHEeDUb9d4dzn0CW0
WtFliie7AnHotNbXWGODvPGk27abVzmR2URTs4xreKAryFW11vzQSMtkc51+OuXh1ra7PiAQJWfA
UmPaQ2Oks9wKdhBPz87o1KlEsRJ1UCrmekndc3wZzX6raUgZ+RWRl47+e7iTWZO10EAP0l4IpqEa
ZPwqK91/ib1CtpVA3CuV8nEwtPEKEkfJ6DnzcYu5gjPXm9YEGLdhvd8azsgLosTpnkYEgfEYjmwm
/LxddpL0Twm8G6N7k2ijlvdblVeQA88Nh931CWpS/mz5c63w6nSxWoMklK1EOhuAsIQbuZN6BrXU
iH6kHQH9sQcoTJ9Wd8oXAiBsr1OvJzi5/xXkMB1fNa2IETtPtn3udwo0fUkbMTuU43j4HGOgmpqR
lgStMejkCl5fVxiOF1DLhwo1/hONlHpsVKpkSXQ77Ypvc4LJSEXhf7+3VUU/OLzTzOFFjyhU3YMG
mEMttBCMUriyvZM0Z/dUizI79Dqv89gIZk4y6z/+EcgiOwEcDlkMLfv1Cb7bn6Pi8EcL7Z8Z8z3Y
y8gCHfImNz1nodZlUaWIVpA6eVRp6lB0E5gilEb7Rmx7iPm0OQWJmW67ZHmSQueec83p5Z+NGWWg
IRTRfutDQ1bDUaxUGPpwDSZ/f2xFiMqEYmrFEb1ZUFZ8IKq9dRBu1tdaOgHSHzARX1OqF8dHES9E
5cWFZvyDqqvtSUuMu57q88MQMKovPDeyEF3kI7i3KOCa92izpButu0y+H800ocD6gJJsdCdWvSmF
GMVZucI5Mnjbx16v3GGE8x97tEGuB+GcLxczh+yksokUD13VH2x0kuPjomYgIh6E9PbgM1npmpFN
QSVGod1tlNAtXzjEDF2xW/MEsr8fHtjAi8XiuZ+QnPRP7it8SH4ZzGbT1RC1QBofS/UAcO59amq0
eVwAEnTTrH7gkzcHHbO/HQpB6ib/Yv9oaac+vq+9WV8pFE/MOreF0Jb+XWCVLpK4K1s+X9B2ARBL
cWRycwFm6DFRoNoi4s6965hPmXfMraaTYF8jryfAe115q2D1FZ5mL8cGxm5oFOaig70j3rBVQfCT
EWtNrerfjBJQdpaHj0NfU25Wmmsv8FC8DUAqswwLiaQaOPgKXtkII6Nr8WRR/af2IXGXRPTaNgoS
PWdH/CgYoxvKQVBkaXQjELKQOF2KGXq3/e235veAshgyCrCtWzf5z9TSmaLuCBcFSfDH7xrOSv1V
b/jJconWIY0WKUwJv1ztG9s/C5QirJexl5gDx6oLYxNVnwpg/eSc6hQL0b0EdtPOMWSqt27GKPl2
dQ+zyf/v/RNH/VwhlnrDswqUuOBi4W+XrdCvyyPgvTMwO0hQH+tdkzc1zzWvimd4nZkQJ9kqY+wc
aVfx/KdHEBm2qCpaigyvypJD4qlcP3AoYhc9oK/lDMLdJ1OT6LCGbxxpCJNRp30PtvMCIJ7hN08e
ki/QIxl69rx0N9dwB6H5Dt7ZsI+lDFRJlQKPv9qZiqMOfWohbYZvl3cEJpM4zCMEObvZRsYcR2Va
gDyYlCTvkiEU96SKm9WbhrkngoqC5ETqTMMOjLZl9sIAe5SezgzO28t0GZpZFg8rFDipd89Fpq8A
FZGQBwyDWhui7AtPQtkCRUYxev/hShED48zfqEuYyi6Xd2GzcWFAZnqURIyxh+/zIP/XL9t81QGN
FXVnV0we3RxbY0LXQErmxUMSFHDT+g0wtRWa1Rg6io4f2rF7Or7fqdbA/BG95YrhsPebDbxbZPir
FI9wXUEuls4oBsnoi0F4QpYFyD51RyYvWybP9+2FwqA3Pq7UIqKVx+ENhjg7K4iz1JcWW8Gq+nrH
Y/ZEetuoHcVoqmP2xgdmv1093kaRYwwIDkamfiQAKhCQyHhiGtN97YWhUiGSpT3P+18gdM/OY4vi
5u6mJOT98gqgcRDaU3B/MElaiLzAl6mu0IAtyUgh9hyWcJ8s2NFYNryxM/Fp2AJsbkehX64aOjfr
zU5KqZ207GQKC0ijf+lCSDnfaHelMgOHcqu3fdSNPwV3mn/kNSR2Ytfdexa6Ge1zVZMrzWiYnagV
MNftBcQFq4Y+DFfexQ2oDcPsf/XLXOCfaXaJjVJTe5B9cHUQvmGalmpzwUCPWpIeyaXpHni39Ccu
zu2tr3ROsBHZWJPLOmg1ZFcD6zOyasExjiX/c+ZAGOJlrK8m/2hdzM2op26MDZ+952V7mKxCyotP
juw/xChHjtZo1XRV99sU/cgdOuvspjeMeu0/cICPYGBS+KVFQ5uCUyzIteokjpSDb8PKeHKG56qQ
DVj5jyc4DeVuqBklvzh0Ek18CbmhkeIJ9e51x4wgDiM7ttuX5912O+vrQW6NArmSFcY1lJn+DhZT
Ihi/px3FPawZvkMjQ44mWeFf0Vu0X9eiJrfgpbc5+VT5c4dFjYAJm2c41KJccDKW4rsKMsmFiH0/
Owpi/jsID9vgXWszmvlwDv+U5Q1DNPl+VDyOqKUWdfyY49rEnypPew9Hx5Z2Al8TFjVz9T5wfWNi
MrgljVnZo6/PwxwS8l/YIFgxdoqsIdjOZFjHfWd2rLD/VL2lsqzZrSu1EIikrvJmU/lcVjn9p989
7Xyq/1xgw2qMZ/S53yLcRJ5fTRrtWFmhBXY/VJIGEfyN7BIEP6/Lf3g5vFICxGFJRAy1yE4C4QL9
17za6CKzzdDtrEUAgBwJjQguXzFsKmpWgHRMCSoSL5lU9MKseh9EfNLf7lAqK6JCZtRF0dncfoTp
U3tTcQwJlbQGFI9D8XS5Nor2x2jKN6NsWtCuX+YPEnsZFqdfYV9jSg/eD3VAaYDukclGOjvmMvxZ
7HKwMEVEou4Zl2uCv3BVs7inG56b00st7SKkgonkVlsgwCUhR8VYECEc2yoI2aKowYiMRYFaFMkJ
bID1tTlEygo09NgMGVkh7KPeowVCIPGwR+ADx/HIad4mbiX/53YNKAcFryqLWkS2sFVhKt8DQfNH
1/90NvS4uJOxXsnIU8MP3G258kkOExh0J0HXd8CgQiMMMKHCN/hzDFwTySgNdSLs0CtKwAUiwfUT
LFqHjfScsG1x+sCWpWaA865M5gYDlTWvZHPTBULTz1hPOZ9h1ihqcrbyJBN0qJmm5DAyWReeYww+
5bd7cHHHFAgmdNOtwsPHoqLQ9HWn+7EpdX22EXDAb1LH34W549huDgLXx6oOOLpP1cefaa0kGBWA
GJt91mdXDJdR0ZYbcQkto3YYABx2zOLMp6vMWc9I+hgffPMO1FJykozQ164GM0KyqClj3NribAlN
0KFF6ykIp1yggbEFl09Pq4d5zEj49WDWnAUoEBwF1ywzlx7bQ09acxg+HE0Qn4+3e1fICvW2bJmZ
nMf3JfYHrDWUpn6eAenOdN9T9R6G+dxPlOnBUDSiF8Fd4/2dLRuBvlla3sFG5giLY0DR4VOpZBYr
5hBOuJEXO/QCxooGCTU5n60tkaD7JwlVEMr0fbB36MTRqDodzHIzPmiZ0zlkZtq4XS9TTtwGz3xe
wjbzxBWwfLUXcJtiAMBuHUc2qQsj0XvmuKTwS/Oi2WjY9WgKgLdpChUl1y/aQqoYLHpMub8gVREd
2iIn3+KRWZb2OW4rnBQoru7JCL2qBvfSMzrYbMfPJCB4an20v7KCXs9GaK4zgSsoyn6WTBmzgI/Y
aLARAk5o5EcNuBXMPFzzEqDHTjAkCXKUiN1NPcNXduWUwnel/Sw5QonFomIssfbyV1W3uAblMFaW
AkECLbjOUEIaGt6aQzBuJe1H09wdvOwv1YbnmQCvZVpCD2vGyJwgFTJ+dfON8AbKLwirw7BVF4l/
CQQxltwEaxRDI5o1XqE8J6QN8inbg0Ag/r37rWmBs06urHWETK/xQTgePrYruqvlL9Tj4Iv6N06E
k1dnLO55G7z4kmnQG55+s6g9Njhnf2B/FIZD58TupBK1IY9IaQhQcCthZEt4PEzo9DkEHbHsCH1/
/4jfuelErWv11E9fwkNA1Y+kMEOUr+FbfL9KzsGtLoi6/7nYqIytB8MCvFvq4h/3zUi9VxZbdKWZ
CEX5KtYN1khPVaqWmQ6jSh6A5CA/dKqrqpupSDmm+Ic65EMyzxjx7YkPyRzPYsr4CqWJweA0R+ru
QrW0BzOO5/RTmIAk+d8T9jUzpkO8w3Mq+NhWM/L1AQZA+7m5lAj+yMHlPRfdNx/9t0nbiQt/JSrQ
/pN4ni81YqfgmIpnNysQ4yryw20GzAR35gpg6+ytL9zhV2mOkIJA8fZ8054ylL4IwkW/JC8tljSJ
VIppHwEA933XD1VH7VBi3ujc5/EHVqszt4h9U8SIIUplxMBEFAq7M5D3VQ6cjn7TSMpY5WWHd4oP
pesR9G6EL0G4UepH3kn0WH6Zrd0a6ahW+YKH09VPkb3akxn4q8YKEk/sRxvs0QYNg9SV5es9QnKN
99hbKbJakCCTE0HKcSHX6R39aj0beGwJJly4kTuE1Jfpm0ZgJ+ZuLLGd8cA4NVBfXzbq1fsvQ/Yb
3JJ59mo0dDgZmhvyvK5/gRV4kYKQDCBQWgCkVVtcaWLV4IRNiWIShjM6bZHZP0Iwf6fnIlYyfgvm
ViWSGWs+LcwacvY+fcp25PoeQ1lVo7EThxbjTql0OBS/K5u/YLmZzEIyOF77/Ov6YeRwkTD5mQeZ
FKs+CsaVGxW87cS+TBGmGLTNYwgpUOWnPES3romUAcFeCkuFGKD3uLR9uuiReFEFdcIXP4NlLtTz
jo2R155QWiQz3D4bjiW5ZCey83CFjrUXxkebh4Y4QXYy2FShZ47/FffrI+hWx2CrrUT+Sw162A4y
PT+M1PRbchQ7qY9VWcooJnAIpk1XogxcKkPwdqrUGpAXuuRMHp6QXj6ryQaHa98RCRA7nsT17WCt
RhL/8HYTSnX+wFue+Rg6XOj2PkhUEFCpCe8sbMQ7BrUZ0Ztu6tKZfnjgOuVI/3aDwX0ouo8AXb7W
hXtBLFnQidWaqYUsq7pZVL/kov+nv4ZrNBJg5gdpd9xd13FWoWZG32oMt8TV4vksArK1EG/b6tmv
TpBw/opcYKTASRnLLadq3RExgAVyrJYYxSCjzjszD72TuXV8hjoo3I5echIK0hdJqdWW7AdGjf2S
FLre/10QIw034v1PmW3i6Y1XWXtB/qLj+XdEsBNmN3YvblKtU2GbFMn+hNdBMCLUlKguN+QVlfdV
DNLPmwFweNcyz+e1c1odefGCNmJ7Q/6+b2OnZbKLfbl8Wts1Betlw4lYppb/yIDvChvOk/ZmncG4
1K9Kc3VdMsU4p+nlF5kIEjO6GviF3eHVY1UJ1fedSYlAcERHSIJHZjdvW0uu/9q7Oh0xhIQ3nUZj
/BrB2N0EkHRm4whxDdXy/bcsWU5AmnYrOjzKBDULTZRxwGLIMm96n362SoES1f1Z6c426+EIwe5y
uZT2QnObYv3jWfsfZoC2oC9yeXIv/Al3zUjHNxfrb3o4U7OxdU7by53caSMaMuaFP6tFKEHpDMPP
IbolbgpNNJZLOmPfN+e734X+Fv1u4MgMyuSSTCSb0NWvrPEUFstcvs4VvUUAx1ANwW4tFhMDYN7m
bAtPM1y1GlrOhR1TemFi7Zdb5HjKraItkexhS3hR+lMFeNDSGA6ViCiWyHh2RA7JTVtUIEF7m23S
D6Kw+RiiW4u9wAM6k1eCwNm1k1ou3Yc7ngnDjNhQAhjwHAePYsgeUHKgoWZA46nDpFabvAjzBO7n
Lxyd5FSSxY/YVaCYooPqF25qQF/QfWVaRl0XyzVxkoiNtbCTpP4EMrtAOtbdw//noJikNag7bQfJ
Jc7ZrNJP154vIolRSWH4vHaqQLpFy8Vz8VvqGb0JoeX1EyK5C5+qgEU3vbubBL2VTJwmBYwiwfxb
W5coG6NLF2cVmZs8HVopyV6MxwZUoQwmRGZKE1PgU6ktq4kHHcNzN9xhn+aj5Dzj8gGhuCTJXg/1
of7VUozGRZgzqGHGVxGP6CtEBspD6gWfrImmkUqgdCBRh1d1daX2oid3rkLNkD74Nsx/Yak0j1BP
bNNMpKjrkcUfvCXqlyQ+0r1ti76cAF9zXTUEmiZWbye0DBjfocYME40g8Zw4NBRTLquQxZSJjxLo
mRki1++AxBJblV+zdYgJFewArbLRx6oWMpuMDmsBBVqJeK5TdhIpjTRfVwCdn4k/HwNQgZRt7hTj
7XZt0GvcbvrO1AeLN5bG1NSPMW/E5up8KBb35/Ey5qjaSGdkUek9y7qD3qQ9GvijZKN1qR0x4Orp
IEDX39moroYTezNTq4S+CZgAxgc8i54iYdj3LMbPUL0KHeIUVBJZM7UZg9wJ8/SWrJaY+gtW6+tU
8gW5yavxrDj5rxMidsGrLyp+EF/ybvYWMHvBWwD5Q5BIDx1u1gn192ngWQ+eRGaSs3cjMxiyeg+S
4A14pyJH4SWiwzrHkC/NPYkuXUCH6MoOrJg6YXuMdjoyRAccOPKZ0V+SvEhVzbDgMWRZn5/nTm9B
2CWpFJ3s9LWC6g/NrJPX8mldjgdSO28Mz7D4bJbBVOjta7IACgTMBltMUD+gMJryDUioa7OFUmV1
2gSHLzXYVVWhp1H+wVfh+JbGQaUeFxA05+DLCCkVQ+tONNHycnryx3brVn3ryU3SrnEdZy/ENGsl
RVXIR2auaVjwPL4YSShQSAb3G4YbQZ2DjCnnDC6XgGBy7TtqMDm0AlRJyDy8hCNRAp/HSW0U0i9k
pLY09QSHrrdHMPa+HzzFSfm96u2NSM+zNNjd7ZpN3O7Omoz2BRpS0Qggr59DFxKeQtn1Znit+xvU
Jg7nGZYiTkU3f5cvWYixnrospJrN4wADiO+BJRRFv21vLqEIG4X344mFn437z9icuV9YHpSfYFV8
ktXXdGoqYfEdJFSij9gFLMkO3hoYOre86L2BwQHyZefKK+DIcg797oCQvEm2jhm7Xpd3mA11pYXS
21/HdCaCjRRPrJqhM02vUjbp4n9xr+kulM7qv1GMbT9OBvuknnYs+leiJ8QsPlVogyy/m5FIwVs/
H3vL95xYOAO1CZ+l2WE8RuHDXhZ1epZt/wSSlDg22PgXVpjTDqHPcVynIo+m0fcUKFEFvqMu+Sx0
a1N5HTjdQ9mlL5v60kgeq0kk/7fVeuYs2p7fw06/qEZWOSMlDm4DOKsXQ2jC9tCCVL7SBrphsoVQ
piHM8MAVyxmrvY1CseVQS+phxxoITuUUx/+parnUycht212K79WMVOIspl8g97WK++ZWCXL8k0hh
vewKYuMObyS7Unf/YVxTj7CDLCZwl3hfFRrh8IdOI6/rxjCv0VKVn1ort/0TALbzmBhhM0FJMj4s
DWFIVakyPJUBGwnGPpQpVN8FUjhYW8qJ9YUjWoLN/t6ho3etRTXFTgOPFSEd6HoabPuVyn9AhIBG
JDqmdxN1f57XLa9TasgAw4eKNRTRbcnh+/ag45ScJgRdti/g1AtwUJpJhRNbga9EIsMN3KvivnFL
PKNx4Q9UHZtyy6yC1ctE4uyqA9Ymh8Kg56LhaTT1lL9r+RxcChCxCKCh/5A9cJ532nmOa9NGJocr
Rj9zGzxHhIF/5CLXOcwe5Xaw8HrEq37g9+ntTF8AHzNX2nU5WUrBTgd9qcbM58ca+C0TBowTB4TL
6Co5lgNQ++xP0fwxmkXKFTkcWw41/nPWtqlCmGitknoTdDzY/YnhmF48IIB09KUqzr0PzjE48KXu
KkROMECFEN0d9iVm86cCLRg7LLlU1WJWtyAMg/UcUCOlkl4UOHxo2V/9G9GP7BYWbyCPqCvp286n
rXCaiC9C4ibspewr+ug1HHzZqoZ1axOHGQqo8eb3V5cZZmGsiJlEtaW6BE07c7iy1FrvGiseVezx
QX9u/joJBxn0h6aPWuPCo1Fz+b3nHqJK8QJHmyJkAFuRqXapL2sPP3lx2kkayAWPFm5JrlDGKIzs
DRlKTvXwwqSJ73In0HcMPHlJlB9uzA3oPgrDe6Xn03oqfxWELdbm3sUsZhLZCIPY/XopwJGsfrQ5
SO5OVXtJzRKmVLg+dFuefn51T5MObPcsnQ1hnfooPOXeiCDsnYhL+HAKKhTlNCRnDJYQm7sM4Eql
Of/UvbbeE82xLwRC3L7p1xJ0EWZVK/BLsZmX9SWxGvrMJtT7UpERsYPnpgQdUbVoguGCfV2JLJ0e
KZZOqnGvO9ijzFtRjc6jayTAGtk5cpv6g3o/scutq3zOY3SJ2WccggxaDoCLoAE7DfZf2jPt9Gt/
HMhzXJTO6YCGRlUw5DcdQLWSX/d+gBiYEyAu+xdEFusBXcmIisNcpRlSre7Fp5l0KkaK/fKAKElL
VEkqxgG209LAMPp21GR4j9vf/ToyPHTAVZpZIgpE5apDz/IO1audCfZkSaTOcgGnnh9xoR1yqQOk
P8BdN+br3BDBVUNls6iPG9Eq8bnuJ9M3VlQmN5cvJ/vXrpEVqWEY8iOo9wisaGUdpN/umdCp+huM
LPwKioqBseJHGKzDPb/fKWJJi9NfLAbraaxTNm3EFcOeoXRHk64l+fUct/dNTTDzT22bMTY6x3KG
5YK320NXRJsL2sl/DtfYuIjbW9okSUVFTtSFV1LJE8QWH7FWD7Vznh12V44aM00JBLvn4dJfgKOY
4yoLLbMFjEMf54qxaHsqWzP8PbjBMMs8H3/d1mOA3LpW4ktRk1cHcup5ZhRmDVPO/wUHXkg+o0fy
ZEQ8VLam3nN58+EbOpEizJDYjCcSS+YSXYOq/d6B/8Fq4zTIKo5GBmYX6E+o4QE4elHhHkpX/Kgt
N7gNHrqW/igjFyudgcziZN+S0LKp4aogpLg8zpi3+xGJilvidBUQ0t/Dsdv6D0UKKhoQ84lxNxpQ
EnKqnCmj6w55MSD+L+1jZW7C0AZ9Y6t3L5q1Pw48Dfxt9mOcWlVjPmw9RLl4wf95pbxJRv5T6rUu
wrqva5PDQNprmcg8Egu6jSPOZmXl3FzCZ2e2veVbDa/LrftJs8rZQQhMfvy/GIUjfxLJLzW/HRuD
NyOtDUjAQqT3RGiwxpW1/DHxOfisL83rqWRIbqbbGDvisaHBBY8JAHHmYU5FNowQlRHBiXNtn0vp
KeSp8RtDHeeDyCLWI1r7wW2Oy0U8ZyAT9b/7D9WccENYRG2J/v3sBfWdDNrpTPOFHim0fiLFQU7M
aWvVbwPparC1C2q/NuT0UIcus2mPyp3yPSdAJBv+Hrc32XANXtQeVFu9UVxsSyAC4qRrzccKkpJd
xdIGupd6CNjxxUGRWU5vnu4r0DYjjIIcrSn6hCkLVtIknt3ccxOwrZSTDyhqzuCluRkDdoEtGt7m
qHNF7LOyuug3YIwmQRwYLT7DScEaeaRT9JKw4Megal5TeFQdWiwUsU5WuSOF8qNqso2X3PD8c4sV
qKbYm5DIIr0qz6EiQnnFGklazqpDkEeag2svY6kvbxnGfYUiA4t3Pe670ekR9SMe2MPzjIzCLGO/
cFsCO0vuYR96UXvWeB4KbKGfZ6h0+V7XuZTA9dn7hTGk/suyF3UTnLfk5g1d59CwNZRIajYHBJoW
R8CdG1KS1mRlyAAteHjn56Ik///MaaBbTXZMHnSXo948Hjn7zIv8O2zK/uJE4GA5ziWU9BZjxBIA
l7VqvMJqp6Orbup2Hfq5/oYqLA2cW4+vFPvMJkYJOBEj88+dI7tBH3QUJbSuwcptAiYKOFUaZhTo
0J/Lm/+9pnP0x5mc7fmK4bDmQLdEUy5aIbFJGvS1545WAV7GAkSVhxeaEQax8yuDgXsk62og7nNS
59HF9QwdmPSItRPo9qqEZuGnEOdLan8FTlf2jLWPi4Ibr43n90PMT9T6rb9SzznSS86R19x4RnTf
PbxhIG+Tkbg/+Waj5gecIDAOO0cMS0B7/aQGwK8ZGF0SO5GCJRnzxO+RS8B8BhTlwCNh+CdiLKE0
i3f0zcaFTPSvEczO2WivEZpl6/fuc7OAiK6gsf0mDbWrWsWvUwZfIozklTfGiOYBBrsbMzJAhZFy
4NnfODQHPQnrjfmhb6CICh+Q2CCnXQhmo4Jh/fRsEN/WqAkPBzSsbaMVAJKKUvjCS0mObMenn2WR
JCzGauOjGEdE+J47cWW0a89XVcG0UbXc+Xm1XWMw67fOVbF20le2dj0fdJ/ED+oua21tzNeNw4ox
MiNxNUlWepUbOfdbmRtVM4H7IKaJKrAWQELKAy0o99Lmpot6b8dSCD9kwVqokmXuVTFXxg6708Qo
6UezRnc8XYdaF6DVsANH+8H1NcTQnHLUh1YlrP1nl+44fpH3nZkZbZte/Y807vqlssubpKB+PoG6
/J5XzeIm3tfseWocAUT/0yuKB/UVyLsi8Efj6PWwenMvvJfp2TYUbT9pdUm7VUhbDkbB7ILAUvn1
gZTdoXAJVPifiriiyKiaN03pyCpKOXKiXfhytJNVUsDySKKMN6rqqzQKRJtn+dqhlrlWfL/DAjh6
AAgPHhXzwm6M1WqFAkLPEsmGMGdBgmkl9vpLADPIceuLLKh2qRESlT49oY7w/GaO1vDqP49vg5nH
wLN0RM4Z7+L9VzRpxir1MaXOCTZdttYEPjdL3l9pBe6drNCFnE92bsKLI5wOcn+LyTcQpHIb4pB2
javiPaZGl4wdTWZhPlhWVOYqGGjyP8CRb7PbltZXHmYpmscdiM8vfXVxHPS0JRuKZv8/uoTMpton
kMZmDuFtqH+bfUw0X8ND/XDgGS8BwsR/040n7ZsvzHtxQfePigppZZ5ye8e8F6Z3WyK4T7ZEWIK5
pB2KfUPPMadG9Vwu4kqYWobioPdz/MaMngl0C5i3Robm+VNGm2PzutjpUkAB/5SKnNVeh3Vq+ft8
6ytWyLGxRi5WrsjCTRjWZG+ZCnVT/8Ko/j5Q21gAcQev+0PlDRQCRikO1bRnEawW+rIDdJTP26iE
mnn1znpk76oXcPqTw056n7ESb8iLtQ82+PY7520YlzqzHmgpSU1RSqOsVE636Ixagot+NbjPzIrv
P3GxfAK31lVJqb/XFbuG0OaD35wLs+33OWjNYg53CLFM4Tt2NmOoQpAUkRl/4v6BHrT39aHqJlv3
lN9ZEcu3dODGW70I2xWIRgCPY50rhgbNhlIOQm35CLHJpNBR8cH604qapN7qRctDHh4U1yO2VnlV
PikZuQ4rtKICgAnWFOFwtihFMaaUKmdwef/4aXKA9B91MCJWj+i24JoO4mK3LQjEo1k45JuXqT35
2tyBMkVSFivC1LxNqWDy7ZpkBS0s4h0Rub0Povd22pOXAVNFT0U9zlEWUUbRRvrtPxjaa42JY9f7
1TkNbNJL6SSUBHgSZtR7mGucRhRL+pOcEC/i2l/nN+AQJhv8g7p+dmErRtTWvaSXosFo+1u3m+Q2
W0HirpqSV4VCdTMiHAwsSO3pkFEqD8rijhB6iNXXED/31tuREEFcVWLlzeovXPSpjWEkoBzelND3
/653tmuZjhX+qVvrbyMICKxQY6OfL8BxCX9pA7UcwdUJLO2whk5ccrmsTbWfOlNmvmk7KQQXP1LK
SR2VLCkF13V/XlvvLppOHkd0f9rCf9CGHb/UtXknSn5GiICilVsOneKkr7z5+412ydigBWKy2n+k
lu/JcwPL6jmQewINTTEkH9PznHxj3RW2H22OvG3J3tLI1Ij5ExB8B++O6ydmOOUie87Bhf/1ov2x
4CRs1Nm0VVmcaEJlLHDE3F0FReaW1ggNvP3miF/k0kl1y34XXCDtVpaDoiWyadqtwCz0NdEQi0cZ
L6OnshOcGqG3z7yjhxlBPwLfsA8CWSqXMxF6s0Vd7uba4IbQ9IZjn5pwzxN9cDC4ydhpyCn43rYM
yUz5XKPUCrvsUWou7UzPVIEJ4eq+FZcuYlXcNbi2prnRGxIM1+5ldGX71JQaTLa0HSBMQBqHCQjV
JUrqF2FPRi2LQyE47Z7gu5TDpEKWKJR6x9gZYG8nllo5lbXinzauKQzZ5/YO6I1IkeJsqoCm3Dxd
bt9uafTL3jbpdqm4Qeq1CHM0yNa25cl6EXrZLKGylXlnJmZsNwQJGB1TG6XMJPmxOVZ6GckpS4Px
RASZ8XiXrKP0Xym7nInSrFuTuiShWb9T/s0FoSNE3AnPLJ+cL601a3nFK42o5bK0rSRc4hJ3VLbl
RxibRyu4bvEuVxP1XCszrMHKdKSIC7tT9ZG+mZ/2KAqVGkle9LDopDiOLaDSS1JAq/u7BnZkQsbl
Es9+BlPauBZZpPPfS91JPDaXRb+Y+JfRH6C19zR8dOKRQBuukEaEAlfAbq2mpIYtC4YcFC7vJalI
NM/5ePYD4H5i2ptIQMAZFzT1a0I1FGGzLmjqzXBibEC0i367x1SYEwuFZpUfUH5hKd1FX6hEgwLl
2wju9hG2CPabyHTChO78bIdVf8+xgZChvQDlmQn1AL4jDI8GuvclPfpqsU3C/XC8piRiYS9KDbyl
uadsF2p0rN8oJEhfjYx/XaNI2/G0XlJBm6JGJ0ALjUt+H4c9jTe4ke6KyS3ix3PCG9aVZSHhBg2u
XtuLanR6J4+sKOP/Spt1yDcUpEEn8hZ6lC43T/Viaoe/hcBW5CqY7JZlJN9GU7PH6tuVJdaBBin0
Q58ZiWtNhBA58dmIQ2MOQrIXOdZjxWtZk91fdQvcw/zUF+ZVbcjU9tNoWd/l144kxg02cH3i4wnm
lReEC/nhOKej9hNyxnmPlpq6gxmAXyUN2VUcUS76Fe8NDfUGQl+z4hyE/m5s4nNixErfloz3RjU0
QUesDPNtwDYFOKZMnOqfmqID+k+ACMM/1/nrTNSQ9KPTxLw4LYM5ln3JMW0/MVN9BmGJ6QpO/TjX
0nPZYLwnmrI9owQxU0oj+YeeAi5bfjvWxOPZlHHTepFcYqJN5muvGlGkMw+N2RWBlsRrlGncrVhG
j2p4B15zFph7p2si7bFsj7KUydEzyNfAFOOj5ZTlKEvMJZpRHW5DxKt8j8OW/P/S6NV9Nkth62Sd
kVE1OXtXqbFy0eRZ7zChHwELOzXi3yNwFOypk3FTSExTk3oechunmEWN/x/I3O/O5jhaOtqHJ6Rt
NM5DEgJlCyo7HiOucAdTFjVR+Db60ESs3VwnT801fdQQZV1nx57GuxEBhCyvUEBeCuriT7egOoL9
VYUevFxyrixmJ877zUgWTKGfCYJsaY4NhCXPBkSa++lXwrIgBtDyKWXGLcSxnOmgU/KkaUnKpw8x
w92dQfZcISDEj+R9gVFr5M5Q2g9ZgLfjT1r11/IUgofpzjF7KoLIDlmOxPILYnZh/7EuUJpKpoIK
L2H0UZhhHz4HYrfgSBuVTNH4NJuGiYq8J6etVpJooJGu6fpqSYOwuNbZ8A/i7ZiVgEw9lrwlFBRo
ZDl2nX4Cd3YxKxg9rFe+y434tW95htsVAixAHFuAYFI336EU/BqLAQ4APvngm4JjgRlCZTIvB/zz
GJj9ekiOGjUtC+MKs5JHuNo5bDOizitb8oBrxQhOWC50btD6k9dZ4hLvKXcqb7HsAZq08rC1D4uc
nraGN4taK4wGoB1aLGlx02lYK0tNEHJfuVvr2+nJa0yB8v9SG3NFw4ckJDgc/T4639UlIKSb0yoZ
bOlAT4uHj1kGag5R4L1pi35K57ZJv2hS5Q65axYWGS0cssWQQgIwmNihwxeRevWVGWfQS9HJQZU5
kV+IYBSEsOdjbSwiRQq2M1/3PGFeiXEGAzDtA8wnmz4OvVL/+BiJt8uflWPTl8EvzMzChnZglIKg
GFDzYsGWATHVvHz2nVaiEfbWfbHaQljVcQ/Mg0qk42lmso/OOmakZSRSFqSU/jOREYjC5cMnbbq3
nnGpvE53NAoxr3/uctDhS0iUoQ5WyfApXb1ofLDvLvmwQvYJIThg34GI50ve7AwL4towIQ74LM35
+EBADLya/FE5Hqxb9tpM400KeuZhm7yM988jII1OBNTKxJq1jovNLh18vOPNFIuOx/g1V2sY07fl
0s7xgW/J4Zd16UlRZ2FaAy3QHZowwpxJ7A7Y3lrWMiYlEiG/6HzACBuqztd99afzVHYhv3jlEmtS
He1DXLO7qmPeQN5dxXybHA4+RufQpghIIMqWxszibsPOgTXRyDJbjJh9O9oNt1MtorwTYgaq+f2S
p+pv/uGt1hDB/b2aR7IGiEpq5DQxbB8/4gI6CbDCcPFhCeGG2yHw0awb9wTCe3vYC7iWev3GAR34
gsTxKxtE2vDQz09+H/RoW/q2DV4tCuWRZJyOkaUIUsNcJ/Dn8uDlWyDnvBpIYzdyE3cMRvMSMNEC
aIYOtav/sH2Fnswy/705qF/4XV/PWMv5FOFxLKpwfuS1QUoYk4e3YrfsCfpauFfZFtdPyf6TNMfb
EJLKyEc3MxPl73hq7Vb/1HmVSDyViS/a5yjSCYZ5nTOJmf19P8BGizMZqywhYAwz90msWLpKDiHQ
R7vO6eaQ4L6A2DH89wy2MlZgJj4CR55e8cddhW6fUHsG54Cu5BXM3cUc4PmN+LuIN6EizW28Q0MB
P4FvwHIAbKYJw685GdmxAaES51AKNZFqABeLmBwTWKyR1LtnprLAxf+/YvWYhfMI73hXIDi4LWFz
4Sxi1oKFe93R53O9ViBsxdATNmj/wgdJr/1EH9izcEFrIy42WadYSTmcJGZ10rwJTT0Dle4ceWII
z7jigL0BHygLC798yKsEc0f9wejVjO/eEy86lB/ANgsTlSp8mb1A/MghIbfJflUPdoXlUETuSxb2
7NVq7hOLQWEqUxtSA1CRiRrQtRNE5466eesFDO13uJC2JerQAQ7g+O7+REUwoLZZWZ23Glq40mme
MkxeMQGpolAXUJMpgbFoa4GLr24ijMTyeHVUJngqErscxqTutXrOSrsI3/AJEa4wnlV7QbiUkNmu
0KoCcj8skf36iNlPfeZf3weDvPYsWat0rC+Gc/AiAGXAjsFdNL9ZM/BzS9/G5ZZdUKIoPCbjjW+Z
mpoc7dpODYu7XmXjCtkA6O+Gq5cYgHuwpXTZG6qVCtCECVBMZpEQDWGNYRFMtoP1S+BMHnEGD9x7
3pS+s7eteKrbfPPnS5gaLI9Bm1BNdK9v4gzkRNx/lSnugPOmJZKqf/f0g60XsybXYT3O+i5ADLgT
dxf3BEFaOz5HLXso0ATfFwWpWT9bNwwKR9O1kVElWqErA6790+j5dA07DAOwQH6KTrHg9nVo64iK
sDoO3rtlDqYHp03jQMcxNeTsa0bgk9g/XizpOohXvz0EdMv5N73J+NI6vm1OhTVShkp5Z95aHzVC
1pDHd693/3HyWebtO3MJohbmNbreU0FDuIXZIzrBhGMQZkiTnXMe+IZh3QXQ9N+79KFd7pyrq9cn
piGqSpgtOeQMM6M8lIqsIMRDjaJT06foNSoGUVUtT5FflQ0d1nsZ/0LuWnEUe6wVe8WgaNuhTncy
ik5PQjmslbn+t+NFzALwAlnIMarjNdxNt75fwPQuC+mEGGbS5MXrq0Pj0yY93l1+9iKR5Qnh7Xtb
wlxSeREpSNC+I21chXCbM7TnflgMgQuGmkkOy1VvoIOX9s+Oo6SU4bi/9YW/z942h+IYOULFQzQB
tLU0k8cqUk+MaP2aMyGke/nkFy+p6k/KkgQVsiA1P+a6ajoyuYA2ORf1/Sdm40LeqDxYEVLWI6sl
1ATnZotsK3KHEMgXg8WkSXNyfiqkveEbKhn/wj+2vOq7XTbrGRlUda7dAGqwyGHRvT26vHVLfZN4
Q3lAwmtgWTvmYw0FauTN1cRvJE4QU0cTDrgUmri78oAZMlY4I1NRFzgn9JJW4VlN8ey0uP3NcSu+
xJR03wM/cEp1HmYqsOfD6BxsNrLOZoH65FNMt5khm/woHPstkETTxrGW+rpNrzm7ZDXHgJWtDkdK
+8Y+iF7FUXg6n+0fnK+RjOibNhD6o5iMaRQtI/cdCXC/bJa4y5zW19zvxopLQNVC1XKhExKkuix2
Po3WBKRHcmSOQA0hmVQ5pZgyQ4ftlqhu34H14iff+e3bEgxHFz9aSXlR+HxCtP1EUJ8ikuhgvSsP
+rsiVZ7V19FZNiOzb2j1tlBQShKSQIp/6wZO3ai8tjJu6IPanh0JypPpVURigyjgVpAThMY5czSX
grUBjtoutyCElE5CKgBEYj+3aIiIiG3nHjOjMDXCFUgiobmuIg4s4AOiwrGpR5NgLaRTb+5oBkOG
MyeSNSMaCW+SzN0GdoCAswdnAtVdF+OQnTaSJXdl2MzhauWbaopTmKeXvd674fl+tIlyIVgnybuP
S+RDF/K6ptnl7eHhT51DrGPVcRBedNW8i+uA9Ot2j4OmhwJqlaAH9il+KxDWQQVTiMRtC+XlHx0d
AdkUyv7lcJbz07sf7HaYjvzYboMMt+UAHdih7RT5H3RyQsHXNVPxV66hVIMClNARSpgbY+4apw5s
h73OCJ4PMlcBk1JQ7J2o7AiTkG2qzmFilel0M0T+fYkaqLFPIMAf2L7aGxGb76i7552RavShgo94
Xb2sVXJom34amFlkeo9pKvK8xRr+cqFGIihtTxzGsL3XEpec3UuRgJ1/B7V/LWnZEDI6BuRfjO3r
S7dRSGEIDQxzcfwD0leZA32NimBPf9+SMuYr/6f2u9j2P9pKM7MRD1XYnEmP/uOePEuLXI3lnmR7
tVOpqR0npiu/YUz1MfkhgEx5ttoJwANAM+nkYTYaKHTuJ6qXH2dbYEMncoWCIUnBmxbP4/84xau+
4wkQBD1ybum7ycpeS8Z8++lZgWftnARhTt+fQMSa4Fm1UaJBjbm19xca2LZ7qcYFaEZ5C7D9zqo7
DtCSb16ZdBHXa+77bMU73Lo69InkjJ3mpnUaK5jC+CuvAKkoe1h8ODAFPvdIBreP1tPwSx5wZXD5
lTaYyCsnnQU3ygKKRv+E60gP33+j5uwAzzkK9ditI6CCcB3hi3ezPuuPPzi02SXWX0FLch21sRo0
Pw9oA7jdKkZZG6JpRLIl2RQhym4xl/HIalKlNvBt2KszMCKgOFtGITHZCNlOLr4OXIJbGsXg3pEZ
AysqwdhZ9+KeSAYCQTjHZeHfOSGvWP8VaI1E4yR0lSp8sKMaDBRZUrsB/gmhaUhnlK0J9dRLww9Z
HQCtVmmU0PN5iMNVgIndLiOQSAiyCoF3W2CKUSuwdXexqAPW7yPH4cformd94ARcpLtADzrIchU3
ZlTkilB/nvSe5KPJQ2fsYlYIfNt1pcLOs5n8ZnRrl7qOToKSQ/aPIeqyPk/c3l3+akVxcNClxqEG
fWvWDz59/jw6bOHj0lKXIMwYwsLwzF4yglw484BrMAZ+MCY7tzLi75y6hx6TFHh8s2UbPvjP+Mke
8f0dTAU5eGUcxNiI40aP+JLN313GiDdDz5RP+Or/HSERf9yGDxRLZqMXokL7hlKvt6tgKy3jWpkv
F1oFFQhGiEnVeo4BlJIlRnDZ8maS98oG5OMCfSN5dPPUvf+atBtMTypNHbhOx70PSX5+6mcNzUy8
XdiztOOCb78mvclcEldNifCAHxb3Ii2Pt2NPb/0gljgNfODcmnkU2Nf8aSurI03rtezuQKrzBDf6
rwIZxdp4r6VRXpfx5xJCrfv8YCJTNlFZhYnTOuym9PoBV4+R0P/PHxVZDV3tDz97yO7DiD4aHTS4
9bFluGfHPIOlz+PPJt3JJsHgf9OsHaoGBqJ5/8I/IR7b3CnydSD1TxTJl3PxBpxDLdtAaw5O0YQ/
1a+so7uvlyIQ8RB0jsaVjZfydOTRMLnMIcvKqrm/clXYavYQpSIFXvCXoSW9E1QExdUpt85Tza9i
lxiyILFnGG1WliRJR60nHtL9eskckO6jNwNkLFl45FkIK9Jd9+P6czRcrD2R00L39goAZ7nJlkcM
2CMT6B+u2AEAtP2yf1ZiQRIVVMvYilwWhJxjhKMcnpNG5dhqWN+lOLentH/axzPwOlTxVJ7yZJlf
lJ6aeNLpdif9Bn5+J2KybkauR2OVE8/gYYCqwx8jApijir5hXIva6QL3k9Hdne4+p36cURt1EwsO
xNm3WBFgH4bM9/hBCJzJHgLMFPKSZZohwnMLpeJJeaVP9amuBuwkt4XmF6+I1ly5VKtoIMJrRhdG
F7JVC0yXgcJ1SNXdeN1eJ7yKtNqk9trqXHQ0HfIJisuV28EQpx1fIhiMUDD5XtS2LaX1QQAZ3AWW
5UuZaYYCk8eePBVINsbAuW7xpAT41dtK/w2X7C3e8WTHcvmvnIAMmCW+lxOkoy4CSif1jxbqLSSW
+ChVUgBy/ojq27TESKCDE2P0B52tMiyfePuhwrcV5ei3KcgxMdzRE4Xy2sLvKiW7RKNmzn9pdVxz
urpHRFwx9ZBtwz8e6DohhkgwzRY+BdJvUdptGylW7cZ87w7Vye/20EKr3MmApdVWeyDJ1a8zFnW/
s9IoKXiRM1EnQkTkmV/xw/lru7Z9HeKpUb/mpVrn1mUWJjv/iANf4reQO4c4WrqQOzffPj2J+K9I
fT0LCgK4fA2azGitvsUJ8Ecimd6wT4JLRjhykKE0biisqOS039pujkPec6bTzZtx6Xx3NgKAOX32
ehbF4KSdDmZOIDPrKY8awXEyTsqiUcDd/8SeVLLBiyiclj5Lu84ekECRfoEkZI3HbtnZoXs4kPaO
mrLKe3PebqS8IhbKyoMzA1iYuu1+0Gxi6FPl7Yn632Y9sIFXAHqqGnFd1twSsLl/eAvOihfPHlWt
X73XecQ+QVx/rDp1QZsji8yy2y2eS/Elya+lt5Hu1LJoQLo7K7+hZXSBFxjYm7wTHVd+KJBXRysL
d3f7qJIeBhZp3Yl8XRto7d69YoHSA7dEg879xwU8kYdhXXRHxRaqJeuPZ93ljvifHf2NtTSwYsVb
V9zeAyJV7UAcIKMeWHW4scKGtozJeHRcb9j9R/DH519Eb5rgg+a4gZbHtX+DVH33IL1wyqwOXzxY
94qk+uY7i3uiRoktsMiCQuh8m/cwfa/P8nUItPjkZ6duCsce08+o+ZbSloMWuWgkCJOWoF67dO1R
eMWQgnN4ouBqZo0Uf7a5E4mIUvEMcmHpVIz0/cEYZOg1UXI371SKnrVDgLHcuGs8OnZJy6hr9+hc
ekGNg6Ngvmbv0ZJ/LWlYKkb11Hg4McV2zPWCnLtfFNPh7twp5LIMLP7IX2fSovgx7YtFxVI4H42g
IYqaFePhYncxmJfmaFpYmYHuDf5FmEJDcuP7y36LS8r08xGyC766jK8A1VCtxim+clos/4bhw6sK
txrydbTLdKO+Z/Zu5BerYDVZcZotko7jiic1jsrZYCq2IEWIJ9xO651qlJnh0YAUhu8v4ok3zfnM
RMULepx4RTga9uFJbV+qEjqni5n0OEFU1Q49CEaVrrR5ItAhHO4Ta1R4KNSLMfqOXo2qja06eDWd
Q1pg6t5/jVykGVgn3+PATJeGf9YAI94jXJSqhdULB8iRlv749m8NbOd2tjc0zUppBshUL3pWR/Pt
YFjgX8qhofn9kEFhhRip4LiQB9TcjKr1feKJpDVmzMqPotr6EaPmvBDBPAuGom/dN+5vRNM34xo3
Qd2SD/wQ36GI5KA7P0W7Tj+IRcXBSAvZSF6Fg3ZkV4vnNyGFgE9AYoTqWHnKkVmX+lix7JiyA8x2
oQ6bfN+FgSbw3RLoBYyh8yi7JKAZW+Gcz2viWaTHLlE6NbkkTJh7zGAOoCcSZVHZRlYg5vHzJgYR
GdMoTsih5ggI8RsBlVYNdcE5aAuT0B5u2+WQ6cudp+0lGZakzKt20KZDkckZ/rrYutF5FHsvWNjr
5z99giDci0fb+O2jBAMwSAu8ZvimDbpmvapb9nDpF1hMemLhqrMN99Cz2Scez39kB4zyZyKl2Mqc
Q+pbzMySDrzqrdAJRvIAkCtIP6SFXhpFy77t4JzOF0JiLQrUz4KtxLkFBdCvTNJzuvW+2phH7bEq
Tve0z1BXiDwBv4EJwk06JJAecL6FWWATGvNyt3VM1JmpH08JcM/Wq5g7c1xeC7uRSWqghLcOZiv7
mW3K/euhAXr6D/v64fuBJT44jf8K5Ni3JIdTfKYh/OnZz3GvTNEYKHcqwTqJmNCG/ntSoZPBmfMq
NOZ658CA0UN3t37YkZTOke/MrcICkzwUibk1R9SEwJs5AsnHl+vNK2zRHZIDAYXTtu/8hHNBAswm
7pEL8eRUW67HEWrGLaXtlRucBkxwb/zId/D+byyBG+SNbA3UGICW/a9W4mzR56ptBPr9q8kfhR0N
/YhmlZDZUXKT/S5Ujs5DKiibv3P6otC6RJcYq5QzKyT+oUPMkSG1QTnwIitK+2t7f1Vla87RjLEX
x4g+zJM+rhrJbcZpLaP8TAenZNX6BsEAyxwqBfywLvgG84hpmMRnTY9mgLtIfQh79WtcFdc7ZgZy
zAi/x6gGvR/fSatZUavlZWcKZ1HGCwl+Ledbo7XgCSHQaSI2zIZ1+b+TXe5MzIGFDg4V/v2FKyG3
lANIvsTiX4pPg5PYThynh7hSlUKbZER6teEZxyuAezjfpZ6Q2KPhNrc6EbiaaxsjoU5Z3d1oERGM
HcRoA+6VHtfVRlod0rDTjW9rFCOcI9TmLxzaK3wtaakOK2frO3E0KPELp5SmR6clGWgqLRQDB22L
MwVGH0+cAb1Xl/1fVEc5osZqoIiPWqQUkOdiZcX7nBausmDZ1R4rNrOZpjz1Jz0V9f105iZlcjNY
4QzAui5xfXtfelHVloL3Py7bHhtk6N7+l3D+IOkG8zv7Ui/9gUbpNvAU4JPpYILVFbLGLJlJCXR/
DRLFzWOjTVQlJW6Kn8AUV+6CCSdhxtrrBKF+YvJQGdwnBbauy6Op1gZmkAihwpbuMTuMcluksGZx
5sJhopzNDl5kMpDpoB5IA5ASKvhUQfVaNQkCaB8qXoZ1jeJnGAOq6wcbqQz9etYMIaJGWdb1DNth
TsMI31BtbO/LHuj9bjwH50of5uCvQaNT0E2SFmYy5HRCl3LAqjH4kssaM/Go7CeZ8e1q3S26I2Zs
xr9gysV4hpP7ZaX21bzCFjAIFA1q+RXuXmFveG0YmWP5/aiddwzRcPE5KQIdpxEXV6GxXtP6ZULj
tgAgYadmfpH7XKnqtOl1stG/uSjSr5IXbErlxi/FtF2oCOmQdwpL+4jYSI5vJD3SHbq/nGvoZNig
PCg1aJS96vpN3vi2k70FWYgXCT+OfLGFMjI2a0o678XJvmHSd1ej/vhckc2w2f5j26N2KlppflLg
vd7Ig+atDVIoMT/1zsDCb56lgjL6ATyYuXyl34LSrBCpjJ+f5hwOQ9WvqvB7Zbx5s8C/S1qSeYmk
SzXtOMFdPJVhONI6Jvs51OM+uyNwLyhIUf9JP/BAtClQMMI58VOQ/v5yrKpm+SKW4KZ/Px+FyY+8
gaA2ZdHjkEJxHoxjQ/p0ePeg7vX5DLmqATQhT51LK133xMkblCe64n28norIEs7lcuI19H/9lPxu
fneGCXBaMzvMWSheQgIMnn0lDFTMfBUys/r3XIGYYKx5LvN3rmdPZ73c6yjeE5CiiYXAAeRM22Ku
JNzIRnrZ4aOBlP2IxWnPXYqp79I0ZI0ILV9LH41KljIKU545jZDnGoLxCcf8sy8DyoVAsXs9Hm+3
qYKXZEW6/9ux8e5WMg1R879yKjJzZu921rnADqtADdCTjdDmf9VNNpMca8WkFChNiNy/EqvgFY2i
RuOYJCMqbL659m0JZvTLhGGXRM0brcodgXMvQzl4j7F6zuhNq+aJT0eeTaA5tWJfIPlOKpwhZZHk
sOmL2of+e3ScxGsxXrapW60QdiHIHWS/j4z6vkgUikONSVWyUmkmZpRtXolwO8Qfu+uVRATwaaCz
r55IcLT8w6Okrk3LVCOg07fmWsL0ze9BuYr0BFM0CT3c3xBuDkleynT9IuFTXJ8UGQulZxAtOA0n
83RspRei9Wct4DDi/AI317+dvaIFQDBHoiYxM1d86ZDv9qaGnfQhw8b/w/ag7wU0LXulJz8FvSVJ
RCAYcNCZAUxgtnlAiuHmdK2ZfWGYHH5Vby6med/S9tcRH2bAK+C0b5kHmnRn7sUa75eKSa72qvBr
2ydxcTSLKW4T3ZWpsX2wATqaQ6WioYxw3ME4gdCFtnGtySfIciUkuQd/pU5pk90BICOstChdeTGo
6QrcwIUSm6k0tK3SpRvKNa3QW7cXpXGLQr+MYe8jp+Mu/Zv0+/Ipt+X9qHWp1nGjezxhly6rXSHQ
i2qXj57WNM8C6jwpTTJro5TKb0PgBUWr9SxISLmg84tjnBnRUfVsn2aauTg2idhIUoBXdR0uilvR
YRKQATHrqWeu/e1cBenrTCHvTwMl1PCymuWYmDFdv6SFwcMGOi4nN65iYAQnjvBYo3EMkEG/Rhv0
/nZZt2M3Hz3OTTxONaHZX8T9um/Gcf6Bv39It7/sypJ8D9IhRSolsU8ZACSDH0R979bZWZ1ITRyJ
wGVI/QLucvZ9SYZ/U3uux+d4os8unB3tLpnTKfNCOLV41LiPzKi24RzgJFlUjcbdW7D2Iz+9UoXf
lz91ezGxV+uptKhgq6e3Q+rmQ1MCvayj8G4ytBNe5oGXPPdXi0pRnlSnETRBnGHGPpw4rR1A8vk/
AtPa/fjcTp4BMCE6TTImNlSsK59mEnX7gY897BSc/34x4PkHnPGEFKZy8/L6k+ypgLwAKJTlXx8m
uLLNUQyMDsFHLAVTXr9M7wxykT5uz3kXSWpKybyEDpE77RdZWPtBIXY/imwsr+yAz/qYLFX/pXyl
gLLryfbjfrILb36SuC+5/lvjTMxHP5NBp4WSWv/c3sUUERu88BeUvBfjXhb0oYm16Id2F5k9IJxx
isvrbOhfUzxeLmudfNvjOeElR4wdLyPVfbk0J58ee7ZLFNFC5pfgnijbsdRsH33EEuRdoJSN3KCA
bYN5mV3DWrCcMOWLSTBFbzoP2Q2T3jSlJV1lL9RIT4Gxa/bMtGLL8qNRCRs1NiepyTC/hV4L5ldZ
ycvtfye3gX3GwZA5UDpN8z1prcC8HvtIkDRkqUY2cNme5zP7+c1Sgm01bzBPRl35ejieVjBIBvLy
VoAbofmBMY3sGOnL83N3u/CY1bbM8exf4jixctMtWzT8OIJYpXDNTgNIFNrwK5qb5NGxXSfqiutI
A/56Zqnk4YMIJS6cha+5XtPfL2j0ou0cIqR8M6RhcGNLwcuD3zuyXXn6BjRJcBqnI1/PrVtabOmH
egx9TOnZJbsxpw1Sn2BgWVhUWt9K0Mi4i/9TWFrFY1i812Z1Ve5h728a1SQa6OWyr8Z/69m6yqp7
IN9yY/cACrQ5XfEFRKVIC+ROs/KN01Fv520fpRaJiDjASTl6b694cOboqYPyplpwgnd23l5GWbsW
K++ymZ5mP27D3LQlvX0sK3bHuMNEVzOY2TOBkT/MHcnlkLtAQjnEav2n/qiTZP+XaWwRGnG0kpmA
KzyC6rCYDJNtaGvuHKKeuXt/cFM5CYxo6py4TNXXt1s4EiT/6TXO77HobT4mQTlZb1v2+kKFvU2l
WNvoRj17Pcid+pX6PNDw48VDhYDCoBUSCx8+oYzkY/oOS5oLPLHdT2Y1Z3bldb6Nf12/BR/UL9ih
/BJZhNIxRBw+Cggy1el7SHD/rKCiJvsrx4HXN0ShIc7mBBIGbq0AEvz+lBb8d5ZChwR1DXgiqOPT
Rjn+S5blDRUYJuqDdofPBTg906XaOqh5MZq2R/LvPpIUkvYUliCBjH8YVH1OGLMyEISLpvIYhG3W
jMIajBOMbg2zbt2gFWNmMaZj56sEt9zMIYgd+pdiZ0V8XlmKi4ne8ASVWhZrqXJn0JVcejuhp364
ssmI4ZQ+OotfDlI5NFF44Qb8EYDEBG5s5+V8Rx46/VDH85dmbJ06RySLcE/zzqPZQiB+QGRs/7re
NKAhWW0c8OoyK3KNwZxFbCIWN0VtV+gn06wJiCZ8chdiC7MbJH7R3lf5WNMTQdqeAq8Ob0relOGH
2svJ2HvBiTywtMznjfDZfHriVeQFlRC2x6JSn+sX3x/8V5hBN4WFEJrKccF0Wwy8TuDt3hDFHTfx
FukRMoOi6YOtn0ozoY5wAnfluPJpncgFdrI7K5SGhQtOrljwGPill0C5zyCc6N7Q9TK4dFJI+x+3
0BYInTGP9tRqbY42WvQ45BN81IKyhjsKrIbvxSYzdLW8WW9LocYLa2iwpIiIIKrxpLbm6K7OWYfQ
Fs/86g1VWHTeCf+/P353rcxFOM3uW6HjEEuT2Fl4tCXBN3yCr0QGh6xfbXQ/o3oG8JSKaGaVLPwx
3onWCVRjbI13EXIy5pFDHRHkd9KnkNDDry1fpkVLTe/VmzX3CBig/2CCDsNnS1tzxVNoAitCE7Sx
whHKHajQ3UBw2KqU8Bb+g1wosevevk5KCiEzdBMOqMMzAqP+toAaKlTjszupITuZ3m7qnnf84pS0
XD6qgQF/9zz5mKcZls383MiuVHJsWDzIzYBOneKo+1Tv2SWlUCLb46NN9BV1Ajz6iiXYc1qgFNP9
XVcsFy92zfrBMzWl36dUBemTOLecGScS8HDQcmZeEa1XY+V5sJNHBfuwut7KK643GAuUmhWzcSU1
E5Em68cS5vTG7I2jsPB4GDlZWdrP2kiN5rzeGc4FAaYqERGd1za/lmFkr40M/yyKUoKqsGzoaWg4
ipknsCCyhASHkUmvO1hI4K8QpxqAzigHJ5GPKo0L65mczA70577e9NEo4FKXSVBkPQODo/Kg5AlX
siRgg/4wDSTBSw5Lkn1kfor+mU2JjAajZzz6WiGbIy+L4fn6SaWcFYo/hO91MAABtlkGoSAIlrqt
qevf6L81hxInhH6JaYg7/wJ1z7NI8KpPizZXM3TxDScbVgxBp7P7mXxYESbWpdIZicD/aocrw2zS
EfdhraUcmp2u4uJL2LBJ/Jz+iDkBzJ5lDMVF31AIxXjWxO0RYOnjSQupZFtTCta6T4601a2zeKDX
g9eG6fdo5+0GRbgFJovoaayHtzLeJIJm0qz9MDV3SsKXldidIPrxJ8yERPF/rO6eWU8dN557bWOR
7otPnSL53v92/JCV9u2XLqKWVxAQHGPBwesvv4FhIQox/3sdaSwA5GXARfXNkot2CPxODSBbfxdX
wsX1FRRvuOwyOpxELqBRG5TDxmtXFt6wYCD+6IM2JLBrXjZfqMOxq5lTYnNsDca4uOLn8hdq7enI
KLIyXthaGJ93kNsL6wDbyL7znR65wfRzjyEoCVlG8hq6VLAZJJWpMg+CLj3kL1RwxtHgNg7XktDO
k6F5nxAYSxKZ3k8uOxq+FXWla1az1l+9gUAT3qZT8EttqhptwIGUCX9c7JaRZNl3M2EzZXLFHyB/
a/ISvcwOEY1GeXEB5CKPnbGn7rPhaWITe3N9ETnVclQImpZGWMMsWzO7x8LyTAiDfcuoSAj+toWf
2sCGU5ZRgeBY2V78oAh5V9d8xGmDycangDbxWwELd6q8GSKpgNpXEMQBK0QIfkzBqwggSmn5R4US
CLR3Qrp8+/NLkdSGIaadf07A30ZnsBWU1oHPmqYHXaG5dNQ6F8YWV2xBT8bq41RBF0hAHqXTqcMq
5zu4AQ/j2B0WzEaDyvJtm03KW40mnMnGdUgLeSZGGMJoQ1MoCE6lnZKl5jyILlPa0qCOJSj6+UAR
E4/eWP64uztJ5pi0iYM/dyevm4NaXn6I7EGunP549Lf50tpGmqfhmCQYv2v1oiR2tWNJf1Q5maQy
vKC5wtV66W4NJTrEpqf4q2ljR/0BGwm5+aUE/H99Up/U3ts60931FWvOMEoBAEAjJ4rr0ob4vXZI
B+sZkQBCvIm9J+SmbO9w/FdiRve2HVu+K+K+DUWVPbd1odiqoXDVa75SLJdaFCuDGgM9oay8Jsut
IhDcyaPUguf8z8kwGokmewxsOB3jKxh6nbgKCxXErhozi+JYTizyd5xmBuwI3ICut1kpOzyeJ+Ck
HrZIHJdq8ZvQ5JOr84WRoEVsOFZfbKY2GxYCbSDU2hFufTKC6sX0RuEEhxisF7yaMTtwHddP+LKF
GeVeLeLHMP/CVMBgQo2FNPbfsajkDkv9xqkNU2aKedevzCEWpUr5oc36KjH38qVKbbPPON8KAlVJ
OQPWhiOoHqHrzHPSGNWDHIqVtPs0QRQ9ICOW0dhzxcQYNCRX7RzkxHf6h3MBOKrXW76f4FiA7ZLx
1y5mp7qseJu4o5zKjm+mOa1Z/cBA0N/gFBD9jZDajXT1R3bxhiT1vzvWVndXqlBiGJHQJBUPMVHD
e5NKuH3gvhJ/TJup4TX2F1RAStOLJYrBXCcVTTZ12mnw0pa4srADElIqTN2wWsCoB0yi4S4AcKiz
0Hj/clP1aiwPkPySDTJJKw7LuZ9aAibCuG/OoZqknEBAZdJbKhLBlt6D6DbYPGqwgU9whDiOuCdi
v5sJZW0LmkVikZvBTXUTbIymWyyvP4cEt/CuzOd/3a2pcvyM027E1reHdaG9WSugAqDFSIVnsDvy
A44WIvfIq1Du9tuFNI3wH6vbLQM5pRDrtRqEJfdtyH5YrTV3/VdNK4+wFgXuCwS8QudPI3IL3e18
GDDUBzDmfl6MIxteZu3lSYaxo0IoyGE68Bu3sOlaPbjIJQ0aCqzRQCz5DN+bC9bE52H4GxeZ+8Y/
+ucJTa+CPt6vwRQIb/TunlV9tAo36sWmglhI/bTcPjdpfKdTfL4E+VSauBU0P2GvMYLtf2xCDAct
l/FnBiPxI1yqL8fehwrRx3szP2BzzfitldG9b2+ZWkn/RPRnvu7cH+S5tCNsTzaQc+E/SXgYExII
XoeWmtST0cajSmydeHdW1D6lQohxMwAxwpFTLaf9OVaurfHkZyBliE/7VK+ZUovvg0vnG6gIWJ7s
e/WpraITwSEaTMjMAxb2kIkAqwpayl3mN2O3pDJ80JytP7bT/dGl34oiuXGO8cx0E3MhkNscIEr3
XeTeKG2cVXS+2cZI5hr9lXuu1eZ26rZ6Uz9eIuo27Tt9L9+mlpBwJLswYXQQwb1yXTxjxtDEO9UZ
tbWgSvB5+JK7gPwielKMnM1CTFo0UCF8ltLtWZorC01k0Z7TcArf4rIH5VIiglcvS54kFa6s4AN9
DjB73200drMvk9ZJmVzYwnhGXefbPvwU8mEkJA2BoTDvixEpkiO//1daZGwBzs6ZVtdRn221YgDG
cPhvnhknn2ve6KZs7SPGH6My4A/Hn07KaiDujzru6ZbS9rWRZ0qCd0AvMZqsUZw90SScuATM/iCu
ZWicpbbH86pm0ER4xnhOWYt9edOk8lfmEVxmBx5A7y3rci2pEcKedjGShCPMYyOanxu8VVgDWKyt
14vbgamCNmtOR+NO/ERf/9593ilU8iCfoEywPWEiM+VkFTTTSXjCCRQsoDw8av0puuVPcfZjjhXK
OPCSlb+nwjQ1n4olFsmmblwlMxXTnky5uk8aix4q52+gRK6jQ8y7YfEvA+M82LTk1qpXmk7dcThm
+wO6JWwEt9KYpKJFjxiFMJwL3vthNHPE2sWMSEFq36SF7bNPt7UuqoMXSFjLqgQEcrxpIWMg8Y+m
VYQp6TIYFnS6OhJTTVoIBIZbdtzN6KmFdDmw9zWdJSyk/hGiod5tteaOtfE1MSK/aC9Jl6h3JC7p
3Ny5bevJ6qgeUEl8aIu1oHaAPwjVacPXeZawDZqNgGXM5tOO/J/j5t/iFO7JWdqdkSqYi9fcK+D/
KJ1f+i2Oh/5V8eDe1vdl/3vMbftmpwpAodLnf4LbL3UPLJTqJa2gIK0RQOCoeiCHFLqzinALUVSa
g29MVChtRZbdjNx5vWfZtPiEkkYqXicFxTdPnsk6cl0gH13yoZfrvBENkSewg70/v+QffFF5y1Yh
8LpnTZ1javTXpgJ665+U1TsOL65hnqZsYgGYzc1P7rQu5KScwZhnrbTgQSasE/n/4SEQOu9tQCv5
DNr6Zb6kKc8AX5NCmjORHbt84rM2jK4sVBggr7Vxblv/OgJaQfqDiKphIUYi+uBiMROS0YrnCaBV
tnWyFiz0vIvlOeHCLO5yFyAB8ja6vidpq6DQoE+at2LYbJGCqGHHvdLcvMDOi1aX58kVqxGc5vmO
cQv8nbvuLPwx4taXPL+Y+X9/DtdFU80KOlyQyKGpCvVmrzO0pan8s23o0BWjXbLUIVf8TtbyXB2L
n5DN7iAzOhcwR7M9KMUmQLNsBbSJsRQvS8rSJjQlJ8m1LMHOvvmMVSAbILHqiBrrICsNoZMUkPvM
WF3gpdgrTxjL8GK4FzHstxclQDUAjFut/P2fFt9SGdJtNLjaQYQkfREHxTFbR/Tzcz6zo5vKCisd
Tsb7JKCy9nHK09Fudq+5qfHe2lfYW61Ug/jz/ULAxYYd/imxcm3E5JRB8qmhBcxN5lTSECz4F6Uk
AC3WAVJWPHjO6xrI8RNQhQ+5gxYKZmDOSg88LEqCUOPQome/wpw6CQV/D9P5IiiHytumQoGNtoTD
4u9a7ub0tSUtrK7SvhkBe69kBNfGXbtWkdSjw8b1wy7Le8zpZZXz7kz+/zyOUUNWxBsw7P/ILrYo
8bCbmiCdjNhiwqRCMU4MPED4Xm+inWtvF/8/lHR4Pgc9P/JRaPHI6LMTtbpY4gsKrXVXnBrp3G8u
oV67qBWWqWs2NDNtarU0Qwj/UWguIMy6dqQpEPzLG+fStZSX/Noym/7C9OQIQYUJGPF7Ntjq9+Yh
Nd3mvrhDrm5oSvzeNc0rNf4Nj4DwnFU7jKNozSD+gtfj6Xo6n9UG9m5Z4E0fjSx8IX4zX0lrcHfZ
3hjRUuhiKUN2kG/Wy5AJqXWKDvG9g+qlNWPZIv0BYzWJmalX5GQtjGevmVbwXTtQkSMt5V0FXHhc
RfjsrOkY+bZaBs6VCv+3IQr8GePjWCxbbueNmkGO9IOLqmjdFtCe89EqM/nLjR4NHhx+goYzsXGc
22ViZZVAiEvTzE3TKp5UJRpun78Hyl5ufSDhBy51lkG5qfNvw9HVDcldiuTncHmPylTLiJb88sdb
VbqksPectkctmYsz7TqJ1OLuYHgib+QthrQwr4n16iwKd9Ox//mtfULDz8CId9P3xhqbhahR2D6r
iYmhR6tFm3xpyAo23DOQgc3yWS79SNfiYo0Vd00jtnRgVgEWqxWPH9fbObrCyEXa6kMswLLquPxe
Ml8JtXcG21kBXjQaxtz6DLENQtRkd5J5aBeAdHI1WtLkln4OhbecvLQpCk3Vfc0GBHYVX3PNNghO
VtmzsZxLIuwBObShJnClLJH3sAZU6hPCD5gxlhXraOR/EO8WZ3x1sgTVjaBKrEpohzTvXyWNBv8D
Y4E8dL/IumZTEiJEhp8NUTXN+41xQS+ifbF2e2sSH1d2GAY0XW125yo8olAW+pEWMtSmvB8MrKDU
XOqKPtPtjILwjvfHyKKkbXV+13LA4dogk/lgtV6E313IMqNEZgkt/z15BHl6jebwaGTBhLNKorCU
4Jzquwu/DDhWNd/iZNtfWDAeYlPyhNoGlckLChOUdp0ofvAl2UbR2RcnbylIpcm2ao7yOEbZ5LA+
LCm3nyeMrCLDjKrTorfI0LwfWBfNJwsVXLPydNe09djtH4xwDV82z6JVZPCR0qfziYKnSGW16WlU
wJeVfzoPLADMmdSBBmn1PXWXpCx+NLjNMl1OpdJPnK1ktltLh0IJI6ELnq38/gH3gxfyN5wHK/lo
CBhHegEyyp+AC9cFRtW/iEypu8xOHo530fRNwlhWdSis+dismfKwE5DkC3emtgeOZIC0YL8Uy15e
ESijipFpZwlyyzz2HNtjpvIw9/XIsvMY4clqX1fJ5lqNTMDamHNYrWRUzeTVZTH38nx+IhNBZH76
1HcocJSmRXI6dFOBUyRx8La+jTEc478vh1cjR5N4lryvzXcIU+/PzxpLB1UXyF7linuPz7tAOR35
Oa5QotrWA5MqKrWwAmzApAKYEonmb+9QVjXKEZuZxkTJSYp0eR+ngFlM93zOHnP7ez+NItmSaUw3
DPJ0yAYtOsvN6KXX/AeIAnnfeGINiIeAj17L/9s+cytha/uCMRi2no1UvWGzEV+bUbHW3ROgNhi5
1TC2MYVgneCc2p3fHLUTlu2yT4a8z1M7eu8t1iNGdpcqEiL8ewz7nXkXRKrHztHZL6dO3UCQj19U
XA96Sik1uYgHOpLbX7nhpqfGYUv94MEk2d2i1Xp8e8eOVkNl1K3UENGGoY6IZgJolnuG2N0NWjxN
IlNeXPMeZDXJVIWCnFr/ktzfPedJGAcmU1MhAuK4WDZAz+ecR8k85QQ1rRRKZvINaTC8E0nZXda1
nOrRR/52DBC1alftlGulYm7JAVMSZMAuEREAkVT/sOLlinTbkPOZXObKH8PLEFgt3CNTZ7jYEjHb
ZMYIVLfQwy5B2vM6rzn5UsPMZSb9JyoS/d/twcJnxtOMOlCFp55c94HEX/0FVWM6mj4/3uS7DyXe
qaxUmrtxC5kRg0m9hnr8zYRghcxyG18nVutaFLTLLVtMf26M5WwSZz0MIQB5wOaXL+1UQxSeP4KR
ThYKlpmDzS2cOpB7jwtBLFr4zIjwaSRKsWZiNqHn8ubmLviqpH2A1ohD46QgQ9K/QWO57H75P3Wr
w1QXSxf8n7C9rp4hmPahhmf57FNuieLVDwh/e8SkGTdsKjH4JrL3fUbdYnHPWDoKt7jrIfLeVw+r
Vz8LIw/DkJs/rj59gTGM4ZquPnovlqseDPlH6S0y9onqAAHDRExLCwIr18dqXtnlJs0/o2WdoxRQ
q4GQr1yve9pquGcxR9V/A57t8MLUSMdEgWxCBTzsEGRNNUp/xnPk6H/RsI4NWnW7C97j0YQUY5jf
dJzi605Yqs20H0BUGLciRFzZ7mJJlMz3ujZv/piqU5dY23KfzzEZC115hvn8pv+zuPN4QaGkYxDV
laiiYLhh7jxVBK2ncYga/5tDwfENAg1TFqhf5D18Bijz2xJId3DGf4u+kDOkWUUl5xMHFQZ9ecel
/mHTmkmyG46WnejJbXmrrrC7PRkPt6MoutA/vryt/bknc0FiARN7k6A7yiylcLBD7ievtX7BVfLj
YpypMnc6ohSFItYSvZ3g+P0DFLBRrJ38UsO3dN78kRsaLnkIWz9ufILyaEZg16JLA9Hw3+wHzmIi
+Utha91oRrglxhEztYOGUxdxKz5q+aYOX8SQJ9bQY1Q4DbtqxrP8XiI05Gbss36lnRynglp+0qHY
C16sCHNkDO+kxzqNaHJvoOnl7vE54AtkQhx3DkYUpnEI+2z3XvEXIl8QxkIuvz7HgRCCVXiY8+Rq
bM7s8c76g+07CcBvm7EgCfyybrCGOttcJb8Ixt9CJTw5bGRgm3GwtCo3naXmKMpwiOvWX6W0V0zW
DeNbPLU2xpgYGjSpvbUVCXHS1bxi+GSXt6lSEQ0iVT2Z7aGe8M6i0WeJrMtnEhV29nDsRbfGXs41
gW55wE2o89V+0fI0SI2rtT1hZC7B+WgWizVHmuyPrB4nZP6YAA9LojLLQ4THBNV5v4v7CbR+NXSJ
4PomEQVlcBKMkoVG5hnZW9MDICb1IF+kUczPRc+j39jfaECMzoCBoQM5WatHtEchxuxmceY2TXEi
25cTFlT1rHLzlkJPXh+nC+go8TgQQp5rZb4LH/2hMaxkJ8iDPV43Bknp8bgGWGxowfN2OKA8CyDm
F8y8rZuNJkgfp/2aau9SQzhOMVqZYGvCfUV0FB+nIL2YUYdsMRZZJxEzckArkCJWLCfMgVRQDWKN
3DgJpQISXV8bOjW3qK7twcmZlTIKxizNMH6N0BTXtZAHKtmSqftv/nQdwguCiUHji8E9l3WgmSHQ
K8JjCsEa5+BsGF3yuCcC/qAkpwrZq0DepzuqF82iDTr+pFlgLg6vwvev2Xff/yH1+kzLIIWS7nge
BUn/cq695NkpK2BAUNq6fKM7Pu+pC80UBryc7lHezeeYPpkVoBUNkNInWLom6YWRVvF2crn9S2Fc
8ARIo29tHzi46bArR1fsU2wRx7I4xH4pXzJe2YLNmDOlPKGdllEGkYuic0v6rH7AYnbX97Iu7PSe
TztECb9IZXzs8J+5ttwoy/LvQce8g37mhrHcW/10KR8em8TduZU8xn2xgeMQwTJ/JmquYn9Q8KoP
sjRJUIBNhVpmr1qAFjSEQHnaR92PA87X20gmCDWl/Gbnw6MwszCneSctPWxJZsAaOAXZFBnJEz0y
eyHEa86Qazsy4V9vJrPV86lODEanB8mSmChMM/QOg0GdPZg3+ApvsAwfCBNmnU71r7mPF8rMFYl5
crYesS9N4BlPjY5UecCCNygC+OwNYxFHVna+NjSFM7gibpROQxeK05zGFPQsNv1FdXBOw06Wpwn+
L+ic87J4lP0I/AZ5C9W3MObGM+OHzqc+9v4UMgYTzMFpg5RR0KnF18aFMd+oP6ZDa1lVoUl/tjQP
YOP//mxC8vwe2GFbmTQkHvcpsKCqI+mt/7ncKAXXgLEDQiW4sjnv9r1fxm6hCQ+mKmD7OsWYilkm
U1pAgiuKb03bkj8ke/NUhfuWoyHLkbG7b69iuiSX2W8nduxuB6UXt9yH3HUlbSdMnvlIBu8OqxQL
kZV8thpkw1aa703pchLowgPkGXrmZo1KsVOo7V9HuQQR7YVbDqWj8i7mev004Baf8bH4Hl9mMVEH
NzFvJNOd37zWIwio8Syewfrt91Bk/SaiIQbLjt+ZfL9lf62Y/n1dcwXKuV16TYgWq2HUSGwVRJHD
IHNcgEQJ+A/jGtkaoknrJu3FU5KLfTqjaEtN6T3irIfpS0uFbaMI4I59KMlHdlgfr6ucrByh+iYz
1YshAaYW5XJiDwo7vkjrnn6GfiIy1VGX3XZAazSRmPwGFQrois11RZ6jx+e5CEAijBQGyH2tfjfa
qk3s7fRNltAyP7Tt/YV/dzuX5BL/zqdcKISp8xGSbxl0yIlVp4eJ6LSsVwdU3OL6NSyfSs3JQaxD
Y2LUiwoxKHaNxwJ45qwm8DD9Pe0ngMrArDy6dB9yijhp6lMHSl38nXLfj96JSfGXXvVEzXodsATU
6yhWZXOXArz9mwcrP/Z8lCDQeJEfuPmzbBH25IXDqqmv5DkR9S1gs3dVZSiDw4pUeS+7UykNuIXf
/IFRquUxiqqf938xLqWYoJyfu7XCzNmlUZPATbtvsMQ69ZoZ1iT98qVaopTQhhYl3LM1XfbDsKsT
t9hLXDdeo2FRucZ1sy18D8uoR1449KidIi+P6c+8XnfXgJSM4lnShkztHeNjl0L7QzaQcG310UkF
HnH0kOL0HQZ0JpnO2e7EX3e9Cu9m7pREHBzyxKsIs1UOINDlyejoG5N5VaMyT2gKwWeQrh1PQQhI
xwcor08ekvjiQ/3aMEhXG14rB28AGkXfnwkCf2ijNMsWaLdWiE2f0PeVZj62bSVhzQY4m0Y9KG6v
29sHnDMCpcFBal5TyTBs9nUOiMenZI49RYHHBN0qE/vAOUTHZRN94rDndCPqyxXyuJ6xu6iK29jd
rbu3GAzZV/COTHuLmp34FrZrCvHeTfTVhp8FCfuA09U4gHVmS10+NxD90TVih310fOQBA+OYXHCS
EP67g6C3s4Gs1/hKSRoKeEbBWMW3BdbL/e5bnS3df19z39gkuYJd9E6TvdRwEy9fYOHRjAXQ5Wa4
2gzxr3zWO0cb/5SMskdMT4ea40n2o8cR4qtY87xVLjdiVzI7gxwYFYk67g/nqtbhZd+TNHy1Q1Xb
Lz7dnpx+r1OKgR3Fd3xXVY5OHRsvkusRsVClWLCWtsycMGrognfK8HshtTgcyH5TsV/0cQwOrUIO
dW/6ynoCELRVf99HBqGZJNy+BvO4cWp2vviSFHuaPysL0eoKb1DEMl/H4xaANAWVjZg9uIOxP/ty
OPlrEgJB3Qpxkf0MpudEAA48fmrCVtKdoVeZ76B+s9se0UkfJLUhxfOz5Ept6rXXSdAGYn1oePGc
VcqiRD0HAEV0UhEIvIubB3ysoi/dm+a/FPGDHDmhzeqjpGQXhP0jLa5nQc4KESf2aSmLMb3ZKom7
Y8/F7yy2gT7jdQNkXoc5y23YO+o0rrxbXBL5GsG1MgRWE20d7Jcet4pKVOOF8102ffO7KzYNOA9z
9sMM8dyjtBcRWGPu7YJ82Nw3RtOvEY+oJAdp0ad/qAXU10ZVaP8OuKwH5CFZ9n+ReXdd2X7PYqIp
XZ5aPOGZaVinZoWHajOiHOZtHr4Vjy75IITV2WxrvgK3v21wS1AVDjiLB58YQAyp7E4z6AVO6k0R
H+d+ZXUvPwYN09WzhZPv784Crxq0hmkpqsm6EtFCO55pWoIhpMQBPTzAuXzhDL0pJIgG3IC8oSA0
uiNwoEY6VMpbhbhczS+Msuyo3NOIKuN4DOHe27CjSMQ3EEl90h6JmzXgaFS6MTTzYAw7khBF7KtV
wGyXimLofyOspwSy5v98rDXIX/sG9A2BNjhmUfoSeH7kBPhlBoT4Fk5cN0AzbVVZnaA/20FZSWe3
zC+3SIG9Tjf77BDT36mXaRf1pExFENQJqHXScEHk7pO0AC7il1InTSLBodXkIm5lXatrS0d4VOox
iuKmJfIEc1L2uVyaBx2bl+c+Fxtn4rRgDy+Q6LYhWtstEtvf6BV++3hBsZLO8rjNELxgkBlmySuS
AbtdlRtbriiuaVdRkj4ToCIHmE0djvxq+MAdPR6CL1HUW/BYgJavY9nj7dPsyxyXQlMNqD3jIpwz
a4JWI+Ct/Y4BH6UEWl+ockSdpFnr4O2p5FdeKJh5xVPWtWsmkN/kzZXIcX0OW+GdSjaREqlGmThh
6auQvEhzcRG1km6HLYiBiCSilHoIXAZjEbrlfknmdE2HRSDLMdpFwZaMWFYyPrw6q0cU1Z5CFSP5
0yg2ATI60KjIe9fyXUW8REaOglN4YuzUZCPlkDMoVIEAqj+rEUQGUUJu7HuYuz6vLCmV4rwM8Ll/
93fiaZ/bEABfSf+VJihovizX2Mt9cFBAcff82Ktr9UA1zgCZoDXyx4812xhkZ9YhbDpOof36BW6o
0a6TaRFVn1KbNQYFhH6ujcuZG/SuIUieKCaPmXU9AqP21TF3/fUaCYgoVAOsbFFzMWQvnqLfONPj
W+HVvgyy4R35EbbWgI6a9TilCh+jM9eHQxqBS3bz9tL/0hjvrASvYMLOeEEDChxy7phv0pspND1o
fM540qpPnoibDpEsvBUpsv9oJBYsPEczkAZaOWuMbDdcsyo234ySU9w04U/KoT6P15G3rGEdzGSG
JlTi3cGn6A+4Sr2RD+hgdLKZ+l3xkbHQQMw0V2SJPrn6NxKep8fsHTf4O2E/tOKEd+mJ1dAt4GJc
SmVrMG07BBQ5HP97qGzeOOf0IuvO0PEPnCwAS+knoWVg0hVcfNluEbuXUnnSSLPtq912uBiTtJw4
dT0jsLMqMsdAVOlaJHAwN+S0Sja1xcqJCE96yCCEb/JalU1u4cpB6wA2FM6FkH3UGnaTAw3Iee0x
VSC9cBY3e+uxqdwJimUSowPJyrk9xmGrxI8xxCz4i8Jsdw9xuvqTUwjgv44yEFh2bjOo6BCbA70K
FZN8pgX6dETeuNeijYhH7FPH9SIjZpjzRDem3oy/eYY11EFkSYQSdDwmbpvtsoqDfCiaiChDbpFB
YIEpnhB11pNvpInl7k8TWFvovcSPVDZVaVJNeamUPJd2QNUd/CS0DRH5wb/eIPiuf1Rbq3idbx3V
THs1yryUkmKfYHpMuHJawafLupEVR68zORFvRtqCEmlGYm+VcgjdK7a3FgzjrvQS/MAAr5xEBFgU
RBHGtvCHsJJvNl+yixCmczYdeuirSh+dVAuXjac2Dy+2BzVYj05rlLzDApyLOgH9TSzp+H3jkcMp
MuxlzKUS8GAGxhj2lF+bmbIp+hu/kyQ1/vvLGt33sDTNI+NCa2/xaZp3uCfcdNmXv5YcDGNKSWWC
wGzvefl5Jh+FEcNsQeplYFkc3Azx+hBi/el9eZ8RKq0k2mIJgvdKw8r6i95Wx5VV8qRf/fEOiDLT
s9siTS9GHrPRfdUAY2nQiozOIEKUFOzgqzRunhvqJVA+L2E92N9zGmyu0qUxqPYkw9pYM9eIsY3+
aYo1ASb4gu8KGNLEAX1QKExzLMkn4Vw2C5Ia+JH/bQZ/HKKzCsuvE1BqGsNnNqdxSNX7sOgIQvUS
7HSxq1TIFSE2eToUBwyzkRr4JKk6ue2qw64WXoHL9SCxvehnHML00dT3Dd77rhDDFPNPNkNJvni3
YjyraubNT0N+HmHOFo76MjuilVKluot4vZ/9QokaaCsncAZRfZtVetyFidA/VRepuUB8KR4yXqM1
QS2rFmRy0z1xoRfFL9jkVOswdLI0bfumbE2GnYYEM9FJLdAwnxik4WfcnbBqxVyCXIBN7o7WgykS
XoryX7NtmU1t34aQgnVXTRrTi5xLSj8P5o3U0QkVtNpkNTUYFGpTm4GSoPGM+7HFiPwWGMTMtR4U
w4lboAkIHC7r7BZefI3RZe9bondLIbgKl+RAe+x8vdwS6vae0HxBsCf2XAKsOHW+8xrtnT8iRS7l
FGadndqm2p28diNmyMav1f17b30AVpkjwL738WT3xKvorYCxZX1n3NFLFTD+oEjpqHZyWA8HOGEe
kYfc6EWLN1TPwaqgymJnavr/yXvXVHaKT4nhzgI0f3nHs+oHjd12rz+KED1lZuRJGm0YXT1/QGUi
Q1q0MLFKlhn8u+LnySj9wOeYkSBGMQu1UibY43dvvZxWYcw6GEL/vye/WswlCEbrbQi6wqrR8XNw
NbTBIFgGKiKiiuE6RoIt13DXB/an3uJ7XI/d/pchOCzBd4JJKsdVaRkqQbJ0Fq0Sew8wry5flygD
hXqzre0CLRncqSaoQdKnSqLVFZrK4IFTJMsbbUJzg215yDLoQC5cZgKbDjBUrZ2xTX6MRL7+cg67
LJVhxpl8x3u6tiuUYtA1KX/JUb7T+LPmEmnVy4/dE+D1mHLLiW4j8AS6dVnlZMxRPQguWh+CJ5wH
P63NX2hkCUM9v2bVpYYUinA80/jx5nrQwKI+o+tUOQQutOaTWiSLCNL6M7fQyxUjSIlQ+jmO+MGN
RUlGk76cTn48ZoSzhreEg6Gs4zNAX2vDqnZbUzVlotXiBmXvRNOJNFUCkpSM/pazvKDR1FbGr98V
33IiN+2B09CQlJIZM7y1Oc0OAdQfhvptlycgqVyBnpj60ITQpgzXKIjva7sWFyFnvKHe7zsCqAx2
Y3/lz6XaP+FCTqR0awcuJpVq7DypE1sCadPDQn12HRpWQgqNcdX2Y4Hwp/RghpZiUqb5l0NMXHxX
EjyveDnhy4Hgg+cLq1UcqL4aLtwPH30sCpaY6WNh/0wbE8JU76QUfZJyo6FuInYzDVuaiIKORXNe
b3WYqGjBqnYyOGa4AVmAQP8ANDbwYquSAYeJKBk739s95g4pJ/AjDxa57zyoCzaXhpGODxCofeuK
w9qvknScDwDmhbXq4yZ6b+VL4Tv+8j9msUR6CG6P2ZQha0zDJBrGiay7Ew7EtSRMXQ78poh79H3n
ClOD5F9FYep2QAhhdrkaLraT2gcUmrEz2s6nG2sUWeL47oE7QMvZcl6hjjkKDL2W0aGt7nbtZY2L
VU5dTALnE0tjP9QblcydulW7Blf9DJV7DEJkT35X6oENfMjyAh6UMZ9Nf50rPwouxEijS8kozdOW
CsJ5UK2WQNsp0ArO7XjD87HCdlK8B3YXePN+/d6ueGHGelCRBiCpUJAqT8ceKWtSne9qp6w4Iznc
hgQ19SdcFmXuE82qBtBMhuY7InR/Xmu1KCJSNqmNyKkqjn7KNNjRIk1RXECMMs8bFzdBP/lSIuA6
zzE1f5k2E735NkXNCKMstjp9RTu4qZ7fynOIqsCa+K1lQ+45tXQ+akpSzAhi1K3RbwJym27+eadK
qIrF7gYpEHjZHJYz5B3xSp//2o8qYcbx+DOECeZ+P8Qp+Kao1wWqi6fIotbBPABzdRYQjWZABMQE
mAPvnOfMMd1cKkWDQYSAki3+GbPKir+5P2hwzsVtiFiRfJT0KA8kziN2w5brAxU/Pv1olhY6a/G7
XRV1TXy977YzG2QtiBfOuG5vX0ZF4/E3/Ej0nCilzmBnQE301ELxZvTJ3tAgwfuCUzr3ltRsS5Bi
zMZihJrgcw0CEjEQqQnYPq4KpWvHf2AQt6YNw4cD7mt+Oqm+w68cjAIy68aotZ4zfFg2twRAsY8f
LgFlFR1fA9S2l8Y+ky4EvTHgMAI65/ukY1UusVjrhNi+0CgkEaxHPjsMDsP/ysTkbjz7ZYb0/tIY
oo4IWioXMgfwztOqgTreZJOQBl9w55YecWeTXDfBaQlrKqtQxzPYb4vrzHCW5imwdR1LrseHZXej
kWF7lBWwAHK+lOU8Gv4HDJS9MSBUvBUYdNuiQ4t8G4MM3FkJFqWD9LKhoJ7nnIxGh8VcEzPoR+2c
bvVCYkY1YX2sI6QGWBJdZQggGeOrFdH/MZvcItz6Pvn11PukPq86XyMih5lrLdkJjRM95PZRZtJs
hB8F87JHAB17Qrmh++XTpGJrzZUxEIiOtIKQhsIkGsQK/8AWJlDQe8J0hERS2eu9rgiiPgxwm1bz
jRuG4xG6WUobNv0okb/95oLi4oXWx6OTqi5p2wQhAts4MRIWyCBapM4ayRp1TqeCWtuD8+WM5o3Q
5j0DrQFnN3NmheL6xr+UVdyqau9X3MHb4WnxR6V2CC5IER246a7HSWUKHFz/2jy851rwbkoNLUPC
4ZOxXFb5Y6Dbbfp9CGVJFJ/VJI2Rv/Y6l2rE4kC3DXBZUgDaPB+v5lpKhXCLgfkWFZVUQuxenl09
528vllAVtb72LH4ctsePzhEU8lLhkCH7hgifDyyQxbgziADOwBxw0YhxspsAEmd3evJ6GtcAYQTU
LGRyQFcIDJw6UQStSX7xmWQRrVSVEjaVVAMaaokG4KjFb2pHX9tBRP95XsbWRCgxPGgLPge99ZYH
qHke/5tcwwm0Aam4uxAEndT1AFsZqONSpBSDSka6k36usZtFZcAz3JLtqG0qOqyOSVLHya/6ekPy
bQ0Wxnr+Dk/z0MVjgvEdviGuy+Jnw4Z4zQUKo+qyDUoHW3PzA3xd569uXPabIVXTiMoXw6vYpHyM
rvz5hBIcBAnSscLpJsvMezd0XlfyHfn4V70ebcXb2NqsoxTSGr2LFzHHSk+aB8oxER9IPwWRvhCr
dCc2wZZ30a71l4n1wtQKhiUnxu1AQLRV0yhYp/CkNN+qJWZiepbVknlL7UpBGKwKOeY3usz0oowh
oaclNeqF+PzAFu1k7TiGZ6Nfa7161VfBr+C/wAAVRoawzPNFvzqkGc2VlxaS9LotdT/R+uHd9G9M
hanBtCGsbRR4nq8ZNifpYwnll6w3fwzYhzoSlGaoj8kYvsxlosxT5/s6quppJaCwfL5NPAL2AarQ
+CC2Wrt8Nl7PjJqDM/s/OffB7JBaaMsMllsw6ER4HVrOJgPWwY9k3tMQCrorTb6u63e7r6InwuWW
pGFSTcEqii/PYV9PtVT3WjqCTe7xUruhEbjrO8AVLmDbA64q9ixqzxPBauq0LvQxLsNlWrN3XuHt
SDlE+iH7NURXWbqDoBCrVlbmkjPMsC7k/IV0pE4RXjUPYeaGF1SfV9tG5B2QMcwDWvqpDNV+ZHHn
8s+0RFmPbtAgXNHO9lmOEdJ3of/tOUx2y8x9onpWcV71RHqKSNQtfH07UwNTNFKdE9ULEYJ8q8Sx
nuHQrEWAnn2vMNx4P7NbRBQjlNThqO0WhDDYoqclpa4dgrhgUzha76WiZ2OfDQtuJIw7cuLc78EV
r3/JJmh4rPE/5zvQlpCTCFuUnHT2LQENxPMF9DFK8n6d3F0cwQmdGfD3ZXWV1aSPPQq+uSOEtpu7
epnP1IgpT2JB+1AFbwu9DsnydXYVByUZHQ8TvjPeSU/yQXSRRivvyMcM5+eHr1qEYKxzf1ElMxPS
byNKIynJDQSCIRLuZoCnApuVZfnHEuV7H8yz8WqplBe1HwoTMXNWCTBKzdzbhLgUVRuxM57lZxuR
ZQ0iEe3WHIaAeB9rriVs03e4AeDZVfENHGUwyvzNE+WAcZt+6ZbqOLgfzX+FdwvySMDtcos896Yx
R0vzOmmRs0yw2hea4VkDkZm9jTRQM5q1QiaUiBh0XJUNTQvSuRDirnhQF4SQb3uQ8ZLQoLa3JpFr
rkhTy2YmqTatwQwZJJHaRcJQGQmq9lOiBz09aGrDDCcOv0I/gqJaRwmk8m3bRN3Tr4RWddTJ2XMQ
nbE7eQ2jpR8KVSLA3VDA1+eP2E+R0pbfA5HXfkM5a6oDKkKr2rU7FNzHwSqTXEjWROjiE9DIeCsV
g6ScRFvQCbBSsML7OmEEIP+di/U2VcaSZVUJVEqI0FdVcqYUE2DU3h7kBJiBQxaa88FsNcTacJsj
B2UxIGJAKqElNIpj7v5se1s3eONS8jr5SODbtsuCC/X63ma35R9BZBOA/1g4E3eONSlVGEVUPnrw
FIRWfV6SA7mrMGMcqXqD8hk0HY7UfnFJWppmyBs4HK+7MGuFD30sgWoCW2evI13X/1HNETgfURh6
VAdcBOMSBwlCifxFkweW9tntMlCfw7pIzSmKlo2cZQUuL1shK+NHgM4+jKkUOxNkj4AGKDbtbbgM
2jT204hvFn6KaJnlsgsKHUuayx8JnnIKU30zjcdtX9jUXlzl0zvdYkFKmQqGzjsFWYfj21czCBC5
YwT05M4AW7lHlOUvD/FLb05IX630nvKluSRKngVSzavVQgJxlxqyqnCw4pi0U3nau3a5iHRCyjKf
sVqxv20c7zM1wuzDua+qpUMKxwgUmptWOFm+5JwRfaJDq8zK9uTGC9/iio/qdBd439yc2qPULEcb
jItmMDUAnNMAG2zZNjUxViHaUYxlJGBHOJXtVh9+dcs/oM9MPJej8QgU/xbxw3PS/ET20NVg8g9x
4Xl+DEhrRXBn7O74RWHXLaD00NfH6YKQOcySKWJsI3qaw8rrUz0JEYrmpcWMeejoDsU/N78dhill
Gt9YBcX0KeRUw7qtrd9HyJ566AoTBUHSH1hBPXwyk8L+3YYidW5RPFCr4m+JG8ECuVAiqnsPWtgO
Ml/R4H1fnCNZR8qlvbafCBt3VqLxBxxMtbnG1qZyRJh7jtuNWRwVDWq3zUWaQPrNqwkdsfg5W8af
GNL6287gNlfUIBxr+0QtaiP/Lx3Hvo34N4H0funQOnMs1Hy0vRf4Qq20j36vvMrsROs1NGhsKmmR
2R5UvRIRbZxlaeg0VU8xJO+bpPNw7irRR6iH8HqSOOPvPYz8QKoLWI/ZkS9UlRymlm1TEuiHt6y9
pRhoZQs5OwQchjD3zsUd8G54VCGbGgInPQabp69akLMSp38ndb7ISsaqcRbVgArb5Bxvldtsv+R2
TzPFiGtJky/o0/dXcwQaPaPnhm3R3A69VxFIr7qQ9cYpIUNNldprej/yQ24/4p8Iica0r7GWeutI
mud6PJYBTTUS587nGtqbCnWFGPAxDh0lmscA4rbaSBesWoN4FR7vkZVQ+0M8BvcF2VbvzoNneHdR
rjHrt+pxxTXEzLSiUtVdgqt5Q2DcY8BtiYsOV8FGq3HJyi5JulXVsTKcz6iGQy5kLwel74LbSyl8
YZGKZR9KYkvDzqS1oSRKMPAnonHheVLluQ6LK583h9o7LCFx7Zae38MNpjFao7Vpe8ZUnDCY/hc3
4nFDj0/wnTtT/ULZgYCQa0sMGlIhOSwbAVJsYqHesh1iEW1wALk15HhBMUiNcpzzRfhkX9PAO4vd
E6UbfMOpABI32FNpl/xa/8e0nTm7AET/STLwYQRrPLCmKuFPocS+R0FX+se8daX2sLRNNplQ6Nh9
2twFT3vLVlFZkgcJlqqpzOs17uBxyZU4WIUJNhUotlHBqB4enc2RDLqvwtZ4MTH02og7eRgskchy
HQwbL+JZk0w2p8GjX6JZ0zZYr4QoKocLuv806W32KFy5b0abRwao0m6kMTOkkjEP1usmzzkLR4kK
1zddHZXNWZoMOetLJnZ/busXZuDZfZW+8Gk6dlvb3bt0wV4ECoYjGgu6wwq6NEBRNrA8TCSiG0VZ
NUhbl/TnSh0SV4M5fxXVxGTRT/JtNl8iK6+Cj6TAnlvP9ZIYOudMgtI+F/dsVbHo5fzUAZij9ADW
8ssxBaedHVJkAB6gPzrs5xxK2HG/vkKH+qJxe8lNlXlfeSh2zvNJc7C/oieSZraWEQ8YUuSV/Xgm
YNJriSkqUqEWVtQHkj6JYESmeh6rqmtEAQGTz5vonxatdfmqzPSEHngFravQ7gKDb5sAXQna7GNo
snpMIzecue9qVxhFB2B4KhNTDjKLwaqcqDu6in3ZqrcJ4sT2DlopO55kkTcE/cx6mHPy6vcgwLNP
gtxlXqZUcdPxlO1XTbM6YFpjGNo2YeiK5JzEpa8DVwX5uwWPVJlYC5t43MQq5BH9gSpeajmBDnEE
izN1x5Akc2Oo7MvLAR7vHaONxroHUq+WEZlJ6UM/LdQSshxOWGJnmVlPAmfWyPXZaJQr/9FlNl7z
6TMrQK/s6sbpWPqhi1U1eAgtZvRR1982NOn2iMRqAWffQyl38pE+1TbNfaRJetMvld3qJ1ZjI5Ur
wd0LYkDpEI6H9IyZ1UNB2HFrdY8DJaRDdiXokPmjxPH1KeO/WcbgDcQY0FeZ4O10/7v0oG/ke1/4
t2gnqPguExX95jxoZNPonJAsV3CsEj+DwzNKe8tksar7jh84ZcujcUOOLVwLmTUjr5wePV76Sp7v
9nPxRLjP6Pu128Od1G2Qa4HW6BYan48jT3+sBQ1AGTnAdlqBTgKJGxifLN4++NfUaCKyjN7m8NIl
Tb2VMtHBMYKgmfwAGCDDalT6bFE35Mqg0dSoPZa+Qj6fEywuz301s2EoWpKttxDiw3SiuUrbKODu
cH//HyJnQ2v1Xhl21Q/E6pVorxr6UooTqYhDeb2pDoOI7rr2rAQztC56+fYHLo7dI7hUmEi2NLML
DUrWXlW40i3ZgmOtrt0J2vWlF8VHpoa4huPPWVlxu+tkvWi+pM8vxsFAEAWpncTv+GPFmEvBN2Mq
fmdkpq8vqBocYWdyMLwTgFeQVWVuKQ/+VEDTYS4KK8QqcpOeJVW4sv333SwU/fqRuyfjsL27VbvU
1XHKR2rcTkdwc2ij76/eb4K6er8rPlLx3CW+FNIUChpu7VFpOz33PJ5GVbiZYiCHSSfqyFQz/Bi6
voobyrvOzzjZ49x6bLiFszvwIwYT0Q8lH0+l6QEq0Ttedtw0uiMaiNBBMX+4hvBCWxc6xgeP6gka
J+fjIgAYcr7prYTizcnCVues/rF/GATAa9iI+QSMm7vaoqP6aP4eB/rqupGGvW0GkVxBH4n9dYfR
8N/UD4QDhObHuWV74hl0fxhf/dpNu/Mj9OkWWMI5DxBYCdN95R5mDB5uTTcdNoZ11cQ2ElgZXLFT
SCRBm5T/6OWLOxPdnRQNCGZrGguXC/NyJyJYmG42XV0cs03tW+y3h5uv9tkABzs7OfbQQnCCh3xP
MBBFDtEkIbX2so+trPSvacIQ48OvnZQsRVzuxcMp+V8YoOMeZsxojZPgpaTc0hL9rnaxNInooQiQ
Uz1fZe3AblhKlAWDwFAKlLRmIIzIFik062ZLOA+IkmrLdQmJmbiJaUz9F0DU5vIC+JpVwTWe1xDG
0AonvN0h/4nrSh2i3gQqLO6Jhn7JA4QW9c1Pc3aLlCeBGA9bOasX87W64QJr10V+IFYJfX5Pcioh
4BiuYCk7RykeqFZo6b0sTk8oOuUd4OEiU+uHvh/OcFb6pyMmyLh/st/of2r+D2BrLXuQAKfXesSU
lZeQDwVlArTb7hvUfti/6j+TJHcbjO7YGiLfMXI1XOu+s0NYSCA4k+UX7O42G5CyxfEa66fSvm8c
EdQElwRvpmJqpRyub+GkHrrRSOzB7GuuJkIdaFMauxAHHjBWjkHlPEgMimpDnGu0FfCwPEStRO7v
6IqIxJTgiMx7QqzpzacwNSKMH6BVsH22LWg1GgAse7kRx+6lKXkUMWZWpKXjoIc1RWLvh5VxnJJs
CHkAMnxY/M1hI/JfFEJXyv1aXY1jLYaGRia3vvA6Dj6jZVPhBWPOzqQb3AQzcUELIwya6+mLnbY7
pb3ds+3s+rHqtvjYmGF/CnDIl1ADZ/2L7rdm1tgEZNIlsUkB6ovQbXeWhtbSE13/+//9pciKEixt
7WGEzciTmMhyDT3x1GpYVq2fJbbyDhxvKIZ7vLclu7SRUhPUY2VKxg51Hz754v68QBzWkZcz27R2
9DRbe+ZTbTlcfmRsetXCs4JaUvEia+eO2PsNuXEPz/U6PBAqtFFRkzvxLKekuiu5TZR8OIPEUrg5
R045eM9XSzRH0EpacabPhFtU7kdVBLpO83fso/Nuvkyhu7kQYMDoR5jw4fZaoW9WuPM0i3LHZkSO
kyZZBPZFEJu8y8YQ6BxTG6ESvTq1ox+EIHSQAB1OfIfK29mo8ODC9JwUPgkJ2qFoSlM7HrVpEQPc
coKEJEFtH7eeLDhYnwpIiQgSMzj9fdXeEHh5s/Tk56sOmEHdXVmimmxY1II8rS/35jtqQPKnyALn
KzcXmNJ60WSw5r7rstsGCO5+hF1gHdrp5R4LUDazeYZzPXT29ESy9BGGDGIv5fmnMNxJ7Vjo7A9J
uBv9fJI91k4gzMbfRgzxFyUh4R8ZspOb1vC9E3mi08Rv0+82BjmaU699LhKFXpUgA6VdBdiSRxnO
NMLC9pNqTCZ6dcbteQkilXU2dDuGAankn6qwwke7hKKApayKS13e0QBv9rMTw6cnXi+WgBYQLJe+
LCBCVJV5mpBmA1FDaVX1gWjD6ERmdkrg6UTOVBUYCa4c6n9K+1NcdqIMohfPJqWkoiL8Vhp/2DvA
q/S8HTzlIwIyxHzB6DfdP4PdaPDwf7s8SmuDRsdp7AKeuk8TOUlQIjmAjSJZiHoxPSHCnjGp2Nz9
iTiItEqWHCHvDDZeUadHu4g3KRlrhwIyECJNFKv+e3aWzt2tFIeWlITpGPNP8xLBNXoreV4palHx
b+xVDZ5ErQMpqQPgPkWO5Cb2YaqxQWxmNxLas6aXcYt740n6Qpt/cTGLi6KnR0osUuHVhNq/OvZk
3XNh905Ecrtl1cANoE66WK3/vZVoM2+7eanacq2B6PUPzrxyV+ljGeAOysvmxCs4gJrXmg6Mhafz
uyZhZDzlBRqOxl1waJwkzTVd7r4fViO+UgyEzi1rqYUfI22oCl5EuXIdlzfhQ1e6rmiXaCfI3Y1z
WFVqOkti3l3KQRb5dlG+b7JG6x4hSe6RV8/v0Oup+IcCjiDqwjJWb/n3ezgFwDsjKAAQbKuf8gGU
r420K5/FE1I5AUeYNU0acsswLyQfhceJBPNZUQ9Cp43SrvsWnjr6bKRi3Eq6Ccq6mz0EiXRAyndH
C6n8uEFb3zfzTN5uS0uitK3eBthiXyAP4Yl5qmmxEJR4lHy5Yki8mKuWfc/3te/B5iqX0vrFQf4M
x9Ks/7UvUDevHcqlh1oBNCWd77lbnQtZ+CdJVh0oGd3NExRPWFBYORxLjMwxB3cupTRN1i8H5B4i
HumUuMTCUVoT8z8SvxttJVHCgChHtXXmS1QGguWObwQeNozdAOQQrlONIgQ8nm7TxYnNU89jsib+
DvrdRC9bQJag/TUT1Ncnq4+02Odr/IP6pyBT76P62Y2UAMDcOLNc/nQNOMaz2zyGGNbOPBU6z9CI
owg2RSAmoaBHMQxYOmKTTbk2nuaT8nHfSNvFXKsxRyS0C+Vdfe6ajiS13U/dzPTDv+dDQlrFOQ8O
yJuDyawsxoCpFqh9bDL9pTxRa+om+dis4A/cMY8OWziDjrYS6pRTV9HiXzEk2NiWI9gGZXNF86Lz
J97uFb8tFrkqJCWha0xqQ5BhNrR5yQZ9j5xsyNoHaQupd+SBYdu8gSg6thdJDc2t/vJ7L0vNjpEX
8f+9zGjaIoJvS8tmTHrn+Vl+3+vTSvaanRYZSZMsLYpPQXFkoND3nA34S0BGKsjJhosE7nA7IQRo
LsMkbDr/W0MpEyw5ntNYD3buodnS2KFkQXVFyi5K+2zbmXRB1BAwHTanOlYIm1z2Qc2P50c/ZpZl
XOdknFd+upeGNEfPCrbtqfwn1FN9qKqnsl/JDdXSXBGggsmF7v03SjnhUSFpyZqvtLPGo6PQRQMv
ECwGQTfCFhvpqq2Yno84drM0zhE/fs9P4c1NZxztSdrTILzlL8rD799cEKfqtElgxINq1Ih+XlG8
bV8b1ZgJpwoNGhT3LEyGt38m76SKK1pcKriHUuNWukktj2KlV2oUDi+unkBW/5AKWMS8Q/Y3a1Pr
mVCA+c4rqMNBqMPvIeSfn31AR7MW0MJ5czvRFK2sL3JO0ogflEsurc7TN1ckZZU+c0eexcwuPqrm
iZYHKLE//9aL5svALFoBBnkGRPxoHeGmKM1K55RdWLgFf78h16rIVrBrIo6pS/NFAGBSK2g3QEmL
wq4aqnbacpZqrLJjnJ4YU8WKCx+G4KyfeCZMaUvkPKMKmKXAwX72HJz8q8OKKDslTElU2/HyP4xg
hmhYAnY5AkhVsbtvIAY9atrEyNrH82luFdeGmpLL5zZ2pWGVyB9Uk9X2w79drejIRfm02v/oU9kf
Kv4C6KNjKHUFwET5EO1MHt8WeFunXNkaBCbdDQr3XXevukiYhyj1/ddQKsrCPZe29QQkQv6Zd4I6
QPM0PCM6i9qYB/rk4pX+PQCZkav/j1D0dhZR/HqafJOej8ju5TfIDeZRZNWeWKJVvgTpKQiwPFRl
jvo0+K9kVe1G3r+VJ9jX+1Jf4tKUFn31x8kOEXYXXVVx/ELlFjNPiFjKibV93wkDSlOzWo/hu/gM
rWwqnOY1NOdqeJFQv7+XWPit925M5JfxxLXjZWypAg6MybqFUNojevYK512MpxEfUtD0ibezCmbD
xXijH1VTOTJcefW0h1/TDyU8C4LsNRbOVa9cErfjrQounw733eRBRU397ZjEOR3/vUho6C/z6Qza
3sipxdri9IA2gHr9ZCk9qVC49gCgeNvkFxXasJwoFXb+X+bMFQAl2+UztueoVBcg+WvD+itpMTyh
qbxaMnnf7r9J4IXFQiRuOT5v7bB3sTc6FaIY+ZgsUXYAuxvVSTf09CqWS/UxUaUEmYd8pYhdMF5z
aR+W1FZQdVYLb5RD4Z/DJM4XyTxqqLlcKCTgXoH6J/SlZO2u5stVuBCPQ5/BDCx4997pzh4IRnAT
ykTVoX2fQPkNmOUYIkr2yhWWtDJMGKlN8818cnYfT29FupUNNCClGwjVHeyuBCNf4C8W697wT2zI
ayzZBnEkisbtVyevOJYcw1yQZz7nAQGm5/w55dg1aHEwSHVKHrNLLzoOCs3uZpI3K/uHO2Lw2NFh
09MPPUsrFUNI6buLF2sardSxLR5FBgQ0X2sHbfI5UxGbyNVYjq1gWvG+LUmcA+/Limz2J7EEjW1F
BjI9YARfPrlPrSrP3IzBzYwHDTT5Rakqqw3mmQzeqQc/+T6gLGAkUDUg1IcoStMbDbAEWONyRMdA
Om5xxXapSDYNKk/6QPpBaHIOcgbWAdnv12NW5YkbHA+156IwePiwat/Q4lcqhZGDcqBXPhZeuwDL
YhS0l+P/DKywaoz9u2U3RNYzJlXfCX0hcHFVMUjaC+JoXQ8/OE7GPSMNCTwfGFaueHUugjYNibd8
+TWd3HKwjq2LLooR5MPUL/Ed21FECTzFhuUkGGmxoaUMO4z7vvBB1MWcFeCmoum2jzCj2fYXucrZ
ldzm1RSXMsOaYczTZB9Pkqq66ZaKLkKhe/jnDzdHziVxNbwfnk2h9nD5XdhqAxDw0JHKLOUlsRfh
yW6syWO9zJHYr9MuzegqBT4AqsO4yyyBlLFGddal+d2bpy/VgEnJw5EPA/DYtqEF30vNxZNofRfp
xzT74Plb0wsmPfd1SAdK0TIIWHCOANfqREqLmq/LC4EjzjFaxIRosMvDlLrHtKFfI+QZgaTeoPdY
U/H0eJvfVzQAKPojNaOfYa9FyV35+Kl8TYlWLvfl6ROihqmyYbcGngOxm+HG645HYtpeIMVjWNps
/J0zqYdsy+1PrEZ3dhHxq06PSpMk1XBTfYYo7kinsOsPW3f1lGEmPhxtIEUgEWKXJzUerq+ty3fk
+6Dt34858JocZo1mfF/qKTs19zhJEwOxrkMB1oMKkz6u12TyT6eVEHBqgbg1JDtebdtjD65HJUN/
175sbVcasOLSd6A5hRRmsQVGADDe0J1FN2iX+HZdxwhi9dqmnWAn3oU1sTiQ3dQcVXi9KQH4t6sw
+aelJZ132qTsLV9ZnZBD+Z/LgVH8LWoHSB66XH3imUOPKaTxzVIWX1otVNqixMOaFJ6p3t2Zwa/R
bOiWEHplX9b+4PC7LP+ZXd4d4JBtdAyPfjgEE5u+Th8cVjtB7Whb6s8CZ62/efBJmKzq0iKD9jFP
ltMVE6HxPb/epnaLKTyvj+v2jt1z6bO3kP7aZg6NSMIaA6m0sMmBGXJXGO8G2tinLcZEIcRaPiZn
70JeO2TkJYH1Gwr82Tpdw/wDDblfYtsBtjZWa3TGxsmlbgm9wsyX+oQ6XrsX/FV0rR8il+qsQToz
9zHb3nKe1AuxzIvMwbbVTaKFFM4iz45hhKLU4WaQpIHDslXmNqZzx02u3h05uScL5MxcoIR/cXar
I/DLsFz6GoF2bbbJXhtgAw65kgs2J55MxdUNBaEpzKQOgY6sV2GCv0UjUYcpAju8KvL09BvK1Xqi
cRzy7gri5ji1/5/xX/SpO/VVFAkYA7wOM40o9Lshvizb0UJhyJ2A7psREFZlYSolTDILfJIAB4ug
AV6EZTHY5H3a4a7LZjhPlTdB3VkjXoaO9lnQt+1qUEWF1EZLAE78YylxcEvgV1ZRcXsLXOYsqoAJ
HyJvdaLFsjNnTASoHCdrcKo6btOp9YlPy/nqgW6MgaJ1un4LSaLS8pgp9zJY4Sw2QTxml8QU7pf/
rAG4RFakd88ekO7MHzomN+jIQcjy+cli7DdND/68L9JiCqprZ6iNMXvmjAPdKrtz2QlFXEJz3IwL
VnpHh8We78bo9ZXV9Cy6zE1+40MpDtE6V0U4P3DNiW+JwM02ZZaBc+tJ54LY+oQ9UHXKjVXmtrBe
kj3/mboEzuz1xPNY0/sgkPSZaCtzumArf/5HHyK9CPTYsev+Az3svMXgQoqDrwTRJrGnXDWw/bZR
4SDu78TLaRezFi/s1LDA7Ll/wUd8JmOLNgFzLCa02jLtqR1N/R6L4fx9z7jjWWKB4tZ4rsOERJgM
+Q7lATxPRQDuSUqh3IlzjC6BPTByeeUn4rsCdmCxNwnrLZ2u0wtWgFRenM//17IUJMXynIi1Sxf4
jrdzEOUGYmZxqOrrLZjz80JnseTwJmP3LW66hvR3WmHU42KzAe26TN/T2kW+7FrZtaEIbqfSXVEF
8kP/2xwd2luGR6uT+aYc/uXAaj1liaQooBuemnwcao1idUAhKSQw+YcciSOIbQMGzJEM6BdHiPOM
pvoPZhoX7sdbgF5pesPJyq9myLNgVaT1hUGnT8OdnATrvc67MV5smLEaVxxj+K9m58e/BIyuMhwJ
oJpYz21XPCR+NlxWAZFNA09WJSz+CANHBNH4M550kXJIUa6lbdFtD07BJn9C6rFxXg83a+Mgmycn
3HSDOTClXFxonbruj5ecmo15QWwEukVh+T9x87Vy4rqcvKock6dlv91eFeDl7TwaC3OLvb8Oh5V9
eXpe6JNugDiNZV2giR70KpOnimQ7U0IdguqzlhMt0+N9wOndZpwPuguXEBdRVR7chkf+HOjIECZY
jfONaiEVemLjcrk7QJnp45FezM82JwTuyf6TxGSAMEd7rQsLIh4m1peCCuTlywZCqKkNDlaof7Hd
YOf6sfpqwF+1Ngs99sSSwRDChq8d4jIfWn1VKoAVdgmfAf7fHPO7Dzvwqaf5vJuMYA0cjVFMY9Qt
aAalcnDUDDtOAj/P6ZlasaPib54GyuE2yPWBqSBT2vKRsrdz/+pOEDFh+uPizi5EFu4DtsAjHUac
KcS6pYCmwYzIhnN0pBvwemmsEcCWJI2jkTvZS6jOyVHTzXWkAem4RUzhfKdFdzLMAh+Z2CyzpRKw
oOTwa3df6FMSYzTABmW9Mj8X24aQCUeOX6K5DSSVkJjovi2S+fd4DmepTFlqU01WSp0YuUp74aHL
Nr0rxTugg1AW4Y3sEyApDPnKo8Q9l6/tlxrQJRyLFwZziIIXqdbabFC43054J5uwko16qfy4AvKh
66vck2lVWLZPMoA8LCNvrBYJgrvhi+Uj+TOrRp9kF5Ai3PEX/XlA45JSQM8XkME16N9QAzTm1Gta
CD3/arHpB0Ufd5SGvascoOIbVVZu7GP0CY9qPlMjn8mJ6gqG6Px0awdQp2hGu+63wx5WhaQAI9Jo
TDpvqrAC/d24V2rGC0U31UqVzXGUDSn+W2hxx4Ewu6Kk0E697GlY7TjtmFe+eUtg+KYOGqbLJ2JI
+GZTalsEeCFcGhEwaz9vxvvrOq6Jvl5srfYNZ1Ti6+07GH0MxYS2S19Wa7iymamtoWZsxdpk9DzW
yH/jPLPae0llWyKCBMDIiW/MX3tirO56tf2fy8QBc+orZxjDfaMKN315UD2QJ6OY7y+YvQ35bo+Q
Ald1VYLgK3VV1PX8NUjNBlTohUSdVKHyLLLMzit2ZTwVkfYXYWG8ebEVzOocU7adFpk8xBQe2CTF
bBxONf4p5LfYnrl/mK4fv4XiIKuO7JsVnbGoEXYpMfGzrXWAnvXCLY1f0kqHW0jkrlwxjDzFFbt3
1ejja7qVxckINmv3C0Qk+xak1HL5mt3WcbolENj8cVYA/tfM/3hhYDchDDgbxVnPa0dhM8zGrB8o
VgYXCh8tzk/z8DSjLdTchD0I8NSUBQbH8mvuurXioomGnrKWjzQ0DDhOUk5uTkeJf47jarWx91wk
JvjPgmPD/SdeFb8sz+Mk5uTl5GW3khRtWJ91l6+vx6OxSRKWtCF7ZnDQZ8p8YO3PuKaKRqcUwFue
wXprvoAT6GhCBEsNfTdOrH0KChUCiZkUpZ3kllbX6rdqY7vZoHVEBqZypDV0ePI1A9lOntJPHOka
hqz4kvgRQsZEo8l21wKuHZ+VWN/6iFwhn6fjLPvQrmxbAkt6B+wcmUzKcuoDvD4uK0JZNhxaHG1H
E91zmEuIfSzqYqZpYbf2VbwF7hFYZOSmK7ZvT+44mr/EsVRQpU6giZQveDV7tCelPBwyq7E09Rmh
2b/w/0HQqcHhAFextVxwGMbcLgw6LMWQX9DSVSqySMszh/EclIhB2l+GjzCqMPGNJKdXprcwgXp/
yyARXrGiot1sUgG4bFlzT4RhxZhzSgMeq71OgteJnthO0MJjhuex098FObVLV5quzVQUTI9dkDzH
9oWZ4Ti7I9Dppec2G/LSPvpwafxr96xD3zw6I7hF7RCaUXwMdPDm39VhJ92zHlmf/5g3E+yXRYwc
Vx1DiXEAKkNmeVeeJejKU1Yt2sBHwYJyuXbDh2xDLOsjA23uYaxUZWwPLFC3F9xcKw0ygwqgr9Wx
Zbi/SQ3xx0d/nL7hzLHAYiRoFBw4RuxV0kq3cfcIrXngwCVxEiJrNhBJABbsnbHUoYHFglDZxVnC
LWTSEi1eEnCTaM8GKUnT+/ICaO0/jRt5P9smW9nZJbZ7ifLYR/ppW+0YmKGAULDtRuI/KQ6sDMBt
pgENCeFoHDR5COsIUgZAfd/jhtiGM5MRDxDciYHvJ2GPHv5mmiRfc4ajvT34PGZ+xNrESAW6V3/L
Jx0zZHSqkXO3z748w/ztYgE8GshPIm9lh41WdRb6OszdowLi/yed1OPp/zUjsBJpiW/qPD9e7Xc/
JecUyyRrW38I9cuqWKwJbrBDzDXASCxl9po0LAr+ovSM70RpscKUgwiVyiwq6NnoosD32IjEzzY6
jsBKzCEI7bKRz8UgjchRCF5X8dCt1T69/A+Ce3H9sbSlGIOx+j1b+yOxqCNbQqePfs4YDNVcXygg
GIwGSZVHVdkrNYwYH1k8M4BShgytMTt13wGrvHXWrbCvKF44QDBWrskAOI9LmYW+VdmK1Iza+VkG
EdaDlVOtytg3evkWaTLHqTVDLYs6hnnqHmJRVDvdIuxyw69zIaPTloMliQkhfpmhYgiqF94xoifL
rvVZHqQFy6s9yQstKANlVhDWXccJZ5+BgYkpwiLOD+OxqSDt4O159+M5occ6hapigaJ1eHBdsIRH
1dlgJe5us+vZfUa0iu8F2Q5Q6mhOGGUcbc/CRbGZO0vwvjfaGTeB9QL8iAj2jLJFFnoYbkz8jWYK
N8TWXmrRMNjkhTgWGzu9JodjHXmxki2LzRM7Wzce1MZlTz46mwjKG95D7gkQa4R6LOAHrI7jWwfM
7DhVmMACXUW2yERbEJubxXPF5H8cDFmEGt4vzbZ1Do/35YVwPB6kzKR1Tb29WTW+YUxk17xdu88S
OFN7Wmsh1n6ES9skA91otQpLq36ph9DcPSzQ8w6DadwpNxC35sdRh12rsmJcfY6mm/W12TpZGjdi
eMKqtH3YwCVQFH6NQHEjszucLoAj1dXRFYFs4dpMaxv56N6rq0t6rr6xrLs45aJeEXeDyJ7WegGe
K32d6QSfVWTlHVdIGU+OWzE+ft/gi8KuOE1X5MC9n4nnOg4a0P2Jx91grGcI42q+ytS4f1pviPKf
C5tiL+m7kEFzQXpyGYPxlkYdxXZD3TBYn/vU9AVlvQ6DbLzqnaz3dlahbACjWXsdRdWchRZt6ggy
xndtOo1PxQGEQSY5WkPXw1jAli9GF1bi9gB632AhM9yvwLmRbSjAlI/XdUBXQQZI2WYqyfZaGY6+
r5RkLMPNTGT9TGIGFnC+7C3M+GMyrEDeyfm/JJO+qZbaTWLF+JtqALshFeLV32W1G0GEilSNRYFS
tvneuId8mXSI5i5cLB3KgOM0ePB8YdpSrwoM6VcO9vl4gPZbeF5MOAPUg0H55s15Q047sP19XFyI
gvJU/ug9XSSc18NotMmeAZY3XXumvY2oVaOb4c8YzoauvzCrWmO3gOH1q9SE0G2bWXJ3UVcIeIhd
ERi8tyoPe9f9Nl/Ben/rTebQrWZKmmeGZfoo49ZiUdieX8FcFl9k/oBFNKGquc2o0Y93hMFvfWlv
C34KAi9NsRdR0iR3EY/D7C38Vxl/0suG+tVf/28WR8PHG3tQoqufkq5w6hrG5csCaAotuLYzF0GN
6QQE4qUEngz8nGfFegWlc6Yx0SrFjhyUtiotaErQbTAZ8mb9pvJDPDcw/zQab/WL7vAPPrUk4ZIN
4Ll8npGvVa6QruYHrcATvj60+lOds62tWSjG6Vxx5iyP8MA0BHbXZp/Ck/eQzpbl3wxiJYSSrfOT
SoOqpkXrkTHdar+bG8yb9i89D3TH2zpu+YfLz2avOMkaEFZu+UV1DusNGmrPcH4XIA/wYph+OSx9
tGuOs+8T13DEZNKepqyvXXrSLa4iTrBUTUS/CLiQ1WptQ8MnwotJaHzCOkRIHuhW8krj+6o+2AcI
+mcvBA5NUu9uvsQduSs8l01z82oC2X/DRCWeh2lkrWWHcgTEH4b2rFy00bKKSUGTu/kTwAWnqHeS
vRBnZEotH1G9GtDOk4C+KTmeHzFZX6dmuDiIIQaG/w0ay7ZbE0dsJqDl8z+pTqS3jda7v7G3gjH1
oZWim6WL2P9UOwvAbAJ2gXlk/3mgsLwUsjWi2rFEc+JedqS1VGi45em7EPzV8ACcUtycuV1EWyim
vSFosyDa0iwOvxOyb0szGN2Y7VyoAfzYbOiBgGnkWQw0XMqwDcbkbaIVEg65Zyvfjvqa19VZLXpE
NQKjaxjTWGGfHpF5Fx5D/oOowJy6bwVFrzLWgMcBssffCy/TRn2y/SXIKqWg4AXTfxaxUplW3sA6
RDFmrkUDIMZiVgK7S44KaQcPqDpYTNuDLDltVbKlwqyJoNoiZTbc1QS+Od/GGoMDIwl9t9epF9FW
x/FwSw+SJd6kyJ8sEYa6EW1mk6khOqHwcfs42zGQUbtXBEtwBTNytIlu5/Wn7nme6iR3tQ65d/qe
3B3Xtc8veAqchPUa57XiB6tf9ld4A5tnQIH54fluMMAuNbnhpuY7+vu7CpboG7o57MA5xBMyseuc
kMUcEf4kPMbpiby3/rLUJOfNR4pYiQkzDHpUjKwNZL7Blvu3g3I5UJhE23994efBAp+Pu9wjKS6Q
+6+mCkHdfcNJiaK/yeiwoOj3rd6M6APG9g4+CwJJjnRZ9GPCIdDBKV6exUUsPLOCffslIevQlc3u
PvIeFfmBa9cTXE5l6gUbNKatn1rTBUPpLftiS9yvLGpst9tYY1zwezGJK0DB+OIoyVUXvhGqYRQa
Uz1LtfCKBHI63CSVVluqys8w9j5n6nXIYGhl2lYTFuEtDz3wF6FFH+LA4QDgzVks0+xeFI//Uf2T
XgkFCp3QIvwk2i9SzVw5uN5rCzsGBKJhQwUjhS+SQULX3f89pTIKhecDoM07avAEVt+bcwzbLFwf
SAob5DAC9u6Yjkk+Sh9h9DTmKYSWfi3SFGpbIhKKaAIVaNBGYX0SJZSkY4MJeNtiYFWXKaiRZgoT
en/rn/WUfpG2Wh3FpBjGbDzivdP63Zu+iS5NTqPU82lNLwBRJvdeShlXFSuFy2uv0VKImzBVTmTe
zRKe70UN38wXHiNB/48no5ERj4bn4jo4BMmf4CiNa4bRwyymSy6SbUF7FPwlgHY5o1fdoGRFDuLe
4ZgrmF2qByjFZLoYnn5fSJ47izXRF+hJ4RnmCIu6RWzV8iZd24WjgXgDHTZXrKIwstxhZBOXFFg7
CQorusYGoVg4PWSEnG12Yiotm4cfQISQBS7/m5EP6jp2ErJXQ9CZP4W3DbYN0K9si5AVrQEnLYjQ
kb8wC9eyEWZFHzaKjUx7NShQXW7/DtvjHEBoEKwNetbM8U4u4fuwrRUBZ68rskB5Scc6RuKqOtnM
j3laypKJMwaZeqtD9ca8yYkToYdtwROKzmcFLgVukXs86zrOEVIhb7BRNHfrvAKzVouGCUGkEjxN
v3tpV2AKsgsru38ZErX9UDNgSlKIOTov91Y7Xh96GpdnL/wqaymXwh0I2XVLUU9e4vtJs2nIgHee
C35AClzafcj4UnZ3yOkkY4klFiDcIHsPYGmZg9NaO1AVAOssSbZNXrw/e/Y+pilwf4VqRSLpLUsw
TOZQWUF3diZ6WCn7SRi7/GyNNR+K1GP0timSIu0FAFM2DSseTqhyTJ2FDIlnrBlLWtWcm3O1xHNf
ArbLlL94zsfApmsOOprQFNX6VEggRdB/6MbXDTadFXwbERP7d4Bpnwxo5fwFryL5WsnT1D+PPpkb
4IKCwDkIoMZ+Nh3mD9lWu+09rixXdpLXFKl8RGaesIaB4zhNCxbkBBHh6UnXlKFcfDEMqNnUxP+U
Iy3pBUZeKkdvi6P7v3WNsRRMT0xFBQ2mL0d4Pr4qgX4/iUUe7J2HAAv9h8T5/zjl3YTjpN8mpDr4
51bwXMNpLtz2y9wMnLWJMmelo0ljeTYD7lPs5TLgkwTCCSVH9q+/A7ljbMiqCWYR53dWJlkAIrCz
EfLYeF08AeyTiDPCySwqi924vrGxQKb3GHk8xdwSrIjylPQm35lbgAcRv05SwnjqjQcaageu9M/l
R2z3p0MlTgGeGEkQWTrm06GBG3T+TBDYsAM5ztsIz1ZgLG3XTSzalifZKwsVbu3GS5UC3xBgF+lQ
azi/wdWC/dkwxIgb7chkUPnH1IXylXhMbu09onaS0NPRT9glD+upO6TK0X0F/5tglcQoCRlEgcC1
4kCRQYLkSlAK5WWluU/INmxKtb8BTWvlA6IVKzI9m6k6vt0argo4od8KLbGu4C3ipVKOCQaFpwhh
p5TYptyNfBefft4Ug5txLNlK2zvhsgBbYQcyCtDRKGUIAsC1ZUXGJeLAiRHykb1sZtpk9b2AWK5L
Ejp8B/Wo4+DoInX/jrFxIiCYu6yl+6isKNbx0tV4BQYQXl6rzpadO+Wlg5k9wNCQUHxlE5LORUBE
2BV8j7HnSJuAZdroE9TV97HXMyBp95zcRWrCwXpXm7YonVY7+sxwek81CYudjOfgzVfZ9wp2Pq8b
640i12zuEbTOhv0Uw+p1k8BdCO/oI9+OuBMLkcaEkLyG+y8U/urn3gobVnOZyPbPhY2uyFE7gZP1
08NMzJCOfES8lSZsphVEsqt6zgDpPJOXZG6TQFWHibqCWGb3BZsiopiYCPm9GIAXoKCnhFvLPHGj
4j7yTWJIqsO+hH5CIbojJc8OqhU+wUuu21gLOCUO9iEwUbXoEOjYeKcfgI336Ad6ATohSUEu6v4v
xYXD1MpThu5pgYiWyVdgkVlkQIO/Gxn7ZsnSSZ5IoThi9jWewn9WKzAG8tFA7BoYtW1RzVNY64M9
i1HAUkKFOpWRVvUHd7XJpVV2Q0pHOgoSbvRqbeYz5qP0kR8QXTYWgxqCZi0slU/pUxZbtRQmlMKm
d1hYEKT0ysaC1N2DtfPRtZlFlRdY5NKpY1MjSFVC5GllIEVAXPhAfrw/dqrKC22mWhtJR/9qOk7l
oZD6K5sAKpZISs3GNO/roV0B1iP5TV04kTLIyaHWS4XxaoRb+IGyPiqDFGLEIWhNamy0Vb5KN08s
Qbt+/DX6ws4DjhGnM6FHvq+gRzpkVsYXHu4I4Jo/DNviJTbtnMb7wKAu5I1aEpTjDb15tN1DJufp
rT2I/uf7Sawl7GkOut6EyCXGtkLhDp+84wuK1h9YT/UtjTug8pUJfV8Moxtp/j6X2qtEuTw4vz60
h6WS85YirdfyNmf9s2MW7O0dvcYbQoyBToNTancLCtewiwpxEiuANqbLJL1vuHuWRQL/ml63nHBg
U2EOYVSK3dHizSrImSrLoizvr3W3OBiWHsj8UFa9i41VwBiYriwU9D5Dq0ZrdWb9PDPRJUySQvNG
9FPx67LiOP7FovFATr/lArxKUgMXoJ3IifiaIzKAmWNozqka9O8wc5/KMdQ6YyVn1JL6ICKVKZhh
snNovEArUwkjhD+d6rD/gKZ8AOKZCfB6AxVAKzzeAmsW/T6umA5y1tJpOVSkfu7fbKE8YPJ1lJRY
0qsyIq1b0FmUi1J+Jx//a7NTDTc1fE68Z12Sn1yJoFaZaZmb0fP68mZ1nQRzd6eyxDlJCUWd1VR/
3GTD/L09iwkvtu55Z9S6fD6/CUHcR/I9dNS32j8AhIPVRBPfn5DhO7tlpOj2UrGJhNHcN58kh2LQ
E5WJkeCBXsLsr2/Xs3ADojy34+BwrTvIBReLZuMyUHnCYq6ycsD+meIBE+uksV8D9VFIui/aoOcX
GJL7WRfKTBKJ0p1lvzyJOtrSKJ6TX7zvQTFTWUZJOwD/PNp0zDrxjwmz6wvsnOJpkJXMM6xzgE9k
EVxRGc/F7DUKZJ/x7CUIst49hdnMpkbzB6oWK7Z1iBEzjrr538ekkO4gsTcDDk0Mm1JnjU1A25xN
OmnE64NqAnSvx2bwi7q1NSufYpzkmG1DW7+LTkTVQGkwTv52CiXPz3XdHpL4zqyL5yaSb1KdZ3xp
SZBagBSb+sE0b2vqNJ4yCE33lRVqgD6FUBNOoymG7E6jUc5zijlTfXkDenV01NAH11ny18VFrqf7
ExuUMWcRgjp5gk2W2cAJlwMHCPj3jeUIriri/ukEn/S5UFDs1EZK11c91PCChEtIWc34759HJAdU
8d0PkgOxACOZbsJTg3aSnfZn3lJIbyRICNvyF+YfPFVuh8/uFDebP25Akalmrncyn4ldCogDqTyX
ShttjqrIAj1VC3Mvc0JQ0SVMQX1+7Qlt6/1zjBGH0GofY9Y/1BlzwsH88oTbRLprIWeOYsIxa67f
pTeUvElg2Psw2Xvzp+pOETdwW+mXvBmOJDYhh1lbpDbXuBOOcvzngdZV1+B/As4k/9A70bfdbq/J
CkEgWYmkQD0oxuFhvVRpbuGB7mwL1tMM3DysSMBM/Q1EMFdrc7UqDTrDDzNfV2bfVigKjX3S6W8J
ZVRsS4fB41DFfFQ0zGWY2yCMjTFEWWXfaBLOPBgGDR8O3XUdp7wCReiwkiyzFTwavDgUf5rOJtQ6
hw0RrT/ax2pdYgRLO/IRGgoBnxH0n3TjQOibLPIuCcgwcaraFYtlpFqELt0tbp4oFetvVkueTzSx
4J36bfaa9p6lNFhLtVGw9b8Gxp02aURfuFCLaVGGpwgr5/ZHMtO4uz7ZgC++m7EPLtO2JHiPxzxg
YFxaTgHZVrj7CnZQ21bk8l8/pbeYLoQLk9KR/9nQ8/3vJsrxdcIoIzjMBpxqz8T6x7SFDq9W73Je
wi1RaWeuIuShmREr6PruRXwwiccvLLsGfFFZPEfNXViDSPcoSPsIT8aumhHsJrlti7nKxAf84loY
FYnmG18rxiCtldhTgBWCb78NMPNIqBnn7VOqTmuACO29KjEHFTyMwseJUH11DqEx/GqYMdxLn/IS
o8ot6/Hjzy4TuhF5BQ/utHw7OD1PUgF6iDZmt6n7BB/V8yuzyN5B2OdQlQP7UtNbxiE2n92V5hmm
Yj/NWOzrMUaF1P7GAprpOR+hIKawnML/pIBz5Z9tWp+iB1JP/dFeITR+7ya0BEzIYnEQ6P8VMF4U
1oxkD4KHrLY07SgtYGg72d7lJyW+Xh1X80OPglCoN4/teF3EcjzQYk/cD6neRcD3G6t8q8Z93dIf
LjKOkWmrqpXANRoIEqkuzxQzsZ2KfPqJDR+dJGzyIZicYySzIn4kfslErwzkyHxVR1+GgB80mZ9R
utDWYuBFbzBxFXUg0bQ0XNQmjk12YrgF8rFfXXVm08tpbFU1QtXX1+9zTFU8kKAQVbc72fArjq+i
bfYsqpMY8cR96WU8tFM8tjqaG15vbWjUEjOwQi+UedxlTkqgzewc6GxVPgyLo10rxDpdfMyqz+Cm
sSDFK1/gVI5JAbl1xufBMMtJJS6nP08l6kpB+G6+Oc+iJ3zjsePysnXpnsaZ7UcRZNhl+ovDZGCZ
O9El3s/AZl9UHplVEwqI0lTQ1duv4AEQBEhqvODBuljsWZlI6b8F8Ewp4U0X5HCGPgzvi1magewQ
I9paJ8kI2HJmuHRJohhfDLfddHa7X9mSx/iRLUJPU+B8Jk2X5shhf37BKG/ZRbIqL3Isy05tzeFx
hHlyihmaFM2VBuvWbvvYQwGqnbA1slpaHHQmZ46IAILqwp1JqItXjt35efmGPktxyEcpDfweGy+A
IUhRf+/L4NquwA7fjzMbDWcsJBV7z90uM4KjN048llTI+i+rTpssV7zlWGpBy6A6RUtG9PJ8OseM
KXsD5qw7mdi6R4CzzfN7JjfQAHf7ibUxDMYzp43fYLWAh2kGnG75UBW5wW/ElOxVILIlQTYRfLfd
46Ez1KjcNIz2mo7X8gxk2vrnxMIL8tIkk9FneLZIJAjvGju374xfKHh5azuzP2diaT2bwVJ2LvMR
Vrz6QPen9U4aTt6W/khBwhETyQ8KSYExmWlhbfUiNFNXZxbwrwXdlQhR10DG2U6Zr5gfA+87o9/m
EjfZc4rKp7QSqBuGhv89rNu49sLD2yOrVjXhXycT02XI9Ck7CPFqxcF/EwKxoVLQj+lJSwlAMhFZ
qe1oEznGHU3prH5gNfXpHfnzu6oR0fgcFVLKmAvELpyB6qC8RfEBSI7yC6TB/9UQNf7IiP9+Afab
O8INDmMWGnnAOcqq2qbGkD1BhL4BlSORmRX4G9QbzVXxyg2VyYjPiPd5jpKL5oJ2Z3++njDb9nec
GPJAZFyaJE9ixSvB1B28z4g1KV04ZxkXnJq86VyQye3pXVEsGcQsq4TSx9Nkm2svo+zrX3BtDqpr
C8WuiYjV9cjrzYXJBytxg8dIQH7JEVssGXkNn/8I+zMySeM8kjcVaS7u+u4qDYdnTmbxiF30F8KT
wEtwrXAMz6lalPXmPr/zyIW0C4LKTgqV6X9Mc2IvLMjeOowf9h+QW42cuUyh6BtJqoVMCyYMH0MX
lQHhy4EyS4OiJAIYBGCzIy2QgeKbo+bTqq8TvBcKqUq5wg0uZ2t54ib+IgsrqwjYALVBAnMzUQ5z
GqUa7f0LQi55CQZbg2Dz6n9YxRfHKl1eSfjfr/BgAa9cXEqN7iptfdaobZJa16UGCU8o+/yUx7B3
20k9vGD08APp6cUg3YYgiq0nEX/ibXrcPTQw0mVomxFom2Qy3OX5kEOiWIhnnMwUGH/BASKS8gAw
bD15HDmiQEgDKfZK8IUbygnD2i4TvWo0dKC6mGwqi9MdjFC1uiMlevaQJXxWqey5SJbf6F9PBeUI
WiYN+IQNdIHBrbfrYrsKIJppEmQIXBhwpyQbb40fIbjhd1JGOnhcbF5fvDNOThlAIdnKxNWOOV2y
OMCfkYfa+ziT+LxTLmXSOIwgDuLZcECJsCdfvAw2lpa44bAiHWnc6imbmS1wbtUXUMyXpDPE4Z/p
ZXA1B32My/GpI+16XtNVkSyt67AnL11bEBnI0DsmJ4zQmDf/UD/1mpimmGAHOsXkKDXycdz8jbBq
u4d2EVybiYb4NcOhFJa6yOU5m3si47Wffeuy86qhWVQfcAe3DPqhGX2mpPUH27i1jHC3btcgizrV
Jrj1RmUow9HMIQYsbplZ/ArZmNeHBekgtPGfTDGCkUdWlcuCl8QBgFLfyE3dsdAzYPHsbZjC5aEU
12vS0tM52NraB2J5Qj2EgfoEMctftdRSlqVGYpfo24ktmXXEFT1jaBCFM5QCG6tH1w1K+FbzLFGv
rS8F5bXfNcFazn7ciyCipTgs4g4Fc52Cob0g8AihjgHLU4o0bAje0m3cxvGx2r1sZ8LUnQI+3V/O
7kf317DwxE93LnsfIkqIUq3dRLEeQYrhGBPg6+l2R5pcbW8hVtqNPRb1hUnmkNOUpYBx7+DNK3mc
DeyxGBI5GrAZL40aKFyOaxvkPey0RZSY7aYV6T7WzzxhsMVnOrfB9/2h+ZcVqjA4aOXR+ZQIBvjn
GsfRi7OQ+gIMtI7O7EaHuYMAu5EX80ZR8IM9Mg4XihbpWTVy/EJKW1axwFBSDFtJyTFRJCQUG3NF
TXWMPwhoYT+Lrj9XkVb87flMKku8Sc3uxQNgVhgj2rOaMkdt7Zkq6VvSFdBYkNBuZdP0+kqr6CpZ
vooUay1Vohzy/CfDWPGaDB2/S0MocSZHS2lZdj7tCu54g3zTveIyqL4AiRVVTntDufo1LbbGphdg
LNhcFCW6YTGLice70Awvg6LEHHifyV74e5kaC7g65JfuhXfWF1YE+3pdXANUUheM4OMMdXyDuXvy
gjbzIWw2eXBQ51bbGWutyug6Tqa7dKj2X8yRWuDaaq/eSvmYkKSxab7tw3SPGhQSZM5kOhjuJdLh
Lyu1Rusw/Wbi9FboAXkcuZaQ745emhCY1FsPNlp4YNIsSUtwSBpulKIa5wY7CwawnvSWV1jPxtCp
YSIRVBiX6EXBkcAd4aA8AT+c9prO7nDiLZaMPk0sGcTmn95UGI6JuI/3sJOEwjvlivprvWMiCHK0
/DZHtAJdMFU5OcQz02gf1nxhG2HxsT/OOezdI2nz3emnX98X/GC1+gzmSRkYD1xv0n9ToseRCAeH
uQPoiT4LXTeKCgcrZHAIU7TW/vmgy2h+fO57/pfVAsj5tYFDU0pBvyvo1phCJmOpr8gyBMNo+Nl2
1U/oit1dsUqZs00AZ2Y4Wo4O6Bv5BwSseyUalT75KfebqnVrFyMWWNiLnddgY1Bn+FUtaIjkEJKc
Hduao3jpmD85tDIYjLCwmcphbx7uhhj4KN5WGUBr9UqLlZrr0w2vaiv3579sbkl4mIA6gQ6a9Czy
9aB+izFH3gFhLcHHL2IVXNrLFNbHL+hz8kMlW/rA8DMnvKbfVLIzCDHOW3gBlKX6VpYkPrt5GQew
rxC5LPunLpNXRfrfnqhv09autcSGD04fMtZCGoKgMca7hNZrHqXMaYuDokxBHMOPvIwEmw7OLgq7
SRDxJpper4Gaql8YgLUZQMs0Q3uHJSzmkbYU7B8lFoWWi9zTWRyz/d4006e3OqHlbhErkZhhIszy
DU8pG97kCTei3SAzlGWCx4m4YRW3RE+E+w9rGhsZEGLULqio4Yk2xba++lwzTncY0hfUI4A3f2mi
2TkGRpgG+2LJH00Cqssb98aqneCkHgCyaero8PgRl/P7J6sMijy7by+obG7VRrYEjvGbqrTTCNfK
I07bzv2Gjt56Jo2XT5diZd7HWxKADKZFaz9ZLOzyKOl+JhFIPjHjjgEjZdRyUC1Vk9pLRqrsbJNV
JGdbkEeIUdzJ4Cc6TXXdv1GJgEGT3nrDQChbOvG7R/AetfoS/kMAc2273doccPr6HZMI0C0klr9J
eWB2veR966ovl1wMSfkEunSwYviAT2aHEe/IuXdJlsy6tGcrFEbz7uPX7/3wheHM6Vb+LJzWNAKL
db8cdZHHvHll+zPKK7Mod93UY34yhep9dZMUdQyK9RrQVwYbW4qVfkr5MV9YDsFGjlPc3eE1I5rL
WLJM7wrGwaSD5RiCwC/C3QfFoM7p8o6ND07fG6cesBUGtpR55WgrVlhewf8GFBrd9gD7aPOR135Q
fgR7n/AcEGaHk/i+2yNe+ojCiXPXY5ahhy4Dl6DmEMwpIglqLIS/gP4mBQI1olWIl7QsIvl35Tqa
7fwyIGQ7tyTQglreNcvYKk4L0yS3Zy+EfbSEozhzA5GaVlgyxcF93p/KyBgFRUmGdwlwwn5lV2Pc
hemLi2h1nUt0rUwutGFKd2n08dDaDbhHnRDeDUgHdDqER/DrHrXbHqUowgrJ/fEgeUIyAK3613jN
5ZWwWrmuK/Ws8qT8eX/Z4mjrwj5pr1/4s6QpUXvsETdDWxGAR2OBFKFXTEWinRiNKvAfLzKjcYuo
LQ/8Gnd83a9Zay7yNfkObtyRQ1wF1bxNFpSjYD231pKopZK1qkaNH03UyZlvUsiVFlYdtB8ZjN/v
D0DLRcNceQ1hXyNaoxO6SLDKPBuWlFMptTkEkb+Wf/RVWbV8EhUNHsoCtfCHiRLTAxdl/uaT0lWd
L9n5qlTt1QVTrYE5FC0wmdjXZnpxAUSoC8c8Muuogaor4mgWLqbjWJz8dRWxud4/Dw0XFrJFVUDz
+5fc70LTA8LaXuSdsQqnbq2hV5goKtPtUuB8UpBVpPlP1XVnaxfE7FRmqwM+vIMqkOC8D/QrOEAE
pxWI8SdaTXpsOLct89wMlkpZIM2OlO3jDhNb484QLeQ7MIZjM9B7dXNVuxHfxrGA7fx7PDDLfhfh
yv7rXylfZbUc+0CN5g0ckOOsBzfNkv5eV/5Bx+cJLkcw2F0gOF9lALngFYlKAfnfWHMP9uFrCDp0
G4Dyv/rDVlUbeswHv8IbTJzWIlB2bpfGp5B8bRW17Sw4OXVZYZPb/sUOeDU2OlxZrOAxTyl07EGZ
8GTZuxZM4r7wNjXrfA0ou1/by6tBYMQP9aorG2M2ZVpNoIBjQZEICh6SwV6Aw4nIyZnxtVeVxSdS
GLZujBd0l7FqdzsF4aSYuQ77Eht1A2Ao5NiX6tQGgmyh4CGGzi+CDdvKZi9ZOqc3z9HljmMldNgB
06YbxL3EwMC+Cgfs9xXStNLepDpAT3hhYeg0FVDiacMTm3KPdTHRCaIXt92ncsOGQH0Sx79Awq0V
sOYThzilrZrzidtUAapbkDr9GtNtEy5uZjG70GyMFK8xOf5wVpNur8ap33ooSXKeWZmqDhWt7hA1
2O/Nnd6KOki3oE5WoavaXvkT6kjGQ5+mekBbPy+WI6SyKWq/+SU69QzWR6/zJV+0Khx60Qau1aS2
r+ANhcteF4+uhBUyjuLOTuGbS/wIEBNyQb/Rko138nH7bzk0D9aSN07iUEIWg3moPiOuHublKU4y
R5b2MSAqS6Lb7dY735Ew8Bpx6zfVqdHSC9UAfNXcXCWsdq6TdQ0JyNHYqGXXLHZofubUXQc0dWj7
O4g3jrZt0Z2efUupaRxVNwXRSTL7dqQ/KRc2NHFW0cNnmfbZJdLpIz7RXTaESnEQAywMP+O6JTRJ
qdzwEJ7YGtC0CZmdA8qYhjRARNXSzALiMQ6JdpVSsXtM9H+llu80JDJCRxy4F7bF4fLhSqEtWZCN
utd/rGnYAHesdBJAed+gU/3V0ABHdSXFvEqxkvOI3Ifo0Dm5qeYomUql+9d/wCKAXAgKuZG4/Jwy
vlx/VyAmNUqMi70WEglsNA1AkyGa0pkx1kWDd8Vkv1SnpqJfUPW8L983g3n33ZDgkkKcOhdzPKcf
D1a27YKk/D1LVort/cD+s/Msq9YOjsTZJEdy/3EfiCuiY0o0vxSsRavUYhCmAWvDc8F6wTEh1dor
WXiPCiFDCf7O+PTo868KVIftYs0ryYrgm9+qCLd4TaE9HoWOeTbjtj5cFsSa9Gz93W1TrW4AL8li
eipqNokUhXABkV6FzSZ0UW/tQmEIOp4bRWN38uNAX9o/takSR3IygQclt99+XLpmMkO1aolbVd/4
96ejXJv04ncbI1ZlJUlWirOVTymBM8UK62TP7BZirVS81gOu0bjTSI+GIuymcFm3wvkD3rAuIBQT
GRXd8FYau022Gfs7e0aDGMCWxvK0hxt7N1xc5zyqqk7Rx154NhqhSsk1UTaBbGhqskuFzFZzgrdh
Cd/lgYML7azKbgCEv2jbDMWl09gQR+UaTvONu2ny4EQRZEKt21IO6bJj670PNmCLz0bi+s4g4Foa
PCPiMkxewyDygL4Vw6vOnVlfPfV6JAuPkUOgBX3GFa7E34JTR9LYMr3t/RAyRgBZJuHuFHHc9xpa
582e7N2UGZYSHKkMcbm60iVMLD9S8Be1RCCccDucqKjBUG2dhbssZn0KVjGjEbdwK1V5t7D+sNzm
1IdLuXfssmecbQmYaQBEwENgye2qW/kzCmHSjOxasZJmG1Cbwcf5g8Jpom5QxddVdYf5aQ5HoWGM
bndOjovfnO2f6Qj82YVc+7cxZSZm2PIjmUMlzBiQ6Wpx7WcqRxroQMHelPaBlKJha8ubFuuiWT37
7uvx8oBieblX+wzg36pyF2UG/zgjTStFlNpHd+yAB6a1bfbpa8AfGQyMDUBw0oYxsI+S5TSdYN0B
VI6lEPazcVz602EQf8S548hGe+sgFY9QSgiMH0iJyGoSuV3ObV/EAGH6wmh5P5pyYNENWXgR9yME
N1JAMU3bT5GuNebfAar3XcfpPBAMC/PlQm1oKQQd7nizsq/qoIhoITxusVPoNnOwC+OKhKqxrbG3
6VlNTd50YD3yxZlXkmO8YRvr+0+ECVBGKyds9b+Fe+MY8kgavS/YzPU7FmbWjOcYwvO/T/eCO/uw
oE8GFLH2EGh7G4KWSsuee41TBsnPFTPTH11ERMkCQP2ewx3orluRWXH1DAoIJgWK5mhDWj9NSYwq
9ObJY3VaJmjmUibvPwn3NHe9km+HQ3gtyOnfC0N5Ig/GrUjqzbY865kKfmCIra5UcU5RrwQJuCK3
JnxloZZxbzmas/+aFHrWP8L6zhnJxe04kcc5fUTuOdysTO76GKkEA+zN0qU6rfNJInprPHMSG08y
dTS6UUIXushguoXBQ4XXSk9DE3hqrVkdIzOh9B6fae2Ei0QGmJHmJ9QRRIdSMytZIjbMuOLsLp4+
/X0VvoviUP6FXR4zkdKf6QTWkT3rV2aws0c4mB1J3RqWDv0NmlHFRewoRQZTnFhVmEbs2A4uJUGF
VQJQADgLPtUlzgV507ICv/aPRKxudU2XL0EkD8TSLvOcdVWvVXQSPGPIHos+iWIyhHTO60Y7Ks7L
GFiQUc+3n1vqe7d3OmzYAa60q8W+Cs/SHp6euKaEJJ22hiIOMxmGFj/JuZqegglnpIKdEPnQyLFz
5n2HCArBdkqdVW+tQk0vaSkFHMjbprChhSjVFGSu21amoUfFT6eZBcSfmSbVTGCZloEL7S1jg5Uk
vKx3K6mdIXxPYMgdSpFYbkQCn/wofBbh1zlYeDaJO++S53TTsd6o+2F2t4DPTTp3Yw0VsvbJS2Fc
G68HWm/2Sb4+Bh0G3NfDWIvNRjIzhhVubNGVIRjbRtWxqjmvhh4RTp0K7m9AlnU1X86IQnEOjgq1
algg17s0DsVVRtSwGHj79xdZJVckQzYDOI1njRV4Mu38C2tdNhMMLp3hnoQstZ77ESNMrQEjjxwV
z/Amu2ou0DLE33GR7x3xk11BdQs4omo5w7lF5MTrPPas7UXtl7QGGBSQ2QoL69DlnP6FkTt547pa
IvyQ17ekJWVTOsHusalW8HK+J4SbWfqGBqMjuoEy0CBOushYTR+DLOS7tXwCgY9Oe1iCr2IPxfQc
Fua4jsqBrivH7l4xytXEAWvvu3/unzpFlKJyoJfeMCnHHwOwVspQX2MQLQmoKKrpvgwdb3M78uwO
1RJzFmTWrQPB3LBXxLlP53WXa3DLYUSzDQ2bR8o7VoEcmMZ4c2iiPccjgsXbku4XUYG2+7rMEuwC
6wZ3Ge3xN8qq8s1lNj7HzyUDOyxObZBwj3P3bgJ7z1lrk6yttodFp7S9dwjqls604L1b5b6bAHZD
xwzZcupN1nHNLg68XU4bh23SQDAcHmqaKycS2LgSIysqmNhO+KCYk5XkK1r2O1imu7iCT2Sv2y47
QGR69QZaQAPJkmelNSRgGnAu5ViYJ/7Jk45m1ASK+WGbYHBbqKohp1Ekr8QHMYfuQYAy3YQyLQC3
5Bq9N6S8DqJoxbrC3ZtTLEI//lluxEqGuk9hNiP/3BP3hdXdEi3u/drJ8yewkILL/ic8vx/iVef8
VlskVGSk3aje6zp+F0arOupBuUgUTrVB69nx68doE7VBKiC0X0Wh95/8bkkPqSt1nuLeqqpZTWn9
PPAL6ohEHD65FIDNFzP5VhYnDR9ES67AXIyVvJVl6m6pqhMn4rqhHyhs1gTMTF7u88xV5XZbxx0O
mEt8lq+WpwHb0wu5gOzj6zIgytkRa7QeQMXSOOXir3jC3amb74MkorcMzspf+LiGiB5CCSRl+BK4
Tq8xbkIbAisx+BNESeq4nripTcTflm7l0NqGTwqPMnsqklB3KR/eZZ2M3yeLyYYqB7hKC/JreIZ6
lGagOyCOvqpj5USvNxWkB5h2hFWT9p8HBaCY6+ASsfwljDK/dGYkNMyDwJtDBOIN8VTil6Oy0JaB
nhG+wUcEoYSxe9Cjx0Dj2yxxI5TZXmyrUjCqP63CwnVg4dgN+Mz622q8qAV47jH5UUQgOnmakTil
4YRMiwZJGDu6czgkFoi5Us1K+cCoQ2jCnL6FiGUXhYjDQXLibXkIRL6+Wpl8/hdD+RzALZsLP1V1
7LxtbRCI4YuqkJbyLz9z9ULsCsME5H18JbLgs8PcTvwQX4Sg9FEaQ1+stglezXRu34W+tbbVASkf
DTG4dNafVpYsXqw3Z+WeTz0U9wJOWO/pmkwKXiBbCCjgECIPljj+YR1UiK8zdX/SpqHjDCbgQWM3
oCHV26rk3e5iQ35nPomcfS7ZcvxAuczO2iZwCk9+VgwHyvfVVu8wv8QhO/7rIYFNk5BN7tsw+DfP
hzbRCZXeeE5IKAcdT5ryFKZXFf9HC1+Uyb7HU5vBfIInhDao+N5qTUNLl2DCpZ8jWhwhR8uqewov
5XFXYYZCmNSD/wIW+dXw8DgHzbB3Vo1zdggCz9mGkjtP/kJIoVemcQRTagmIVYu02jwkHne8t1Eb
Qvf+GZrsDzseRGWCiiX2U/4Rcghq8oYJhl+BTrUQ2Yl6h39V8jIlX04ToAcu2JrvwEuUbdEUfiHR
wnG3hQKtzy/JIYEaUYm3km4o1caKsu9modFR0dkrlnPd0Fv/dm3Vun0oCdf1IIi08r1L3ty7T4C3
Zhyu5TvcWWpcHYu40Ynj96KRZNtpXNa1lnBBCZjXscL947gi168ETKW5Wybl5bG1ANDlURj0LUCY
0+TfK+nWUHgkq+4xs2fnMwxw201K5XhwM0jFsdAR3QNYPzflzKab3OXyNHJ5KaHydIKhQsL1uGE4
5Abl4eA+8NpZ7WF126nZLfAChxED0q4qvPkOpmlBrbWqTCBiUPqD8J7NK2KlInvuw3gf6EcRwsd0
sRX4xL+kfOmqrsu435VwIquikNaMMEjaZbuhCogRvOmRIE0IsSynXzxBiGD/Y/NYh8En5V53eqGn
wOu7Vk/h1pLD8sMwNV9+E0NYDnmJ8IQavZsWDIv9ddLUP2AYpkELk1EO6Kdr2FCN+HneMCvAfVbt
PII4dUbYEhdlYOvphkhDltshbHFhjsP/V8hkR+KKiQxM/w8o8gSURSAaMBFw2qbAmuwmA6xu0JIz
6xAUFKaYQp2OhukLr/CYGiYHyZl2334htpNWyZVAlYydQUsmhRtXB2m/ACp7JnfPNHvM3nH7OZ2M
Y7EGV960qIZdzfRvkcIk8gSZiszaBJCf9BCTmIfx8SEoPj/XeNagqVY3RZLYlD4wyg/8bYBj0o0Z
c2NA4s0PJ+eNbQ+jlY6rHn6jZVNsCpoPRkGWH2Rb7jcDAy/YTJcxUhM5+//PCCnS3DpHiG0t6Ie/
6U9vkWFPCbwGRA1HlzwXYnx3UfdC2MK9nOAOBguPzZpFRnpJkxWbT45sj7X9D/6/ilOZegzgK9SP
SViUemKcE502QXyF0jrQtc9BUpOnvuI4NTVZvADLmTbGa+6PcPXklcH1qMo3QQXQtSvrhmFYmrke
hTZPE50BfEbj8JKzckxyyH+9kUjPmpDwuwRTHHd1i5LRQb4IVKRncgcAFLJBVpBG/FonwSIler8G
3bEzB7+CIOH7mAdAH8DE8MYqLbOiCXxBtM+qKlAMudHRJeUFEEA0y2WwQEjZU7X2wCjLX3IYI4dk
aegNFD2EK/Zv/g6cudvgvDeI7XNDwOqFfLQ/pDZ3mC0s4E94BH3xQBQXxUCzCVCd28OX5p02zD7d
49rhucDQ6RvO/LR/IR4e4sPlq8A0O2kxeh5PeLA+H7O2ITnlNq1odg3yg7/p5Cjx+UhUsD5p9cqk
mIwrhqPG6+AL5cjgplh5LMUcoomTcQY4NsguNoMJ4y6oI1pjIT7av1W/hZ40vJ5RiIc5HYCN0t+R
Xze4RWryDl0jvZIdovHznYoZGEvGXP3Ru03vZK2W2wl5tK1JuajY0cdnSJ5K9HYzOCgOzeuxdA9Z
veN4HPpJWvf3q36inLAJnodUcRSbU+h5CCuOqBotxnqhZNDo6wIyqYsqLrp73PYWyz4ui6pOmuFn
PmtRjgWgOqVvmDi+zH4g8ULB7AegIkPr7Mof6t8omU7iUq3SmJXWBL9oU+413fkvggOpu5nEgGhp
nKdhKd8gojzf/Fy/t/bdG17lLhi5c3qn0vrFuD13u20fujMX1FWNJR+W/7yKn1qnaoNDVDEl1YRt
SBvWANsHfHPYWP+tBo7d46LUvcIiR5q+sLKabqUYGT+nDUzLth/lRKcK2baJjfSXCpoStkdTbsdf
W+Uzx60VRo1b0Xb3hjAI99c7hr2Lvxaxmb/3eH6OTU/Dj1Lt+CELwMnjeTZFEx3UA6MEYelaldZI
ZSPfPw5YrwYoTwUHv1lghgbdRrsN6afAMSlJ4sDxRrTtIPtFoPgVWaTLhz9e0Ps/t+ILjZqHMNOy
UYDFZs6bBqLGQdR//gUA/OMWbvY0L3XIDgBeiqbMk58SFQ4ziTbbYo7QYwp24p0OGxpR4bia/1nQ
gNQ77JdiNQujWH54acbsCGB+xiM/rKatikBdhcR2R+0p7/IHTwLn78kmmb+rqa8VQnqA/SbToYxX
54E9K48457g4/HY0tDuVOljRJuRXSk3bQ0radobD77hG0X93E3klXL0Y6JFWKvtYN7o+chIZI1q8
7KFN5jzi0V1C4bPSItpiWNfCoWzw3VOKe9UVc0YSdLnZEHjiorTFjTVOkxq4pVDSdH/7PAsmSXm9
snYbb7wcZY5yHPB58GHA0umkh83vQgnIK1nLsq2jA5ELVSt1pb4WN9fjY113IHuqx9WAakTHH1B8
QLYuCxAMnBI3hWwLHEA+UkuUyJlwdwKSLIEPG4dYvhw3ce+yBW60bec5EqKgZApjmmNGhFB4BvKF
Bx9Z70Ya+6TWc8RhXyb0Sel2KKG/McCybTUr8GNkjlvnNvQNVElHfs/nAH2/IMtuTbSmD+ClXppO
LTSm4K9haL6WOLoTatzenSDMSaqFos2wYUJer2rfEETYnDNXQaz80Hv/GVYk7ITA4GXlIXLB5rNy
Tysd4m7OI7nzQdl1weisZoR53rDy9c+AQzlQn+aFPimlfqEDQbjEho1N2tQHJry4uDEkxoEHb+lO
6k4yDMNpGIo1XE9w6ETs+RvG6cgFqgSgPnfMnh4Oydsz8PT6f81xHqJBBJb0yxOIrVF0Iz8PCRRM
HADwHFFnQtwPTMKH8mSJ06KEEfufTenlQ8mLNd3IPuxmNU/O+7GfNZ317drVTC6QM8mB1lyRZVyj
XSzt5PYjJlaXjibBOGdjht8OC0s4Oeev1uIWuDaTLKFZS+x2Tf/wNIB0/+mvFqhA3PgcuOSW0Ubs
Bdb6KXftGRvX/+0yuHaYT7rRR5lnwaeV3nBhnBHgtUwUzVnpFBYZJuUAWDZkAbb2/p0UPbAGytn8
zyUt5j3+Y8tyInNemrlZX25C/RCV9lEP+Xd5Bj2CtbuF9Nx4l1WsMUI2AbaUHhqYCcquocCMkALS
vu3w2cfT5c5s2qQtE+wOYNlhsyozEBvIZTqGtslnAanZyijkNEvlSbh0QcMIl/WILo7VweR/0+di
X6gQIonWr+4Eh85kWLjxb2OqSi/Y9JUqBX48StOGlBK10tQC4CnyumxEu1aI+6/7+jthVpQirp5n
IyQ90wUo03lcZtfUcxreEChJLyDjLpOlh5k3GlCeRoyq+IjB1AbQiRLSwzTKqsVoPnKKE6Bxe+Oo
m6OLygW0jgOT/jJSoC198gIPbGeu9matxMjiQ9/5w4+JnxRdXUDdRz9Is0B+gFkJvRYD1pgGnt1i
2MovXDxsoMlGjhzNo00K7P0AKkLe4kDVGacd1XsAGBaMCfO4wMVgtVUkjAIOe4hnf+6mlSMLIaCJ
u8Sqzgr9c/alYCPU1Otz1FTn1a6UUFHLU2lKHTtYAzziV5BzqbR6YyRJ027D7tWNes+NbPa/n3hm
Pn0ImkPE3JxCuMXjGzcDOitUIWHjXtn1z1oXu6IvqprIjARa/+7XsaQ0LPTEE5yAR5JpwscKMffB
DlHUNgIvMdWrhqJXRTDakS57TTXt/shsk8nEvKDyZY3+PxBwj91Ac87pYxVAAFziQyqCsmNvAo0Q
NeOWVspX/NCd4ble1JnlqXwJ7sfHyamkAlMXLh3f0Ut8pddwhkBIqJhuz3mcDSKdEVwfHUTNkpaF
PhF6qji/N1O5RloDV04i20aL6xiGFhWV6JhXe4IqbO398/fPvVp6Y9lgZ9Ifp/6xaQMvqoVDjzwz
qfx8UPwtXMx1KzmgyVxDd7iol7KmVntVNIlfZcR7VTMAlhby6tqn4p92r+F1MebxsYuGUIr97+r2
wKdyQoLlerCxsXLjSfy+KA2DqjTXkGa6EzxuPeDSOpYW81iiyq9Y3lvsYFFDVoeBAqGkHSLoTYGW
daDfbV6xN4XXnxIE1KyRYAEckXgGFaSYPkQsEJ4o6OQaZ+87ZmfqdLg9pLTxaC+0BRmkUOAc6eDH
OkUR1foxcfbOJc6OWpAsZUuVEfYkvFYFPa9y6NXYN3/jzHhu4XHeKyh4mgPCjRsEyfXHKyXOz1mk
T1cp2zy0sSkCkfHJK0h0EHNKbRXlSQk4CtwHn7fCc/dTT02vpDZjkoxlzQQ7IQhCZuc4pe1/j45L
GlPAMplgJU5N2m1b0aMHw9bjgEpLhW5g0e4Iq0FsFYmddaA4SzZibQdRl+3JG03FFl3d1jdNTJSp
Y8ODCJMkjmk8+U+KHVvPJ8Owa5LRKrJ9/XkIgRyVmaJuQEL0xRdi8b3DN/Dvswg5Wkng+0g9uxu8
FxaRRZhFV1D6KfUjS5z1vUxcDQqmyxVPOEGzQJdac8JjKs6N7bIE/Ffw+SoXFnoZE3we/y+NEEM8
MkDNm0j+Jv4qEkv2TAFlyCQCWWXQ/osti+zWlVOAi1dj9l59a16lXr78SrBpKAGkHy0nhm12VZQ9
2b+pqxYcINIWr2WbWHO9hj5cK9A+bEmGKxvKGBLBApl2ac8+9glvsBElpyfwAsa1UOScdWH5IUmx
30Npx3yO00co2e0cA6PmIxAOi2n/9ML9RCAr2jNvI86dAbYtfumMhyEby1ShOUyBZMBmC8UsIPGf
3HWKOyp2OjZ1o0srzclnx41c7RH68lkfuDaMt1jhekOPimFZvBLgHBSyMCZS0RZbCb9EBHfKla76
x4FV8ybwAKCwVglI0OyY0JqsMknRfxoueJ+jgPGBGuahWxKaE+DuTJjyIMEdc10rAAuru95j21x/
ASFAIjuhKTaxr1YIHQGttsje/Xna3LLsJE1hcW4cvWHPG+irztT3tPPjNTXMR/9m50230vOVtHmL
jlsayAQNQhi9G5+D3n9lDio/8JE0ECp+shxQrYfu5au1s0D9QXibxoj+z7D+zzHn6sPBgldH+ND8
zESoJNTOrbKsIUVokWxJIo5sUpvf0zh9vEY1yiHj0oQCsoay6tV1f+In7jbZJvU+5F54eiRRv1P+
Dp/JaNvsVwE2dUHrn6gIPgwyowr3rSttrALTJTwlthL3VjTniFfk0HOHvz8UrcE5WarbVfxRUfoy
GTILMZYouPwcGPGFkpII+Od7M7JfEwNf9r6Dt0qcFDLpW/zADrkFcC1lvSFKVOXR6Q8PXaL9+Tzw
PdxBDJ9DM3qc+jQcj0m4YILowuPABgIgmD1ecFrBqw2f4UnsdCbpBKWi9yRHuwCyMlH1TvLRYnLT
6ZVf9PzdrqeOCOfWbKysTICta+h4tGX4l4C704nDCyzyaVQYIUJRm1AR2phG/BvmKoUUS6gdW6QE
ertzf9uhpcgJVgrUJDSJN0yEbxBEBDFvYgnsORPhA4T3w+be18QhqtXu0soocX69nyiD5VovKOPJ
wGL04PRsG8keoPAH2W9fse9ibfKrOg2aBtrMH0I9NReye7qr9o6fbKep7OGX8tfdSmoGfl1rO1IK
eNpH+O5ZYZHvFi9LFn+5IKpoSSYyOrRaUcS7VWksJuKkiAziuwpenQ1drN2SkpSe8mHgNWCphOgO
Bp2NLrS9OQKeWOhu0V5BqpnInooMqrJxCokp6h/mJ8x0mkR4uBgJ088hdLkM0e7D96neOmoA7cjy
F7QOqkEfc+RCBb9RqTmeDVKBV2sZtJG9q8q8tWE6Tl2xeF+58Eym9b7CWeSpdulYJR7/pYI0bNAc
5RZUX+ItC4X3NAaLl/GF8F7oS3RuZLM0HOgEdWmz6WsC+EIPFJRkqEpPBuDtCelm13jAQgXt9DAo
F9LZk+10mqbt9pzrc5R0C15goGUzWTZmDWAKq1FQu8BT/ACXhA1ZgfQcxe3DZscwVI0YzNbGd9z2
IuMDKCltBh72b00LBpjW1NDRAcVVoMz7G3SCYkO60dQi2zhLtvliUhBAG1IywGPHjFG+WDjhuW0z
g8XF03pygWG3aLA8GlJxdUuIdtsVWMMLiLM1PCezOBzex+WXcxpjWtYlbSYd1rzrcJ4YvSiOnU/t
I3u/XrZ+U+BJp7Q+q+krjjBNkhW9vCRIwGH6P1/JKO+do296VY4TkcWzswMJwc/4yoGxSZi8QyMj
y1403DC4RjzQmb8sVSJ0mZ9CKpVeC9qPayfVKcXdWGsoJlVnEBp1f4FYb2PV3YyocJ0O/ZsILa8S
h7cjqqizV7qGqpCsAeo23Hoe0hjZ2mRaFqVo2lbVWrtR4o6TbMY5WFqXDT3omEGftRKXpnf1AFs8
Xz1g1YtAHkFjx3hO1IV73SX3x11+CLgs8o+EWpUBSvLHlT1G51v/F8IGGcJqx6oY/dl2fYJ+U59G
LqyfQDbv1xekPHp6N+VtpVzit9aFLCyN+246B9g+ZzO4CTCoTZhsbIarwN3ecwnZ3fjbnA/GCSVo
hXMpe4/QXB0IeK1n7F1lo1TWcPBp19b5PL2fA6bjgUDdOuMCdImOzLvP1FBh9wT0KAtThcTpP5RQ
Ykh/QvHdo4Pr83zGnQ0QCuNElsZR3PC2gjOnlSMOfyZpPbNLttRG/LQprtsOIZ0qowikGaaBSlRM
TAWdExJ8tX6aldkJrs0Bu2/cBbuQI+nkESybOz95lKM14I2YnH7V11nIs60/CuAl/aMdhxs6YYvu
zGGu0OSEWyM+GCMEXnZoZL1oB2qfTS4W9KV0QIIf7a2bw5fKtQh+c6nwt5nIadC0ugwVKRDjYISA
2JMbeFdT4+xJWWJbu8qrRBEFQNgCWV6dLQqudVQ/+zYAfYQ+WQm30Hz/vnpO3E11pqNhH0dCWZPq
9bgyqZqd6rdLQcDZFUBAft4JcWrHrkxqPhJp+Uq2+9KF3QSvlIDi2brpuZdXFeNikOgzMQ/dj8mS
1hz5vXiRaTmIIKI2m1Y6ristnV4zjqUurAoQNna1LrCud2tXgB01hIHHyXplzgBVyoT4ABfrdH/g
H+EOZ10hpfSmThuga1k0wBCzZHGWqf1XJJTbGf3twSPNrCJUKn/wjJLqkwDSJ4+kyKX26/K2viIA
P70XqCdiLNwrrvC7ubmJh4OKSJpBCqdjzXvj/WfOrjgEqrxaPg+Ap7KQtytodsIx+zW40HzF+MnJ
WMcfx8aVHD0bfW9PobpeOEmswndM1ps8NJepjcC3QZpv/21MT7/eliZ4Cw6gonus77jWTTJR7We0
d2xZCqy3KU48jfGYtTzhdewkANxwW5fSba7EYxWCxJSmFMhRrNO8nFzLvc7dOE4Nqu2hEHtTTJDK
1/eeFXNSYhLjTr8qH/UxQbYqgPb0eg3YBp2aY/fa3/Z31G3HOuy6njHSkkdALq4u8BE6hgSJmIga
xJd77p2eoGbP1xo/TWH+mHhP87jbayVyeTuylVN/omos8Ho/CGTtz3XWr5sGiMrBUzlDbdakp5yT
HT8rRKhqYOheLnRDwCu2KYb39xs4be61EwwUp0DFLo9SplxURHsiHJFT7WBdu3c3wYTLxKKtNlsn
2qmq4hYMGAjsrBgK5FS4QZXmex610xvAG2Put/CdHZVlWqHvugYRooYXE/1Pnit2SviQyYwZui3r
NCwJF5jE5XXqf5vzYCsNHqOF+GEe0WXw8DbUwKzpT5gj7AerfHtT7BLfb7KOfttCkNft4nhvjN3t
mnT9F7fmGYWv2khWNzLHU1NKu1FVtJtG0zwfxFORNic0PGOVmWvJLb05ELfhsSrga+WXTFWAPaUh
MScnGH83LRUkgiphdbdjYBU7S7JZWd8xncHEeLZVH1EDvAQCm7UNoXhHs7dlUMcs07aQomZ2pvNM
wF6s22V3L68b26FN8g23ZEjcVHN9pJnwDQz9plV37bHnNm6ZO/DbYBShI3pXDjj4s+J/J/4R/Bkz
rS7+MikjuTbNM3mqFCihvJTWEYPHRaSpgY2NT2sQSKc+sxtXOWe/73dK6ocubTY8URsFiGT7+GMQ
23+oLF3Eumrr9KT61Xm5vKsTSnWGbTU8/VlNLmZ2Elew3vYRw09J1X8EislQNUvl1KANZtgSatch
8vwC6q5R3DJFj+TeiezhYzA9EuW3OGkY6Zi57nTTOvgxwCDjHe3ww8e1ckyl7bZw6a5v8gE+qgA4
QkXKZXtLqQB/Ji6Se29ZvfZZ1p7VhfYcmDP9qOeFXiDpyiSdknb75so6WGmP2KCcT0Dq9dDwthLA
mqxffuN73Iut3pupbmHJPlbHtZUuXQuPBYTveeMgZvHS1pnS0K5yim0iEws+lVkkWMM9b70nfm2p
Xxzh/WHgyAihw5MI7q2p1H9620LhULYdlLM4xrN5ELnOV1mDGbaBV/0U+6prLcuF9XUxolyHdp4d
jFTAMfmwGwsxGBCGmXhQvpm8wShOPOtp2L/uQsassIBSA6Q6fK9jEIS5m1D9DBdx5tOLJiQsXMPu
ZU2VWAOizVJXsU8Dy7Gwq3GHFXYVddpNGutlliKuiPv5WktshSeCGeM1xraw6slZHJ2EJSTs6z8E
hQMtW4ajuWJWqxeR+QSo4Zv3trTnm01NFgi5Klt9CimEyvW90+BOsaDbUgDUKRibtqnmxyPBc1Re
JZO2UE8eO/SKMpcUuxkEJg/KttTNgIS/LW21YiMrxQP3rKC3o8oxyd4TdFKDFM8GcSkRGGmtBKhB
/JTfKWPY1BBRzZSHI2Eoh/uWdA/DGxiWCcqhhv3ZTWxvDXSGv6cVN4QP6uE8sTIIr+SOYA7iG1QA
uWQprV04F1Fgr+PTeV1Q5uVzb7mQynmZn2IK3pVOZuIFwWRKmAIMtWLA5J6/Rt9fPGz0AU3eddIq
LVjLolPV1iNZt+q1yzWtwRjw0GHi4QxiFcBN3T+QYg/zuqydYwEPhAb9YGhU98O2CLmEV77FC667
8JAoysN46/etVONdlPu8XMvjQcprVswWkTJT0fFwHxdSp7fDwwkkdXQk7IuFNwiBuEgkdErNPcCH
Qu/nz3DDsuboT/FIi/h9XJ4jshbwEs2gj65MF/cd/KPrfhTQ29+o7xdcdRk6XGxiFo5RY9A8M8qx
de2+7SBSfUgvKvreWva7E6eTnGLLtMrj7vjYPxV3uOjaAlSp7BQNav6hQLzzJ7bxggzxVvboW2zv
Lj+s2B891dEOQckqVCFi04jJhPq94dsGzrTtp2H7u9iFS66AkC6TB3r0A11xBjrV5qbXkBKuqu9R
i2MOiN2I9mPQqUmGFnkQGiSm0OXd5TWcpu2RqtzdJcyhYI+G8NyhKz6e3MKjkPsd12WrZuGHz9h7
erpuy7mn8V3sLJMDUrZXOdtOxaDyXWeg9FXRbctcC3XR7G+qbyGkNHZI5JOayx4LLpH38e1ZZolc
cEHBnlsn/781XBi7MAkQycymiXsa1E/CXAW8KrsoWOog2uWI6vYU/mBByLJYKNpQOSkk5/FjhTWm
8KC5l8eO+pEpZSWbdT2mRyGUKWS6l/R5XPc1ZhFL926QDC36oY41XwkBKQw9TPjqfSobMuuKAQ7A
/HJgEwT2WarBpk1+byRHLEP4DCBniT/YEVKB6oRT62M86oLomZXllco9qMHUGiVi4NfRTet7Z4py
Xg+T3GW/U3iPIG8vSrIVtJylHqT1e5AkYyPv0wQz+bKpQuNG2Wgg7qqCiE52G8j91a+mKVRxonHU
JBtE4gp7Hwh+0HTVlKnpoOnBQcBgBkmrq50pcmCt78zy4GZZZ29mp77ic45rdo3Gz202E+Q79fgC
15KC8NfubKkDeZI1Lc/FtyyMiZUcOmSe5YwneQwxxiN6I55WOwGAHNji83u9i8rCtBCexwxOsJcT
NOfORnv8mU7s6bFPjdRn5Tze2ZV5ejhNRUIy43wxxYR7f7WyPA6oXs3xg/j1UsKzYZI7vvCslZ1C
AKs62dmVJMQgZkBNCGPvFKYr+T8JXkTx4ECu82m2Ce1bs7/YKYd+YLm+yFxYpfAH1RA++hr4Irwj
OlAlyvYJsoBoegO7PWZUeXkM9zXzAIOYlA+ueIhOkwol8gqh07As0cRuLdvDlQqZDNh9EXrtdbFO
nuaAwJux5/9cuPhvu1R/Ec+SJjrK1KnqD+HwPnPG2Bq6x5D2ZWXtMaRfj0nZ9e58Y+fqMmMP8XpM
o11Zkum/phK/yB+Y0jaEHz6qFWA46LVp3CwaGRfdhgx0HWFMDmWuveo9fy4nki9BCwdbfX4OARyK
SPTThn5Qq4yKyKGD+4F9rNBOYOzCbexgykQ5Dcffk7fDU+XJI7xuSgk/OHE9tgKtFgg7gP4zKMLC
2lY7uxtykdjqYC7iTjqvFope3dH1HvolCgzwkLgF3Bxt2qaG7Md3n65ocNbk3Ogsa1yMZSPZX47t
xu7ICrAnAz0rcuYnpxv0x/NtGgVrct6WMjbxHSDR00B716J9ehHxART8Ru+8qxRA2x534WUuZsEd
zwj9jJFfH/Fax0XxJWXWjlBTxwF2tLK8WSl/Jut2fA2NwUgQpTaE9F+ajni5KToSR5sHkuK8OxXd
iMomp10HgwVqbQnE61v7K39RBtJgpsh+7eFARKxq/GwspHPkyvbZgwnJVBMgbq37eyiyk6/T6oLi
xKsoH70VN3LQr9/m19dwmPXCe1WFwyIB2p5+b5ewSgwlCK4Q+RLhnAj23/x5EvSRNzYR5w6fSCka
5RFpqcsR4gBzxZkmEcIqkdhI398QDGuIzTZnrHaiPhC/HQeDLtFQOILs6aPXo5ZbjWYlIk/xn0wm
mY8HhC9ewa8RX3oNbcON4IoH5Knej1yNA0Ur4wixHPnkX+rYnPouL4Fhq+N++mIYMaYKPJvOokxB
alLkb9KRVzdDIO6b6hPMp69CTtuyoA3NqoSrK8z8D9un2wTmBiF4tTKZdIe4Ku1qq1HLNRFMSrUF
/OUTyvbJOBEjPr3Kc8Hv5pOK9a/9o568fXUR6GpQyIuY3XRWe7ncisq92EmvRzA8Lvc3R/Lc4NUd
8yiYZw0kaxKEo3rMQkW2nK9JgevnGIkrcLtsyWU2cx5QDjzYhJYenjS7z/sysovcpenVH+iiAp6x
gxTVzEWyVDAPVR7OcujXj3QeZPhr0K2IYr2x9spm5dLRdpgHTMNI5yeeoxgPNipa7Ana995ZG50C
l06US1omALI9vxidCjUV2rY3oWKKEqK2mH6a0XXl6bv2BuV0b/cMRbYckfXfMN7l5Kyfen4dWz9+
DeSfyXTtZb0vpRN/LIBaiY+s7rzQ3yme4TVo6J0LrLiNBPmF+dHcDjX2alnh5blP4Revw5MEQzkx
06LfOA4hZRJ4A6QrdRhnd8STfs/3nN8hEdPhfOXqsuRb4W9iiA24RJ4ekd/jO48FH3tFT5FBrNsr
pW0J+WoPZH5MNLHbCXCVNqktD5nP4wGu2C78I8zASAvVteUU6iMD9TNTO7V0QD5Zee8facQziwaR
goEzp0981kXoVR8bsbb77nGJCnJGu8PyS5/AukNtWPC4I65IshwEYXg1Qre6U3iHIuIrbOEY+PFn
0SA3GLigoyM17dmVHRRaG3jb5mnlKcn22lt5N7Jf3KXDde0T0uFFW0HQVZX5pVYp2U1wAjVlpIRn
WjYJCEV634iTBYXvmFEetTjM0pHmldRYqSGmLCi50Nh9hyIpWA2VjdpDcrpiMcgs4S+fwlD+6exl
sTa4VBn3Eo0rjTJdfJeBl+A+eY37UzEyWkVtCbPkieD+eF3znSoZSEJ5w564ify8FImn0d1FPrO6
ESKQwGF/CzPi0ylkmx/NKvMnJr6XJtX2tTl3ar0FgiqXugKv5QCONkCDU5t0ggSFyq32et0Dh4Gv
/Ihr3ctvy8G9n3m3B3uBr2UygW5ubW4zV7204yqRfCxn/U1HL31TQErzNplHZ7AH+QsqJYjTlQ5r
OvM9DiTWkhP67GWKyQMbF5LWP89IJAuFt8zaEnBmjjzvOa/CpEhj2Jk0hfw//q/w6xn5G5Kvw+ch
qlwkESmJZvFuAK8mLUC04UhNvj148MnswXOKdCPqjeTjzkDuaUP8I3q2NhbKSBFGtgf6pdlbL8yM
ZrlOsINdx7v/VrCgnnX75yTMM8Cg3oPEl/K93uebllgQ70pGr8h0Uue7YJHHo1o4s2PmerPTJr5h
wCZyzBPJqufplryMmiDiKazFK+W6EnNWRgg+7+CLOHcd6L+D1fcD/ZATa9NWJMN0mgrwzU+79kbh
XMMprHT6dgA4t6kPUiSKSmx9Lv0i0NUF3GeLtr8ymuyI9ujEtpkm1bSqojUzcooHS9/x8NMwmJkG
EiVEefHavkh6w9Gr1tjMm8JPXn6CF+1n2N2j9KhwKlY2F8TatttqWdn1i3a23x+o7NxBAGhCtLpS
qW16Vbfx61iuHrI/e/s59jnU6UTJhjORpzppdPbcutUYdZ3EuHgF7JTR0mw1sgK2uoOKUuA1vtqx
7tPCdR4r8kwUpjeUIhI6ZQUOKYXplBv4JUZJNU0bZoiuMzKOXZ1NOqkvFn232dbtVxa7sPXgjG5Q
cRZ/RVQ/4ZRYgmmsKl5NqEFdxKDjveJplx+NSmVQJ6/kSOKYpNyDxpHrkuCAyhIP6bLsmwAbkU8x
U5us+Smq+Xt8PwmJk/S3kE0VbIgVJ8aHfXIuLOqp8ENrdhoxMkXaXUAEjfhezZLEJSNOcZSryBef
KEFbKQxDTbyUUiq4bWATA7VizFu3J1QyXOKOfR10DufqufLihYMbdbIe3lLw/lIVnyKhwLdkUgyO
Ye7xHVDQEWfXCPJY6AqDsxG1KEF5NoLmtaQ5mAA3H31w+BCpO7e+Aef2eXRhW1w5dZ/nuo7kBH2w
ohXZ6vnLwsNKdogyo66/g30jvDhBi+KeJGwTZlleov8VRf8EWfL2pGeLp0Xczar2+VqZ4IkcQiOU
eWrAzrB+cWgTC0zNoHkv1BDMd3ifRSuY1dhNG+5SwaitFPBTmx27vJnfH7GK2gDKlUQHP5wD3fBe
6mnmWEES78tVstUx8S8zJz0NBmhDFRo/inQT1lvVPPa0KvcexdDvAKgtJPzRvZcaKRG546+r33WJ
wSqCwIpHo91XzprRbx4fIhokoQYqc0xpQSGlpR+oQd+PCIRzqIrq94fwXNexujRcKItdw/A4L0ft
pU/G1cvAaeVdF0650nKJqXQ+B1ic+vdjL6XOB1Fi7e7B8/iL9Jx17eNHg+Pmq8524q/lnSTucfRu
9pY9NZBbJPea1SNFXK4NV3e4lGhNog2gnp0gBu4YVUd0RORhMDhpVnRskNDotK5viHTZ8moiDhtN
6YKdK2UWxUrZ7f1pZpdV5oMzi33U05eVVocBwXel/LdHKa+gqsGnCNH2z9fjw2yqAibEhucBhxlS
nZ2/fTzt7sDzH4zS4I1yPJgs0SuBjum2Pw+0oqAnr5LkqGhAtZG27juvAfj9Xpu2J0uBbVzoAK4R
tomOItbEX/zx3RBRbNOmyed2g0qUJUQ0KBcqezq/kLfKDYG9XvkY1V+9SDpX4sT9tdxfh98HJ4WY
i8XhVW6H+2zsM/hzNk9bIm3Mq/uBOUJ6vitH3IDOze8tEmcZqalANcRBSx34A2hlyp2aF99cPyx0
Oi1uqv82x2bD2SOYSHyrOB9mtjnz+eoZ6UJ9BhK7MUi1/i4emQvdZpyOsZ6uE77uZIcL1MFqPcAA
TUAS+YKLuKy5ueSSUb4fQgo0siM2EIjuWkEraIdSuOqQdL3Poff6t7tPUZCC8hTE+/u0mmSdwm6e
XkKNz6lhU+G7bmXfqezwshIai95MSG9ipRxMGRXbhJ1HYL+B1ubx5FT8kuHkw5LBPBgHCnBrRvG0
KoZLYGbmyQ3gjV+jROWDu7zKf++wfmnX0y02EOpFtSvKNUOfO0L9uHTcIyTye6Gp2QCPKRejYYqZ
hkbL9aw2IgVA7gzAcnQRm3TYEfvtfyqHOLhsrsD4XxY5DlJ5Hb8MrVylPryx8bRr9q9qqMrCKclp
f1o6OP3e0OUTqAs6N7IM+ftxuv0PWogi3pQ25M00n+d5CLNlX1mdYAhyyRnbnD1vFo+lfeYj+o/N
Y9Y4LF9l8R9DMFsc4XcQ+jeM0xtCbj93SEA4lASQnL+4B5S2VM1GqBY8W1euJSafscNnvy2Z2yzH
ehwcZpnYE/HVt6fOTNCCjhPZDzLOEUw2qmhZtKP/sti+2OXByeSSBrmCo3xbW3lC62y1BGwhyh8o
/g2PDvfdpRsFbbOzOc9LajTz5s8WiA+KE3/7zco6y2i3tcJfPFpzsGYRNH9CoFOh3BN8P+NUF06+
QkG2eukSxhHqCS7krudkNktBp9Eo0FGc/2eoVEZVP6P+IplP2KM0rQ43Mx2NCWcn3/0ss3/eFEHq
5Gi+nDQcn5bC9rKvXPpl+GQm4g0m3nXb5JE+xqYik820Gpg6P4uweB6OzvN9zTUkW42/pq6GyFdB
R3p5EItSg1uEQ88A7Q7G3nLKJ4aQ2S6xdv6eGAzMe6CBwIedvLhmFcJntDQMzpFYCd7pZqDnmf9d
0xvclo9yPbVctMhrFVckVhLTg72PQy0uLaJC0hpIhHpTEX3pwAsid/oQ6geR8D/Acihgdlj6p9b8
P+yimJ58dFUl9kD/9Ya9kRQbd0/RJIxif1v7BZuJXosOLP5cROIET3UaXJC4VwcnwubgtrplUlp+
ZvlEMyEfvzqXrzwfA2EuCeuPe/NhWxNBtitzn+nYlRr9f8jbtEJ5blANbc23/eDW5mYVAcCmpP0X
sEwoSW9c7sJC5vWFyg09ICby+SWsFS6Y+ge3SbnlkL4HuZOUFtO4LOj9fQnB5VHVo2IjYchTljQr
UrtXAVautTKZ0YKa3ALszkWS12ZEoxUgI2sdSfumZZsATkk3tpI4eAb7SK7axNxZ2ZERB0eXBLHQ
6wjb8hcPzKQr5vNLgxqSBzXFXHGPklubRmjoAtjDpcss+Asf0MXH0ce0jHk7TVHVqt5A+S3tgBUs
ajl39Z2L7hghk1kq7rzIEMZqWcWA6aqd6K3Mt622b5p/Ca9IyFWajM9hZpNPBXtUVa6cQq2ZAvyb
TTLGPhozeZ2wRHftNyTNn7GZcDd7iZVC0WHqWyB+PvYVVw818ts+QONRmAWFgDdSoURIYUK4iY37
HbWHyzZvCSA4Zxb510nmKp4nGLsUsyHCARv4o/mjpSNsLx6wxRMZfIkV4DveVZ9TTJ93a2YPssAn
L8DZl2wScQCAV9lN0YLcg0Au258sNwGE6c7XFyWFosPUfjTa0FR9HQs3Z0u0AhRLPMSqWr7hAa0f
jg2Fd1oTRSXIOJfSOCDCAW/azBlG/BQm+ZJ2PQh03TsSQMHf7izVDS4z5AL5MOp199G3mYCD1gH7
zLWZyF1Fm/UtlAx86AJ1hz5943PpUbGCQGzJ+3lz0iWV33VZIHFh8lkN9DjwyZEZvrEQfQdasty6
oW55Jzz/xt4sylP2YMzi9arjB6nqKkLMwf6bSlwbPOlYR39Nr5JfLm9L3x/MRV0XxwU6JosJaxRA
EwP7GzJrb+IZ7/Q+NJNCuy5iIfE+739xViFBSPva1PtEIPRrzrJrcxH4q2cCkDFpVFtn9VBkGJMj
oEYBNTj3Nz2UgP97JdgyAe/IAI/6MQM7phw57Ij+CPX8M1RGmLwyq2fogMf4yuphXgAivUqrd3Ec
DjqIZ5CMo6gfSPv396bVKKprvSCxrRFSlYiXVDXJFqT+mvuEN3Pdn3nEJGV8CBpxS14hqZnTmhUI
PE+NNarloVsL4lwN1Zn6pOhPquOjnUkBUhDCfuCGZJhhPw9K0ei/Td2ioUcM2w1pBedCQP3e4A8j
J7wvaUSzcUx9v3nc+OtiIvhToy93iycXcXcj+LoSKb+Yb0e0eG4AGo44KQlDOeiNkEg6fyuqgrpL
i1gQhoCR9hrdsfr1kp6DsJyZtsYUzrXjSsk0V14ER35zwPKzQyH1g6Hdja0Hy6bptvloVlw2aw5m
L53brgzv4NeNTWMn6BY7drfNVCZprlBBvBgMCwMnnmzwNv1QXufUUSzQXJGbUQ1KSjaBnJJZ9rj9
IDEqGPl5hF7kNO55q+OABgl9CI36xa3+0tVeew7k0IBLlAln5CLYRYnJtiDiZ8+jqUrAypqYUH7y
yapCxkI173shwml5TgmnS4Ub/wAHYDZd9abqGYnRTYxOB0au0OvhZRyhjM2LP7R55x7rgILbv3H7
MWKO47GU7rArvZpxy32F18hMsFlV2aFT+vhv1uLth40Ta255Odovgxxl23OPRFLabFW96QqDo1o/
en2yJ32aUvM0bB/dVmZB1nGd/94SLAohtu37a3upHu7MRin9BKW3x/w9rbnieYw7cxKzWDVyKOok
WFibT5YqTkqrBGK6tjKPjvrjG86wd4Q1GKzcxnutNwznr2Bi6JpF3dLAMhZA4upcVv9Yux4oP/9X
JiIBdqnpS7SPUBC8csb9eI8PZHndgroGQqYeZ3W170EADQ89g0SelKORIwoHDz+Cmbf7R0qEE/m9
oIg+eJ+GqgqxNTzidN7XT8p7weMP2d/UTVQqTB1yMVQZzYpXIXzOBoIrcm0G0rsPI2sq6SCJkm3+
sGiFw8LZopoGqtd1SRnNSrz3nHg56w0Hca8htSdIyOBFRwK/nbXN4wBSEcAqt5Vxm8qK7sJALUpY
e5F040wIWI2hNGp+EHbY+0UdCgoSPHBo6yX6VzcPFpiOY9tg1DdtyhUKVLXbG0+ue6riwtTRY9DN
sdJxLodgPGT4Rp5/2A83C2KbNz+/ogzRdSmOsiZNM0n+edsvM1xDldwZSFF7ZYaH/WtgLm7cTOJy
msrBXnpNntLTtM360JpQy2KaL3aCO2r4HhMsW+Rhmvht/E0LwU1YI7PIjzTa+uL16TP0BGULkytH
mDLembYl/PxaGScWcXcEwSuB+YYs49tjPkAhOY9NZw8j5IJK+omKs247BrnJcC1uRz+Pr0AEmMpb
12qvIppiLdt1rle3ognaGeo/ObrUBZGvD06jziVOCaBNq+tHNf1iXy6hyK4mKvJjWY4ORvVcrCHA
9IQ5qths+X1dsv7jmFIyucwr7DKIkWh1weYU5dknvmZOB7GBztNHbX+MSE8ZL/hQU8/9fMEkyEqg
tUs4QbtG7RP9BadjReP2vmoPd6q5ziHtvKHiDnW8aqebPXiNPU5AcO35XpibBSVGFFFpDTuwWET9
kmbKweZxcu9YCTWrfAGsmSw5EOCVV1hYpF1lULJZxKzGT2tQlFyVxKmXpHDLJQJANCgRL/1QEsKO
Gueas6ay/WqdQDy9pyxNhfDb3zStEuYSZ8BQBAr/uxB+YQtHoq1NTqWTPDO8+0wzFh2+qJEtI4ND
aRCl3ExJwNSi83PFSbB+5MuefwGafrGQOYrxo3rLU9nZSy//J3eEzBxBL48Aa/nRUGdOCefxNNL5
sB4jZpdX8c8/TiLVmuh3pgeEmaPj3BxVo2VwKpxs67IA4o5XFXP3q4OStlVrl05ZVYSI8Z4oFp//
bqMwXKkUIG1Y8+EH7DyjjYNXU+4ycFuzL4Y948Un4gKw875ga6pXLHBcW3irPBvCX7xgUOYXHODY
CNSUA534eMRAJwb2uWAUXQwqObkfBPstPcKPQ6ImcP/vQOYxpxNzgt91vWGGyiyLU3XozXhjL7vc
C3Anc7bbJ6eadyFNy1WkyeLHtyhkJnhpiHdpvg4D7RMTNbamYvSA7n+xcH2f8Z2S9mas64GCvtIj
tQKehrSi0DsciGftykz3iku7AeYCw1w6z8TEK3Q9dByWjOTnoL92O99VHJUwIoK3tGUqH0kfQcGF
BFmD9PD3ZQlRt5GWU1nxOmpwUCiysDais+sQSBjjMt7rj1nHXriWktH7D06E/BJ7U4mcukUvc4WX
sl2gmHyD6xyuk0rOxWT+MbrPPjZR3VI6VFMCBJPgJ/owB6vo/Vm3xcjMDpT+QVAwg11M5SMp3Ys+
kRc1dpcxdQkxH/3QzD8G5gOb8ytrDzn3Kwz1Pvu8uOTl/vk75nGcFfRZOGtLXYA7Spk7UUv0bIty
axoK77na7VrK5Rkad1O0vcETt+jMuxz0FR8riBshK+zQUKeKg3t3BgjE0l+K+/ynHkowQpU78hGP
SyqKRl2SLMWCKwk0G7IGrNwmDXMxaujTdPv1G54RR6ps06S/8hvCQkYcQhek9kADiXjiN1j5nLXJ
IkBbBAKtHQb3uXztUvuHsGcphbKmWHNtORCOCfiovKwx2ppzeZZ2fR1acYX7qfhAVcfBEq1MZMPE
Ezhw42r87YhTEJkfGIzZDfiHXibN9NuSHbl7wYr/RhW0GJI26CBTrKTBH/u20IVxg/d/GkkKDm+6
envhcb2I83CL0EjdtMMaGGcSY+KhKi+ez2qy5h0DH1bU3bUr1+eDf1qKUXzmrJsarAZpNOx2Fw0i
7IrwMbzXn2SageAudJl0On1UjGQbgRx/rayFBLAHuAGzpLFSBZHbbNNPGBPtMmvHkuPhfI8OOAES
P6B9j32DlblA0ncrk33BPUe8YcaHxlUbOukCWWhxZlzjKhT2nnDqbavYaKjPJySkMoA0Jfqg6RTC
Uk0K0vZ9g2c6wpz3w/NIVWJ7e6LGhFKNjiNG49p3KwcnQfECx+xRdJXXsEyPNf+VQ4NoIc1pjZJe
FQFNrJUGtn5rKS/V0hIh86qGHFXBWIF6Scp/uYijFPbiGgEZWDqydbv/Hjg+Nbw4wUr2zXFG/Wcx
drIhGxjH+k3PAha7DmnNKeg05Q2SwuwDRE3nM30zFdud3GmVxSGmDpDOMiVEjF2Srla9r8aWQoGS
ZV/drQYPpSBurHmtWYW/nj63mUifHZfLPGSMER9DwTIhO2IbG1GA0tY8K+jhFQrNKt2iAZ1YLzoW
gYEFtj7qLOS+mUsQo0DwZHrHxZUPurf1ROthyNtWwfH42vdC557gpvbfu8Y+JQL+P2bgEM5UdHbI
hJQkRy7zpY8a8hL3DZm1Ypw2B4qbQZvP9q1lkysaWmay76/J4URm450tN9rUftw4BFWEIn1erblB
6ksin5xG6UUnehs9svYhvAArh3+vcbrgZth2hV4ByUh6/gMsCxBJBfwrmQz3yDZJqb3yaeAU9F5Y
EqWS4nS99wFyNHJ4wtvBmUYl9+WcjrkY/lx+1lZO/jgw+ON6WJ6nVQcOcPOdJ1r+qN84Y+KZ6aOI
n0NTWAHFrK9Qh8ZgfHU/bsHnaOmMEAh+rQ7puDe3io2ctazBMrVAvGGP7mgM/TGRD6Uba3lt8xzz
iqhVEXXxnDw++y3qVnUCemAcdLrnXXrN8AZOSlhhMvTZw3ODZHMq0u0A2czDg1+wjhwV8zqTYUuU
Is6IHw+4Gw8adAWp1zzQEm3d9qDBmxAQQ6Prq4mvWnVxRv872/cXgdRn3MottYJ0CexMFx6zj2+j
Hrt8r66RGioBdz6hxto2OHfGBwB9bRxJJ/4X1GOvSSvSgOqN3mLzkSo7ws8R0I9LiYncsSF5K4I1
hQRSoGmrw2qiEKJTCkCrJD59FqEzzmQXSzg8AUP9WNy2q3fXPnTV5lLiHKaI/pNa3rQgaAktoZIV
oZA0apjs7Fx8BUh6BAx6wq4/n2t2rA2lLwk5fsIIMqUaGsYEu84VjbsnJl0reSrhgCjXdQfoY6t4
6awGuq4+NXhAVSUDGWWO0+6/StdsPr6u39p14aTszWyIxdF1GPtPo0cclBqEBP2eKvoJD5nSfsu2
eqk7rT0HsDGce3Ja3YajjWjpg9b/CWwhhdH0U7Z40IfGj+WeYZ4mWny6oGXcxzr2yQLa+GPAYYl+
dsgKyb98Q9nNBOYkDltxHX1ihHh2dm+i+KpUBP+8mmaKhSXkOYVxr/MT7/ziEBGJuqs5dfzUSVi6
fSiFhtWEHt9DdEVQqhTX9het3Nuz2prZmLCLJceVzF1tjGmrja0z3DTauM5Fw9Igwbm2iV91jHwP
wkXmWQZhnjLTMOll9sm5xoYCt6bIpVynSqrOQ5ITDvtl4YV550sX1nMuuXdLNL9g7BsCfraDwHUu
UtsmB5efgVxYjJg7qMxP/ZMZQ6dwFCt8JhktT1DR1tzRPMc4WGSR2Cu8x2rtzmPiIcME4LdOaLWd
tpI7oNq6htFcBgvgvpESCsBi4krXVAigUW15nzU3f8Q/ok38TYrX9IIwUo2mPLQK+874WHYybf3E
NQeO4kuUX/DGGzuAOp8NL7NVyrFEfv0/xng4z+uA6U/1xraI3FuNPbfKYG0V7mD6m7tPucPzFDFV
k/hUlMs2Mj/K+ou3OUa0Jk9+T2U7naUtFWxBVECvXCUPCmTzPnidvt5q0bsowq6r1xfZtXATR+Sg
85gMe1FJEFea/8PHgKvFVxFl8yEcToREFPW9kCs3I4o24ozVoimwsm7HSnU7DNjn9csctBj5kVxL
V/+LjcUFhOV7WqzRRgrloYaBc5fY4rVidhXV8Rx9TPZXAtVELINXICxp4BH0XlqK6fQQZYBXH+gr
Kd+a+w/xVGcbitNTupIzVzbEh1ozZB/1cExGhC2xkW/+5VH2HIsqAKuSTc2mN300F7mwOSsYElR0
RSppENDs0hv4kkDsSDCvSh9tWZinRwX+vhOd2rermuT9uBVxhxw1TQT1ndkDBbvRG/NGxNZOxHzN
HXKZhjXGzMzC6AAxKOgpdeH+e6LrwHbb69LziPm6WTzxGB0G0WJwzAmwX0NP5mRNzf0qucclOIqw
QKbutCgXuRiVWY4exeM3SeeTDq8/+rN3i2cXMofuDro6kUtYnSEhgNuBFrrB+wPnLf5JJyqN5Xcs
1F2MD4mYd4KAkJ/5oRZoR1XiUwdwjEl8kvIl3fOZEAFly7hyvoN4FXozuv1uopJyShyflvDYpZDV
zrRQ+Qa5jPkx3WOdnK23fKeFTBx90kzwJ/O1NQYOQnTuX2/+1XsEyK3wqkZTap9RmItOD25m1fdG
83jH/7O2zcG8iY1viQIGbJb1/qErNrE/kCeWQ5UKZRlKgV5qIGedX6aqivc43H91mEiUY2c4cn/5
oZj1xwg/wEKZDfStd7qZnJfLcf1iGWWy5XxpHOaerWqIVOevh7vlZpfoayZoI7rjSWsPLtzdFvi7
kq7wtlnI3npIXPisJ7Tjnx4PveWLdkz3W5+RPsbd36JwsdwfwmjWXmQ5rH/HoG4A33t9yrSslQ5q
61H4t1VbG2y+Cv91YgySA3sjlpDcJCJ3h5HZpPcyvPRdFs9dFix6etJPp1WMYWiEjk5x6imMx0aD
kn+UodGacB0tY2hyqnY+uGDhfkt/XOMHU5wYQs12SNyEHQvQ8NKMeC7lmUqPq2zjy2M0Aba/uY8J
8m5JloGfHw3fJ1K/3BZRZNyFtXMOqx7Pkz7v5S+V2ZSqR6PRiaGHOmhrff9wPTkBZo9JbekLR/Ug
Ar0f3sJNBUvXLtsPQ5w02kef7saXdi8OoAkrlupIwVYioaBEAA3/bE1sHXYGRv1cS1VwhOsiKEvm
8rueQqqyJscr1j2AhtNHdrL68GiEZYNk0Z4NA8eRvU5g47LPUjM11h6AWM5AlqyHTUPsg73mAvWd
J0FtZkK6Y9ZD19/LXwD45VVjLu6mnQDJ0gNmMZIGw5Z4IOyixFP1kCnre4AzPB4TRbeOwAQnbcbb
H5j5WlBfKDuuZwWR1U3yitz9c8Q3/pXL2xSV4lPZnJaeANkvi/+ioKr61YRy4qevEG9nceAEkhNG
UwXbmn+AbsdJcJLDXlmLVGDhBJkDXxep6/agp4Qq32ETpaw/A15a6fSlru1huEevKbGA4MS+fCwI
vNxd+9gMazyBueihywPbX45A1pFnDYT7V66szyqV624e0f8dfZtcCaAmOUDllZx2pCk8DuusIpJI
9bza4P6owf/fjyPA1vYTUtX4jWZ3xjhOxQZESieDkyFspBIhd9pyvEyOiijmECxkRBZseWqAhyjq
HLMk369CBnrxwhRHhqbcmDwvezGlZ/w3ljUHguUEH3Cz+0qBRTnutEeWCC0Bo4twdrfdZ+0ZcbX/
MhUYkp4NUJIAd4OhFXu82MtoZzjh3cd9B2AqE+8dWXBgLMZ3kh3OBnu127LAiGQSGwY9Bf7F1JTM
Hb7x5laKCHE7R+H72WLjSRPqw64N8WY0Ae3chzmlPsRBp1QmSLybUDEqym3JND5C0fhbxKaeYDrx
4HOR2JSHuN364IzcxamU3D6gq0z6LNmwjd57pAqmy7UZDQMRtQFsOJc9OKxQRrPBnoMXRyci685b
U9vC4DUHDUdwarauLf69QwcdQRCTXzkREFnNRPal2LIU1SvzCJOZoDO8mreq4YohBgRJjo+bHeO2
67+jBYaFsACYOtsHHKIJar0V7t1BOL6c1PoSMBXrva7adsukEkGt+VutoeDmiL/3oWuFlz4x6xTS
esjVqOxlS0afKU0m/aXIQtDRhCknft35ttpigBCiW5d3bOvbdidCNP73A1ig1r+BfKoz4riXHnPm
CdooJAf6VYWvxnQddzy8Hc7w20eYJRIKsHgyfr8X4uzp4k7FDhEk1Fj375sSRKUOCj6G0XPCVu5I
BoH94rCgjqDb6hxaxnx5AvfnedEt5wygwCVs8LkTFTJUPuAtViReMDtUpr8s/0M2XNm/PtT5Cbxa
xyIqvksYci3KBld192WgDLFkM7kq/nBti/boJCmhX9tvFDTWxeFDxodsB6/MutuP4w1ej2+F+x9d
cJiEjsyRjK/QbwDQHju0yWWovnqeEa5n21jZKup7nMITktIyqL0afg3OeZReu2d8umPJrPV0nG+Q
kcLoK6ruv8W5+V98B5eYq7oNRIjthojnCq2AWnK4d3CPrhaw/EP/2F6K2v7h/WPCx/PG9q14BOEr
oX87gruuoLrCdI21EM38Nz563fnb8Qla44vud/NJ0LgiWIKrVN5TFODc/clx/DA3JNAJ4OjGCI//
4mmlac06lMme5fSwla3y9CdMvj2TnOEEp9Wq7KYuBr+3imeD0pHPvOK8Mwxd4yK9MllVxkK9wGKo
CrELTMfYohg1WQfpg5S6k8tPdil1yCGmTMpqTbxLpBci/2YuSM+8K1XYF8AzBaHg6ZJOAFMwo65v
hrrBd5UOoqmUlEn/iBKRmW2LYxDxLj7BOilHfHq66OLMXntaYh58LJZnCP4PNzPk7YrOXRyt/jx1
OPAzdZKtKIUXUBtaZfvu0tEn/PL9qyt6/9D4gpwogai7nPlhOz3imUb1C4GekdRDMbb1LVArVU6a
hvUkg6405H1F0J7PYnW6bnS87ZpGEpOXkBPz+uTa1RpFuxqVRN+sOQgSl1joRoaNGN/iSCqH8Ubx
vBY529jbvniMqaevImq+ZByjho0rabiQ/ZBrgoqgPpjPrfNRPnDlTW3Db2UNPYpBvUh4+HwRV5b+
ohaBwxsJdNNqYiT0jgzS1q+OqSCVcPRyKTnnqgPt7oRTV1XwKccMoL19VPE+zFYOwf7QH46tZg3T
xZ7D9+jDDwmkATZUZX0ZWb/4W0rUt3WjRTrvWI55RePOutkUjtl+3bHBbhp2OS/oDVRJ6ZpOZgXz
QD7H3pK4X9eax/0gZIETBCRfijhQTgzR1tfc6LxkWmIw9uk4DyMtwMctw3D53SlCjxQx6vpotVjb
mJFQtltnnWMJ2fD1K7q/HoOBVtCYJOh7+q54GTcdEPnqTtj4senKiY4GsF5oH++3YppLmPuSwvvz
DSUGku2ofGaCoZdCI7D+j+x2bdyiQdtOxxwIsp2M6+GYbtAjGIxqZB3SL6YkLyWnukxjM1QoDFWr
pNyhGEK7AIM6q2vXOaBN9hk6HDkW9gRJnwWvWtE7ray+9AbtTPmQVxWRavyYhZFy923uWw4hrP9l
rvR4Tms8H5zNdOQ4ddABcVuCclt93DwjRXAZLuk9IrUQpZkWzBbsLWPohlAwCK18hLhelTSg6AHf
njCdb6WPyFuzNOqc8V4n7W0a15WPdReCUsXsE52oxX6jXJDEtnhHvvhfO9RwV7g5GpMSyjv9MWgF
HLSMUktGlaFgN9IXgP0z7BouLw+QHgaAy2iBnEK3yGBBbLL91y9lSr3sK5NNZUJYUobyE7w9PNEX
I6SlmXeyTjJhy5MSlCsfaXlrnQ0FfFsQrk5ezjZdjio4H//SANCwkZhnydlss6ibEA5CCQs4/wM6
Tg+pXQ2hXOnIlEx76Ym/oIpDLbs52q8oTBS1lk2ptIovHX1s5ACpx0TGVBwiVB97dLVqmD6F15uk
cVuIBEbbMzBkN0U9nlvKrVUXF+ZSs4UnELuJvX5Di2FAL/wFSPaT/WJ+4Lsye8mjQHQNubZGefbe
K94Q4M7Jnoz8JjfpKU16tCuMDqZK05C9VFGNCGjkitp+h23QkrSROt+6Xhp0irnuZFI5HfwEy24B
iYVeggTGItofXt+/cIyZHcEpk5Bu3qAfrb/4IVIT6mfTa/c8HC7+QXNamlghlihD4mrueLpstCYa
Xdp3iDE+0QbVnqxgNIPfBHMeNvnZiV/mO+p6bEX1Cf9Er0M7NLxyFF1rtcChchGr0TScp6i60Aqz
9ks6FsB5GpdxV8GMpeOGK0anhWYzkJ/cSdwiZ3BhhnkQnhEBRjNCJdw20nl5wVVjQ7WQQZON4JDL
+SXNOUzRZUtqBcWnRy7dz9Nitz07PEgN+bvBqx2gIQ4JcMBw7at1hSRVhZAHDzt8XLWdkk+nR8KN
6fdNoEiJ9YxQWZD38XPjmedSlkYpzCX27ZYjyiIbemAgwjbWu1HAml4FKf5Fawzp+UTen70g7vym
6rHh1OUej5wjQfOki7ruaPEeu4Hk6rELrbUSMrISUy0mm42C5KWjKFLo/u5NzIE2AZq1OgrjA3Y4
QjVXa07G88TqXp5G8I1PuE8Y4NmsYAhs1N+vuSlwb3sazhodgr+crrYCgyDwcvnlGROe04/0bTlK
/XN7OKXbiTSELC6aWFFyHjZ28R4QfeqYKLydgYwgV+ewefa9+T5PJ3azhDKDQwZjJ6svtCvwyMEL
U+IfRgiBPrPt/O1DtN7dynjNnokZfKBFjbx3fUFgSSgzn9nLN+phwGq/qGdrYvJGFSYx/UzE2tI8
4Q76Ayx6X303pTgFd6L/KvZ25R9kmA8FGMfukvpgiYtKWG1ldL7cuNO8JbXYQdb7wSqFoX3g6ksF
AFI2iOGsxMhVkKRIgfyiPxa6UWzS4ZI+dcFFN4mFlnol/uUAmuVOcRbcGQbVU476fxdJTJhTrsLo
sG19onNcCVV5rCj4XAulBkq/z/Gp0JFN9SJfW/IOCrJM6lTHpBS+PhuJD+oNYJwyjuMTswK2Bv5H
nwsr0H0gtIxd2Ai32l5yZ6KMXrTRoHSAOZ3RrRE3Qz5hj9yohljbsVSiiQcvY7yXnMc0pvZiT34w
DjRlbn6V8hmlF56svQEE6zmssL4bj7WMSIVC188kV+rNb3lJaZd7z9ipPty8i07f7ReUwx17RqAI
x9nolXYEJY9BUyUn6byhP+3BPjPGrS2+ThfuLTXSc0IEdWqZDu3IcT18yekPxbjJ3IWQ0+AKY/qF
ylQ444HJvqhczjLIrdmEliyQF7nUTpUp14Q589JKwcnn2c6U4UY6nHj1qBzAANqwqfmVwEgn4wy5
/fJEd8/J5saSpWEy/keMZ1oim0ECmQlekC2K2dfoXxiJrKv0Lgyqj94Dr0mF5wRcXcM/l0GXDJVO
/q+7b8JOscisXh2J5h0SqqH/6jU/mcsVHV+KbTsNswM89ffYCeLc8rbvUtr4qzvgVrzr1qnWY7j+
ltFZJ0Y11IvxCI7iJ/3cZ7XAreOWUmobP0qcQwNf4YK0VPgf7vGigCzVVxC0pm+aW0Nzi66dDYBF
KqblnkixUvusgJ3FoWr8ACSrXy6yAResa6R2evAYqlEhMNzZC2rFfTrbFdCFlmwQfGkEZ+xqUr9Q
6S1mfBd65cb0HYjniaJpPxUlJQaG+A20GDtwvUSXfylvF8xfvncO9bfONC4KK/2Yg3uu6SJypkDk
WP6D2PUFIBBTI9M8pV52u7uuTIMWs/oxKY1PyVuFNE9UAeHmaWvm/w/4HHE4J8cU4rBoqHCw0X9r
V7Fz7hxRusMzD8bOzhmouRJ3qgpdOwQI7xrq5GtacGj+dTUkDtKhWJfA0yZwaCWPiq2bYhof0DWl
GyzSeN0cY8z6XjqgyZcNqXJ9A8aN++8vujTO9Oy3AcICe4841VQ9Vz1kmNKasdNoX0cdNYYSnXgf
6Rn6GNNhfqJJp/jva9BbWAcYmKxqQKzokDcZT/Bdif+AdIkFbhSeqW8KiaXAws+Wf3r0SRAmMXsu
Urw3o/aV2ssNxv9zs7GB5gRyb9FygmgIEBy74KLRbOZqhckT7c5BK78ALxfxuV+3QvBRh2GLoKuD
3IZJHJVDx0nlR8sSwV9kGqbz1Tm2O9RX+7m1WKO6d3Uw52mTDo4gqfw1rEfb5NblsGMvHHOVD+8W
jPnv/CMBzEvUiDRM6NSbtQ+B5hc0MdO+Xn0KvK1gF+edCAuj0MDhUmg2gRHvts7XbeImg47NPVVD
lKOSx3HDKQt6M8k/ZRYDer0L3dqORPBGY+bSRPS8kwzrgM7cwNDernPkH+rfQfwWuhVlYyV7yOpV
ZnaHayM7idUaJUIHtLD9ByWKzN5BejQ5aEL/z9YcdaNCGcEk8CcDjnR5sWLhLfcIbujS8MfyeXAd
iD59fM97IEgIAEWWF8VZkXT/82+R6ZOh2af8MOWkBEU3CkdS/h/zOSJgLzajlZl9iYFWW2++Bi6C
94uErHr5CEp3QK1cy1L5xOwpjKv8vmQLhYeN8KjmsiWB/rnp0rIyByoL2UVuaiGuLGnin5stS/oe
dt8MWt2F0uFGonMzFomfuea0Zxxi93JqHMdhXn2TBPcsEKuCaUYVo6LhR/QaIxjN2OWRw1lLLyhO
PY1F6AC613LL4TFnyeER85OPoGeS+P0D5XkQNfXrcz1gmPRloxX+CP1v0MF1qySBPw9JR9UIHJ1p
ezbKTjB3zfQl8UVwePo/qh8byPlmVcZSdTbwXpBlKvi1Ga8mMUF/47UUCv4oQuOwBj82I/i7jRVk
ZvJI6s+7ifdBEDqJBAviNDj70lDUixbH2GMTc1fhMSrQ9uTq5bBFvBoR63MLOlfk7/5tKKyhkYck
axsmgV6PRyK0obS2FYc1ho4DeZJa7o2DaThfC3UfNXlMRmmWMLvXQH4V0NwmNxsBvaD39Ko5qUmk
zy/lVGAPZ01PuPDBrynzowg2FXj0wUH0RzO7KD8KWnORRS7/yPIw7MWT5EXjIYxJbUf1TUe10G79
66s1WCGRbIfW7NEy0dm0Xn4e+GAs/zmEOdQIyQLQxLwnQ+QXYz5qgd1wK3yvtuTLtDwTFu2sKtUB
4BosN3BUbxpTg1ZTw1ogMz7fL+R2rjY9d+jWPHV2dUVVLF9KAP+HsaFJjX9tKmosVE3BW+rH0Xsc
46DaYB2CHgQKfA32C/QlE05VokTiZ2cGxYPtXBdP/4kkANrOxpw7iF8xGFltZj70qbHlssne2Rjw
OVhBmlNi1nfSIQp/91C4XZlTjJ/TZiqYpqGcdfW+/E+cSppMQoPUGmOyytamuRk3izuRJHwPrmuX
C3MDZosvPoSkh7ZVsVqtpjbN+bFhLLhgdneGcZdE4XGTyWYDQT2kfk7AUsXVQqJ8ixCAkZNEO+/4
1DuYJo7aXyWmlG1MT4t8vuBSjNwi1tFUJM4pVI0kAVDDMO2nJW8ZNLfs1+MXH9miPWUrlz0h7iKx
tHfKBVQX8aqOwHYL3xt/iWedlINn5WN7xepb2oDGpyx0x8C5bJZzhKkq07XM/GCmdLgulNGOj6Xv
9e9EReJKkJV6M4hVTATK1IO7MY9anblyP/e3k7JyXaFsbCN0tmQGzWCLVylvJerY8i4S5UHczfX6
7Wtlvn5t7eCfpgGwWgN5IoUOyXdNOArf86HGqdtnPTNxBt9Smp0x0mKaQz7DsDGqToMFacM6KqMj
VLa08T7yMcczs+2+oTgWt3McJlgQV3yL03F4K8uWrZsx/kBovwZlq74oz6Iv+OHzIiu9+/rCmchp
DMTK6TCf0Q0dwCuiK6R1CQbUPeFnwdzob22VYRv3ap6JHvBKFKzZ4+VTDlx9Je2vn8VS1xrvX+FW
48pzS9T1kNo1lC/nBgOlzqmqXPmfkTzjbDoGp49UcJqFxR7BuMRljZ90ffa3TS+Q6cQvecWn5pGY
uoDrHj8TCSIW0dALa8T84NMRXxMV/kpJmJhUNPdByGo+flls1VSTRoNB6PkIoFCLbzBaip7dap4q
Ho9D0gkt5PBk+gSD9EFJyuJD6QVMGzkgSeA1FBE+M3fEt9On7MjsiW57O0H7CNeLIZkH4EuFwuWu
YC7Z5f1YH4mLyVzJxfkTtOJYA+NyZkFR7eRsRddQQkaRSwILbbgdJw7xBoPOVypclNUYJr2/5EV+
XMAMue+OAvJBLueKJo5nAnJPkfKDI7Tu8bYM8UVYY16oz6D60iUtzqj+NSwkGjBzH7vtj+w4fou8
AOCFHkp5d2iSQUVK3Lo2cjKmBzjs81ioRNJsRxo/oB5sHVuY75S0cctlPwWM/W5fiSD6Zxk9+vrq
k8lfjkuiiIHAyN+BleITmtDp7ZsSAxQwg5Z7gRdAMmcI3uETkC9NlcUoWsZmL5Njhzi2zTXv9eMf
GRzhoXmbHjp+hLLUhAAwrIWFYedbVGhK2zZjtD0rfveLFtVwZEviBNeiWwO1RKj3a2VKm6naZdAw
equV6bq7d/AYL60xR8FWm3MhNEXozSYOeQcfEq5sCW3BeJOSrIuAEsBtOYVGS7qYWus9FH3ZMCi4
B0XLD9QwsXA5/ldVNJdvqPhPDl9v+VNygaESa1PGOk0ojQzIVyNXvEEV5jKhw86P0PH2SZDjgJcz
Idsx/v9m2i7g7plONnQmMOpZZHxDzj9u0CHRif10VIIfwN5BCcHSsy3P1vc4yZCxC9v1kjSqUx5H
lrzsjQCiuIj+xcjzisdatBbLYerN9VtTGu0034phDppWqlCDXGxSoAcY1Xb6oQZzxnqkpij37D7s
OD1tZm4RmvNnQ3qhKNcX4wM1e50tYHGoNe0eambqAVcl4y6omgbp3aropVcndieTM25cJdbvwblV
HfOfK6PLrW2i4VX3cuxlIZwb/YmkW4/TKyzmoIoJiWUVfNXum4wbCyLtVYunDXCO2zq1uN3JwPZe
b3ggS6HKc+zKNGnNfOcXVmyYen4LndyT0yUuPD8KhW5jpFIhTz77i9tH+c7vErgTVCtcHEM8GeWW
E0AXA3Ubi/KKwwVV563VsWWvau/26f2aIYLume9sRmMz8iY52zDIN95ZDLnJz8zaH01a2iv7LutT
Rn8hxwBZTxguHQpUlzG3nZG4eMw0mYI9EkuD2V6Q8TOI5QjIqoXrI3YCMpsacYCNQAST4CUXAoqV
YOz1H72ssxZ42q6W5DQT2w7+wunDKQaB7LEE4Ws2A/an0l9cCsLsqZLMLyaptEGQgMBn8lg/zhZV
Tz2XgkhAO8A/luiwcfOZKahi9zllCsh3ENwcBaZr2oQBHl7c7qrpIpqE56Pa8VD+lAXDQdyMAS9H
2ouOPIUKzm6op3KYAN0eMwejVeTSa641sREkePaKdwxorEHmepk0pZsU0+CX6VJfV8f8pBpd24LD
g8s7kHVaMlus8AKRkgMAb1Pc6jImehr+qAIiSKPJXqCXBvTnqj54hFlLnQuu4XH0I7Xyawqfn/Us
TQBdewFIehd93bTeyRp1vy7eIax5s/3/G4dRG4FJtl3XLMlG8Jy1VOFjTAaxVM37KXXT1v4GnNi7
tw/XF9KbeXra3zpcRg6gzLCB1Ej7wFYGimZnlayex5BcIE8Liraf+BOBdclm7mW4agIegpxtfLP2
lmkMiDxU+ZPX3r0Ry5bzP47D5zUDXScC1pw/AsvBfUhX0HpHn4rucI55Fce26CNlzH9GL87fZO5P
K/gFROUQD/JHYf+Vcr5aiGwnu8VB3HVUK2zFqYSlwsPV3N/Zsolt0cxXlUnv9XZFH9L3kW90fkVE
0lJ/0wxDC/uc8FX5kpPW8R9m4z6RGJ8eSDb+J4iV7x46eiLNykO6uAPLyUNN4Iog8BlBx/J3YUc/
HecLmLJwJFzF9tIsiSxTcbTIBjNl1EFiibm4OkPeRw9cuVkWlAGvVF2LB4NsBz053s8BNhdIHfrI
K4JOomresbVStIVtSydbE6lECFyapXFrawbhZU/cpTAQMb9uk+LF7TfVqJvphYHzKWjV9JUHZ86t
pP0mhqHdLtMUd5TZMkLbDkZm6iXJu8My9rMkTeURHTzzrAyGcRpzFefHPKiinAAkPALeSYPO6axF
R6BBY5SpabWXSkKvbnweTyJ4T54v6Vup876Jcv/tvI++CT7xA97Vjon8oYuS3IctznoJnJoDi6uH
Qd5zXliyMTlwcXGMn18/YobNONx+yiMDkd04c2Ub2YSZ8Y/XIaRbR1/mdKvadQ3/YwmWVdb+yqym
M2q2FTavSuRwPv8SuNi5FD/JjIwPsewA/cbFtDpbEbSGfv5saL4Tf/5hdR/roEAhk2aTP8/8uWRv
FZGumr6ohhnt2jKuCgbjfA/HHDf1Ur3/9OF/KMWRVOOBrUTfy8nYYyL0/rXxf71cQgp1sI3Xf90L
wwTC8aNgVwUtlA9CopeRg/jhMepBvNaEu3YhRzaI1w82XT2+PxYVMXEAWJjay+Z8I4Ug4Md0C8Bx
f6CX2WIXDBrZ+VlfVKkTKeoWDGVwfPIjDk0yyvZCWnQUYhoArrcduwXPoPSy0p4XmAnkcRIeeK98
RnPcDW5Yfh50FwKjiy8gDlJlXhGJxphEHJdt0nRUUQDMO5HYi1i5M0CSf3XVrwrsV+CHNk6XujmD
BTeN75u7BkyBIKGiKmbUBgZWbeiDCb3GNSA75ncGk1Z2vRU3W8+buZtKOebQFhCP5jsrrNG/qvnN
H6YPFqTrdGctr1Jay7BFOGJIpyfr5G2wfeJn4Mf+5Tt9y7JxjxRidgPf0E8xstIT6fgtIL5+1skJ
OZ4N9iJ5eXJYaqmDFBltr+m0qzVFKetU3DzjUgblR2ciaku7V2RoN0K2sKECgpEWx0MQcqn823ae
tZh1bNc2TUi3+k1poouCtQKQiX371OtjGT3I5ZjPEkzPwRY3ffo67nE5E26OYtmtufASrQRQU49T
TsVdCC+vBxmaRbXo/BnoII6P1jvxrXip2v7Y0NR0ympLdS49vua/JaumwVVW+PPH9eDOA5MEMSq5
OfQs8pECp3R7tiYYj6FJ2kY8vA/WD07EU38zpKXRwpzgga2kxi2AcviLUDgg2ga5p4R+E5EX+qhR
CgFYvuHwxDy91VKlmfKAXne1jGwwYpcrr7mh0qkZ3wFkTqMTsbzlx0qJnXP5Nh7zyKjfFHVwbddA
lKY1f1tiNXvoHmkLxK7/7j4tKS3Bc09fgmziA3VEKnBlscblh60WK2L4OndV1O1EjbmrK12t8Bph
CZB5lcFE99A0Ih4YJ3vvJAL3MocaP7ERZzP72IpJQfHjVOUCKDSbTmY+DlCwS6qHbvB9mW4oM77W
Q2hHL353WZgWHSiAzYjOuPyEWyZbjyY0sYnRdWhWc57D444vRQigh/QoGCFeATQIVl8KsVVWT9m7
PYixX9StM5t/c45L3U0uX+UnM+LRM9I/rQNkBGY00VQgfIbQkYf3pQFW3SJ+1xljD15UF8P0sr/N
YX2muszfz1qbRoeOMmCsiWTDCaxw94Bw/yr5TbYqBGyV227J14uSvkPrHYCibzmg9An5OmL0ZITG
o105Fix7qWYDyixNgso/QygNwOLfvGKbLMnji7R2WqKWpckrfHktaBTlDpyH1HzC4qOVdPiYaq9k
Ugo8iA7byO/rMRoMHmq+lVqJze3ZNGq1WdcgtwErn7H34EOnRP0KaiEUorQtCqyEKBgaImZb2c+b
gHEAeCw97whbqk2aJ0YK1XXz/8PEm5VC5STgpCiwqlbHOBjYJxL0hej36nw7s6D7nN3zgftY8OU2
2/kO9fELbg3Z//aEdOb9NiFClbGuZgc5vrv7o8gI6mZYtNSngnIa5D8mZbL6HtTaemQ+cMaLEF/G
TD+eZ/D+GkSAMD7h3kywrpMtzvLaTRMIShXd+28CHAkjzpXezY2P7QF+WUa9B7gFOQJazfwqwqxW
VTLNu0fX4Lb5wjthUfDMw3BCd6On8u040IQn9W4vZl4utHt0y/cP1UM7GI+9srG3gA+hsn+bymvf
FxBzqjaZw8pE+7Z/Et0qKcaAlOXcpIReOLoiNtMWfbK6Q37EpXtHm5FSSNNskFHPjILF4/A4wc7p
nxJW+Fc/Vq/bGicpvaBujMoH8vSOFbYPCoxY50/NGNYkyckxkOWUJFQVhlqMvg1+ulHXSS5UaU4c
bCv9EEY8xxM6x5q1HF+XFJsG7ZmaSEl14ZW/qNXKSGX2FzHIb69Hl1mmn5c/aApLnqn47A6l41Bk
PYK/pOWoaJflxOA288aR6CcuPfZ09Pcz+keA9V5rHwsIDejCXLTQexLv2Dxjd0eyIcFWUPxxFf4+
Qw7mLSlRx8jQOK6W0WtiW2P78aOdYlJVrdZ3OUN7YWpKc7YpMT+j3axIUsJboFuj8KHNhKAQeoUt
Dl6IRExVb+DW+jc0BqBeZM/3PA8xyDQEG+Wm4Gg/dKwsvH2aE0Yvy8suAMud4QYRUA6DdXYD62ON
NVpLyjdLyf9gdrOlUX0ChELrS2CTLVGZTrjPoNw6YmaZDVXV7sjaUVfnsqCr0t0NIUU+mH+G7h7y
LAatLM0/B0usQmDGDnHFNTHbfc9wqfI9jQTx8Rbp6S1Trk7KLrX/5b38Uj0m5K2eJjUQljhOon8l
iLik1Xf6ZMtn8/JytwS6UfuWOAOH/eabiU8ovGrvtFB0MlIU9PrqM4A53GnOzqqIeI2x3JxLtwe+
u7a4b0E6PPJ1jiNkVRvWEJfIrnMdK/aZ0WTXAJ3g45khp3aZk4vyTDqxIuxFSLSbbAUDUOAXRFCJ
WFWZcP8awckle1NdJXyZ5MrCDQqEXomCi8BH0GGi1TAaQ/txLcSlwSlJS+eK9f5cjOnevtG6U8qH
uwm2v6udQ3GDeRll9y4gPK68CYmacuwglLiTAZYXiVodFrBALmAT8pASSZxDyBV73TGOQQvUEuje
yC1AK0YyNHGJbCrBbO/dKtRoaa88L+d99Pr5dbXQ1PHvacYj2Yfup6mQd5s3n85j61x5NifLBibr
jVPOgVstZc33SjKz3i/b5TftGQjr6CFfseWZ2hno9qlk3npKNIMaZjM4EDsYdcdBPq0Y0y4pVHqi
0nj2HNaVbbEIxq0NiimKqKn4quVcMnkZF1/D6Ld0Wt4XhirR4M5uLt4eAIMfWgJ8XSGGwa16G/Tr
zNy6m7lYmsVIuuWsmLnGjeW/65zfz38x/AtYr9we/Bx1kUfBvYAbgrKvZXRE8QKE60hvHJ31ZNvx
hs0GuW5zlGbj1yrggi4EI1XYCkH/ZjW6NDV2PwiAgSIbd7pmo7ApIaZfaMVze+OVxaOEXmJUHKoT
Mgy5Es+Q4NTpD38XbfRZWC8I0j6eyWKU6RTxwWY396b1D839G8ypFXd/ifIZVJq0VW0HvBr1VJTm
G3V42+ozHw8l0IWU6rYA2chQwmvaXGBBCAWl/lRTLVFPQlp3kLC99e2SMm2N4ec/xK9c4Hk4po7f
OpEE5nRK4bpfPGDDZI5BYAHPl45u4/fKBKTkfxplrj1ZxDtL86Z21bMMN7AWjHgm139SxK/vKl6u
T+DEqfGkc6GMHE0Z59OlPp5se7eHjJO12UaY2gdB3j835pntF98kaDYxk6C6uNFGyBw3mJPSKjKW
OXi4OPweGhvqMtp4R06hHi75v07mPab3ZjZ2KZpReP6I43aztyAocLxpIbuUUUhAhfz6MixlWiSq
mFMln5IY/cc5pkWWCN8hxlCbZ7NertOTYQJq22bk0V52jHjQ6hOzjs8D7yuLxXlDmpoDJwJEXOhZ
/whEaBieIDREW8HyuOGkg3O9LhYvKsH3w6zMFealnd/O6WUsyz0w4IRRIsoEOcau8f9X27xWF8cT
zP/n8yi4R3rCtrn3uhXdWru6vqUFe+ehGqc6/LlDc9FW0vF15BDLySv81t2pn9bTntwEiLexu6rS
xsULPIjaSXyp6k4Bi2pNueaQOC0ujU15vTYKoOlE36k84ne1kFJDyOI+PCdG2fAyKrkjTDlOIF5a
fozZ3+F9DcxlHKOS9u42j+jg+62H5KOTo/eD1pj5giCRdWTu/4DptWp0zVxCaTkmtaUGUgJVfELn
MJnAoLy+qVTz6QYF0Bf0Dcy21asbhCSrqQ3BaR/GjNu7W3fRatkNc7MKrUTsQAkciChhewbqzfjA
ex2UUt0ZXW0QhyYzWaWsM118NdDEf6bVepfCZCnWYPv4Kf3A+EvToCQGIM+7UdtIaTzTo7W56LBC
nmsYWS53mJimwPHEI4/RvoCQOrrPEJOTYs29oUaQAT47wN3lcQ1fVFRsbCVvGtp8VcSt18Ec+kl7
S9+4NxD2KMoSIsNG+7AURnFLZfAp39dRRpe5ncingwzCvfxgXjcoWmisoCGJLv3niBohxiunVD1R
FWgAwHLzIbIXhvmzHvc8RXIX07nDr9Qc287CBrnzjS4JjXX0J8PhJ6M47DElIOwA2tYxwI8IP0+W
3m3VhU0IBqVON+3hnI5BRCeVz6TU0R7MyRkmN0MbdcFIXKHkIH+a/AJkU9Cvn5nHySBtu4wxK8Ms
GLNXg0VhCZNVdDsWTozfuM7c5koTBingrdQYHRGczwDmKE8e+KMn7XNmDUE/+HUBHqOYESKj2qIi
Q4fL/OJjGNE07ToMvz+xIksC51nlkHrQv7Z/HAjLbhublsfoqX4Au+ZR+FwrT+5t5VMg0l4Z6Nz6
bVD+rVTU/HDDiliRfa2++AU0Mgf6E3qO4V7UtjReadwgEZLBvWjegZ4CbSU2Yx5J/hM01dvvUO47
T3ENhtTTemYut8JbmxoGSVzN7N4fi0wlVBjRrem1vibaJ7tiSF179MAlnorBEpNBolEPIoILa/39
H5kKypQ0ECcZG/m75AV/3ztWzdc7dLtUYq7dVqfKFi8D8YGTLy7vS355t1iPBJGFhAoCJmAi9/gh
u1rKff8Uw4jMva1fTh3chMjD/MOsMoQ7iYAZ7bkNUq0aeI2ejWXoBkA3jpeYYTeRxG97Cnly/wZl
xeocd8ot+OHhzhORFOeD6NETSMW1wM+LWaFKUKSRwQO0GacY0Pck/MjBkjInUY3JEMGoOreAWShr
o7p0G0q8oer8q/nYmlY7qP8YZYFbInMz9485WCi4VkDTbYmuCoE5ixmd7ChemXY8dX+7JvrMWS2S
Gy2s/8mAUtKfKRB3xpoWwSOY8GhsDeWenmCh8y1Hv7W/bnsoKQYOBLuE7XM/odfBaXxp9TDUEVPf
XP5HmMxBU+rappe6RhrfDh7GGCKU+VSFZEPMINhRozr4ULa7uaQsu6xNUZRas2tB9+g5NTCz5fQW
IaxBb+3518u4BN2nzkr0RMRLeJVo+MWKEx9EoaD+j9n9mXfVguP9S1vRO966ypF+aHnFM6ZiZrYC
i6tC8uZ3qa/jxyITDom40NmSU+H2e5bd4JI2F0X9QktKRwMhvawozUaH0MGmdnwlNMVK1FXGUEg4
T+S1K6QLy6Jbq6APtTI1XsqJRNB3j1k37PZqVB7bPvt58XwjWNkGwODSmiyEW6BCr46PjNGh3BN8
Pc+WwT+y3l5BiSF7WtG79mIpKCXJw6g+za9Vr3m3oIKdSousVi4n9NaXg9mZpjJTICuMSQtlMw2O
3w46v+NleomvKHniEBmvp0iM4aWpZGeA1LP/+Lgtns0N7heTOoNs02/dwB4X7rcyGt16GX0R+XTn
aBgfiOov5le2uAZ+AJLeVjTk4Z7TIgOS8EmblR36rH8dB6r7eGCtnN9HgwrBgPYd8L83iRdxJlXp
Hk4OMCv1lfOR2fcNAK3zjPCckj8OFUR167DXz2eYB4PdcFMGzjNWkKHDdHBaQRzSM/fY+FIiCnvY
1/8I5Q28svF3/9yGKef8RwTiJe1M1swqSt4kfgFSjI9Kc+bcpneLdkNgVXf7i6cZYq/+6073iYZ0
w4QtwCwFXt26Ah8nbJrHeqxOi50ZnZWiyfUpdZYmVFHpO683G31m2dg0X8olUP+PckjNu/5vQic6
EW79Q+ECnnxC7/cDnR5oXH/1/5jEHi4gMAcL3FgA8pgukiMjvm2DLRkGXRZqsO0PcJq+r1wKZEr0
UR9ahan7nK12+mm4EUIdPfF1PR3yBDPJdbUvPCkzQHlfgYaspbAfFNgV9NZEag/loWFqdov9SLHg
ovjbAqLbebjNkMu3DmGrPUookvwzcJ2ts7vMyDDm7WgNHu28Uy2e7JwLTNFdwrRBPt5u6C01Xb7C
kKgS124UgBDEQOTwF+stad98O5s3n1HVxGG3UW7mOvGwU2NWSRGl6sam5gmj2GLiWlwdh2OjUt27
J9gc/csewI5flNr6Cp5MK53kDeIWHtPtpHDawmYk21IPBiW7aMSa55OL4/5Sc/9eulw94BZaTfe2
NzLR/d9lOnRwkMoJjCqGctDJ5fpV4denyVp6+8VzApwhtXud96rpK/GrNrKqvydyICzMLT62yXw1
TJ8KWkLn84t3R/vGGOUJy8oEV8s0WuG9NQ9hQXyFIpptVguNz+2ctJsMS5qOxmA7nubRs59HL7mn
2hN6QePn73KKky15g7AXlHhY9SMN+Fa39PAqI1Q8rqPpHF9Qf6iskxBStJaOPeNoxB1Ba/mYlubm
N9m4gK32oz8qegZi1YL3GjSfsvmMrqtfWP/a5cB+LX5ZkfaDYvC4Nw4A/VSDR2eyeWhAKwPRO6Oz
PHC+ZdilRUMqlO55+PEeA9dLfgMfqb2xFziqI/xopt6RHMlkLh44h6tTP7UG8ToaPij7mnzbCISR
87kfUf4EwkyssPY1HJrplAra8i61lMQwJO8BeqpCj6IlkokT9WLmtC0nCVz+nWsygNVKiFoxhdIZ
yxqFcyejMPCHX15zxKh6UJJnSU4EyI3+99WJYsFZUYJEcb32zTNEUUCeCaCFCCw2OYzS+bvsanws
9JjeHCSl/kZEoEslvdcHFh7rYYxTqnATLEPyWty6c5CpBnPgpTHO1sihu1xbsxIFK4JpSIGhb4wF
OwBQzFeN3QrkzYaGc/q2cwsyIGX1WH8zM/eiX3mnsFLfOWmPfiZvTWj140gmpWdBJlPoGNq1zbYc
HagdGx84FvghWlJudKPLKokgKp+rnTDxmmy75XZw81bVmFclGZsamJhT/KHKjy2bf37M58AYXmxV
R9+GaP3oU5yTD1IRZVPTngCSbkdjXFdfkASRieUtu9DUG3jbXbk5NNeSOk0GzkDVLbxhqokGBQ8o
F6A15+KLiw2nJEE4doKiFMrAVdvW0tesc53BuusWPDXfymuGABRw+T4eS5DTVmpV4cO9+purJrrA
hutXU8LiHb+arJOTekec49s2Omq7sQjMbZ1lPeSCA69yMy3t/3I11isptp7DEzn1Ehcft0DN7WCU
OqVy5nXy1uEwUhFyOzTM3EetRY0/fyTywFiCEOgNaos/CHd/e9DoaqF9X0Am/2GpK4kZ573r2lep
UdhdDRPOfTH+NqMaR2AFkLwY76TFcrY+RsAaN3TicLYGnW7dWNgVzqEiKgaw9DGx+iEhPQag3iqV
bvfrozmymGzYoM00n70WUnrFJGWSfRgNyCGdYbwYnHWf9WrYlZ5CIPXe+k/vn27OIrc61jaN0u4L
LXe9iK4KsaiDxSZpmN34BPCOResVs/nSCTB9OhPeZlrMzco1TwcbidXCxIwRQnlxq+SeJ4Zcwo+f
zC1QrxMjJ8YtMzwYp0MpN471VWaR/u7L36EPcJVGPvPB35YYpG7KHegvR+dixVe6kUmK5SnZbCdJ
yv8gXcUl8ZaNvAD2pNkxh6lUpwirb8SSzTafoIfvb/iUTiR1iEEJp69daOGt+7bvRUiPsA+3pIKK
FEIa4xp7NTjBUrjn8FK1Bjw1KQ9PFZc+GUmO63WFBceixd4/nb5d2V7uG9cj/dkrkE1y02uVPqPg
GvQ0k2GzCCsxbrhzdcxhqiKg9JVPsCxnEEMcAPYhE+8LtsYR9kkocr1Vig7910qV6nczzBGu50Na
W0RN659cxbLN0V7sR6Wua5lrjJfJxjB68PIV3SzyAxLnbXiBTlIGb3UmSQSYWqOc6mc/EVbTPHTH
TJ+CoXYD4pqFeDYbrI3LdRGwaxmJNdSjz8BrIjmB2p57GTBF0InOlNmXGTigt6Cjktbj/CGO5uBa
t5DlaHUG1iKph9rFucINTeDBrLcYF8rOGEa0mBAzQOV22jTteUUEMQAgHC6HN17gc829UnfaBeNM
fljaTuBvpyra+UW57bFUGCKEcaHlg8R6taWSyKT1cQQRPgzzFUv9BrCNncLyreMAWS7FrI55hRRP
aoW155KsntBWE6RZQ9lQVUEkne50fXrWmiVGAGUlTU5PQ+L0zC1fx3pu3aZriM2IlH/ZJAY/eSGs
WUmMoRL/mUXDV7GXyqofJ7sGDqpgDXsuqAtULbAUE7C3Pgh2VjcrkaNdCYRvfkexchVJKDLdP5fg
08AeCPCGP3gEzleWWkiyHKPiLJRbFob1KA8TZuD7A5pNkBKfpDkHX0gt7jzsplLBRiguxpyN6X8z
XtgYKZPKJMEXHj1QPAqFkekQF2DlnVnH/xixNBNMYVkU1vPIYem45Rd6u+AgyG7dPOdXbASTMko1
nJ+9FjiyZN3zD7BJlPWBL1GI3xeqg/oV1xUFIJ6WezdG3FD2GP4BBXb037ik4we+J699dTp7ITLb
Q8vPbLliraxuC6jS9344MUsS+I6D/6EsMW5+5aqF0MODkczOFPBVmzMXENMenKMSjTQvR7HYW1Je
0O42UKfyeWPXubYfDf2mdzZYlzK55y/a6yD24L4JRlOzjigzuHYHSTUBWBS2eUFy7tpJ/dHvKDAn
na+7AGI7NVzDMHqKjySabd6tPSIvKgkbbP57Ms4fQ9AW1UCQNeLKpmIPxrZuILgGtemj/2c6CFDP
cdbQM2nO4S8/PhbCxbHZ4BDnqcPAtNLPgyayicmmxs3ksl1C6JydnNpBrm6NB7Nkl2fUQMfa0C8l
yjQ2bEkxiKPaQuR62H/KRGsU1frkqZPKmTyx+zLCWpzXRy/rL6Fbf7vOWakGtAhNE80zJLdSjq/S
E90gji1eBNatp3OoSlbJpimkMyEv040kTOo9RIFR8RyqOfiF3yVi9ZJ+Kk+/dcGN9kUmpXSVmvhN
+8+6sW23TNvFCkGN1rrFL6E2xj7Iz7i0+fJ0r6SUJyEy5iPW2/eB7YQHk+ddYbdvXIRYFyOat3sp
BWV9Y4d2YyLmNZC2J9i92nmsynw69WsxMTtZe02r9xwdXY+hGzrtfG1g7MRaysJjjSUa+EFAsnx2
cT3f0ApYKC6zk0ZZvDqQzQKCx/MB/ecqOVDfhx+x5gxhZWmZPZKyQFniFKMXhwWc++Fm1YwujMT8
HtbMMw9AcZKf3VIqAoiRDxA5h6hq5O2Hhy2/XsZEm+R8mNG84O9xsEityn4Ql0XSUxpO+V2vxmkX
I19sJVTCLNb6jNa+GAkHiNQmu/dQDlxbpJMsm5Zz6At6mKw7V64CKA04TKyzl/QVACB0yncu8KAE
0GJ57RoFdu30w90ke9thbYpdgAbe/SS9r8xGux+DxGwtE0NEFYpvInex70LY4hdDx1WWW5FbhTCF
i3ZesX8ub/TUMQ0kVqPsmFIfF/ZWVNYd0kdZgO+Bk9hX48ZS7/F4xs/58CexYhelQdtHqQPXR0v3
9vHCowgllMkOp5Z/I0XJs14rqVjvufKi0cGII2KS/KSO+Wf5DvPlNBiEyGkA+LYGl9XtnjJA9RxA
Ervn0GOH7BxRWeOTQrOZbExJfrBIbkt7d27lq1xDxnBb9WIGf9MjoYlQ7Tvzho9kgH5Ot6jcm5x9
CVPEyFbDlywIFx3w8S7ux5r2ihRw7Qjk0wl4o4U6oeFPkBFTRJIh/bkKo9/j2ayHK3wO8B0hR2D1
w5SHaGTLhWxoEIRlI9WxA+wd6hFHiLZxPNDK9aqV2hjNOZNZf0RrY87kNrmySN0PZNVbtqgbIQ41
3XxPHNW/ZJKuRCIitU2dqFkkJ3Gd3DZYEIAygE5GC6dvAA7uYpCHmHB0QwhZZHmeVvctKf772+Tx
F3b/8WMxs1xda6WdaGLW4CBwaXqeox+XQ5ukgeWUjvdePI6HF/+1x5GcQKf4PayzsyTYUGdLH413
JsmzNRYNpACTvpkTi7KIHXNu47S7cHSTA+TPxcZPc+/DPHmzFq6K8d7SbrctC27MIUV0dtR9XPDr
D4ZeoFLXMkIO8aFHjZeFOieUP3KcEFk6EhUXgWf2SwfRHPYZt8pjPoWZkJU3ht69KkD6s8bz+MWu
r+pU8aIf4JRl9DhmmonTskN/brF2oR27L+kpwSgVmniZiWkVI325RLcxvzNpwyLKG+Y7ltP6luU8
xGLCSHt4a8N/WbSc9uiH5XTRDmKHEqivtBSPzQE5WXQT588rK+Aj+kQa10KMX7/8smXlKqbGsqqB
3P3m6Ni+876Ryh5QY+xKMNZ+FN4kf4VFpDFJ8Fm37IWsfk8pIwCyYxwl6YSKxwfh4U5xjq1u2lCP
5NVvmqDSAbbLlmf97/amNwvff08SQVruERFEmep3Rzci1ckNSb45uujvODNDU/C06+NQ8q/arhgJ
83uQoysVYGFNOO1nJ2pKxXmSRXIYRdyeb7sWpTm6XKJwytFswxmUr9nAfQnyHH+7DCb2Nlxv2Vzf
20m56u5gGU9Sj8ssakzOWC1QU1DGLB82PiXI3LDP95z0xlP5FS1bjGc07xpCI5141D5gWTUwyOw3
SdqEPClVNxqetrxpjzaTbp3oYBDKY7A/t+G4YGgjWulE0OQ7fcYrPZyVnVrTxy/6+YsCnxRgcHH0
GrMw3dtwsBxAmLTOPSZiXuD+uZLR3vum8XI9u70BErUBKeovEJwwhCtOtsvMb01acaJ9jjpYTL7z
IP/Gy34fINxgb24G0goqRem66SLnVRul0/ETwrYGq9iDKT6Mfle+gBWeWMiEpWhVTTFyKc2C33NK
lYnLTy8DHthTRxh7Hclx2tIAUFXOsx1Y0k1Ix7vS7K8IgN+M2DN48OHLnM65NygOXpTCTS5BpRkB
Wtj59zOqXCGxV5yOY5wkXdUWBS0KBadug9kTT3evHNOIkJ2M2TuqTEQKvIewteNE12eeYYbbqy7V
8RH7Y43OG+tStcA1sKdpsyus+7+Oprno0CP6CfvggdPhDc/EBMmhCU3spCS+9hfZ+Q3uDL5iYwFo
f9dNf4S3WVP5zMQtsstOPCWFVkdonGl/dbDLvMUX0WT9QlZsdUlhLQ2ifjDvlTKdDs6+rqfXhaPQ
0gmbgfjdbcbiUQ6PjQu01Vmpbr0xSpKnfi0aF648q/IEWn318khTNKT3w/evNStu/31ACOx8vPZf
jbCnUWLYNRf+RM1g3/1ZJMjKXPK79JFMSw0vqieboUpSkIul+/PcToZa6UaGO44S74QZ9Qam84z3
HEjcgvEqqwI3oJzJ3n2XG3hOOL+bPk9et/+QEBIbdB0efhd5joso5b1w9JhFR1q6IOG6Qxia8IJz
IYcMTfTxt/hqRqbxaR0+JASh8wKHc8TuPSOMIJgp3N/HXmFbaSJ2yEwCF5HFznh7ResDrB7ibTZa
RLn9j/A/so+SVOtCWoMSlnb9SQis3SQcVBu7s8e8pceZ91adP7cvNW2ILF+xoSuciwkxJzAxd2bh
KPhDQIOwGdW3VNp41nN46RW0r42f9hFxGnp9w548G5Z25ADwnO2bYmCTtuaxC3JADS0lJJH8VR3o
+MYgsor9bvx37MISrBeu8uotsfF0Ohk0jb3bn8zzKdvBlMrFv6jYw4/Ec0jqR0CSpxVIZuGKgRDY
CuzEz1gglT4uM8CK4fs7mTjts6+ZnT9i5YYs4L6f3T6A6aIfKrNubS9k3FlKudfKbApMAVuKyZ8y
RqYWAq1nPF7s2UOcYgINBbrOS3inU4Uq2u1MYAM+/2hIL3r06OwxA4aIkHPhq2XgPhWUikYXeOj9
x+/s3LGhMubP2LFH5hFib2n5ctwvspc3Ozjj0wqJNLXWPKJkjQWKiiQsA4OJaMiWmJX/3xBg84XB
ya2jDXeBp5gJbkb/2LIOKcuBZhObHGdvr69doMMlPr+7JLCjm2YIn0NQdKqFLw71vrlMxoM/piVH
hkL1zSkkhLoMHFWmivjQ7PZGMGuP1P1oVBWBWa5McumwVgGo63ne++afyWDw0jmUjlzdqLYuCyua
s8j1Gqq5rw/cbVRTSnD5tgkjTnWLpr8Yp9XksaiRdLhacE/ca2552jSDYB4BiJMkQnPzZiV82ToE
NN/D/6EOOQoEPCitr+weKbsLrtexD6RGr9tyEZJK2fejU0WF8/Br+agpwmiXzd6eSMiF58LPaJ69
WtGWRFdrThoW0rI3tpW231kRsSTxzAhVn0wTJ+vwkVcNpVpzQf/rFTtZnnM8XqSB2QWbJIaIe62N
RGYtWY+YrZ/+tHREO/8Lio2W2bfzEsU63m45MJ69RUXNCBkkS5VJJptEKG+/SHe06TmTyAn2dv9x
Jp44pOda2xW+KdXbitCaD7j9UI9l1gBIAnMZzRHqnYjtEs2tLSj4vZZgdJ0jBsTDMHkde3Cb3VvC
xOZNMcppBAhOcc61X/1AuRcHUdtbGb7r7efbmiXANe2JFoV71cv9Q6tWVedEnFqlaVPuTIUwpWG2
iMlrip1xpmBMOG3N6Bpf6PxfxxJ4DZ+Tvt0cZ3x8i+KGRGB+X/6jpXXxCUpSlxt4aW2+qHfeTsp0
5sRFbNXJlOxG5nKRUMmCPl5MuMW8Jor3BQUUkZ7uOZcKotsk2npAGvB/xur3X1BBEx4wx0O6A8Sl
fXwmXlSAerIeosN7K4jgcGe/rHStbmrpYVRNK4TE8mOzK3P2H8UQE9JpMtO835D3Nx+NBiFAvOxq
fFciq7xLt38En9B7KXGg7fP15/1WXJi1Vo+rJEe6kQpCF4w65uEGYFWEIWoPxUCCxsHgeIobX4R4
PdQ9RqlCxGkqRfEQ4LuyQT2elLzbrsO9vreSMxpkjo1034KDa+pZQIAdQAL+JHUCZU5hXMkOiyAE
TtfrT3wMq8fYGfwvujc5AjwZbiyqUaFKiZxHy1mTjJZ+49JpNCfP8UQcAFkrirbTtFY9MIlw/7jc
PG5KZm9xEWNNBphqN2cgFjH8NgCLXNjnO1g8t0s+qXIooai5cs+fj9y0ev4z+ALfc+KF+a6eOX6+
LV4yF4G3ACk3eOhmsa+mNdxC61k1jFefK8zKMYqUxyRBz/i76A4kOUKopL6iHqBkENzNSuxPEwu5
so/Ze66LzNdjCNRC3AI8WfzXhPCPT2ABpos5N5gOJzM8PvQuPY0rR7utFEj2+Eyxfx6ANGMUx2WM
RpZOsyMamt63AZkn4G4lzNZNyC3NKWbxVHPZYDE+LnXX+2hw6NIh9Sx/+RlJpEnAgF69F+hT/AMG
5W8v2T9uHQZoKOTEvIgwHSA5ICUqTJvYUgB/RFHqXuKjSCngcaoDLgIF/jgjOeoLV6WNRtgJaEt8
97sdATo9h7cEce2Ll+PD8rqanhLsFwbZAO5tK2NW/F0Emdj0KTDaiYthVjmC720xda/EnIIQw+A6
Q+d9tcnJRyF9QMvRbASqNRSGVsD3bt3dR4eu42lzCH1LR59eXYKcIEaIjv4ejxsr5KCFQq4FI/Pa
g0NuvW8EMwDpHpWsj9XGT1SHakkAoRFoke5eL3shQc4ILY4wDIsQabDgqQjmGFg9ci7wIy6na06p
Aus5vr1mUuy0C8mZPo78THezBgwQdITE7yC36x2BoJGxJCKG7SJ9sFh3XykCsE9vY5Ogs3apDmyL
zh/TBejoLKsm0JW1DAXTaSo7TSJFGrJGPgY2gxAraSmvwUWcwVroNfIzmSprboeqhgE3t1RZG5m+
DpfTMk0iIRM/UmQE8NbQ1hvxOmLflteUorCjoJdcFBfTqdgH6GKRo/QVzpIFvnmKQmuldvKD+mI5
kg51rRa882/shd/7NJ3nYo7yUyryG2z/KxoNV5aihFhkRvy20fALOXJsq6hY9/Cn3MPXtYONJfoe
OQWd9K3gbKr5IPFv3xNQAtvJODv48yLpkEIrYNNETFhZBgEi7I2Br/hyzL9LS/Vazz/YTv15L3Xs
oJiwRtuQvVQN63Z8dZZCUXyX43NDEoQjlhasZ4TH/yWPB8ARiNsbvKFoXdfj0O79KvSbzBBzNziE
Gne0KU0Y60ExPZe/eyECmu+eiHV5cTmOSTTjbAmhuizXAoXrFnqgjRGV82tKIc2IyYJYPVWsCo5N
ThN1TmZ5v8lOiSsd7/a4me7XtAunTAY7JplewX0d8j127KyPPD6f2g4ZiRpoaMjyHkozjfPIw+sn
afXAn1sCtMdke9cXEDX66yfvCEoK4/I8iGh87FfWRKwrMusimH8TMR3ah+CQ8+VCDMreU5JM07lU
gU2T3v6E+eKgS785P2imW5Ti6gmVx7+GW9mDt3O5Shj49yIBzkxWr8+Eorx3dqztzuvcPEYM4B9r
Ia7/ZtrE6TkXMuiSGhNznr3ZXjMHTuEIpLOTDMujpMlaP+SD/EjUaWR7ixbVhrSbNfdSO1rhYpMs
OZnT+exwwwbvi5JGH0sRUJx0EFGzchzCTYPGHjSuyYRfxg4+vaqO7l5POcgeqxZBBr8x3tRr+rrJ
KkDjyHX5CsQitVgewZj65DkpHP0iv2TS8tPcCjjeBt7aKTOzno/Vf5qxOMUmUEQGilVcQXsguZ2e
8cr9d1Mdh8bCgMo6YNCn14e+4JqElVGHufVqLOm4/bTHc85euh0CT4GoQsksIRyRIjh9DcenxF2x
vQQdixrC91wFJfJeyZQ4iCXwSLjyVdz5aAAvy0bWzYaRd4AKsZKWQaCCytRIsgwWcXDM+nzXRJ85
qI07fS/xORBnjAG/l3GcjjiGvLXllVBb/4vhH++1o2E8jfRTOY8QFpDQ+z0PJR3Z/ad0Gi2EOF88
zlKIYrcSVEsPmZiB61+hDl+AJAMlJuaAKARN+xshJJ4xuAtGlnIFMxg6/PkHQ+c6hXDTolVqZAyL
DnjbDzrJ7c69oG6Z8e7Jny8KLLAaT797Dz4ji8D3JNY9z4aPtjK5tJczlTnu2oD0nEBivlnHqO4T
d45kWXUvXfPuhQ1dTFfOXcU8005/gdAdvXbFMWJD9cLX9SwM0C9LInlS6R5svSOAi7A8yUahBa0z
D+MvVhKLOFZadZbQksOomjlTOTN3h2I7bmIfC/fS3f99RIMqyZ2gUylrU+zH7KanAdTongvORraK
HfE/6YDoci5xVYc6AyF2nO3TH+Ig3XciqjXrn83nVZrTAxytmblAudw1hTUiUhCUDJb33Y3x6nQA
5pje0z4e1YyJDEngDpyTiiUODlT2eIjfFfqS2rNhVM+NTWKQGaPhs2i5VF4H+3u2RzuQ8musnSFB
keOt1/Z8+cQLEpIBr7leqH00dLqqx0T7hWkEL/EL9r0TJdvVR7kJPOHYVYuEefjmGTTSD8Fxlv0M
NoSWsTUjAvTJM+jvBiC2FgHk4Whp/aOr4KjOhdAjCTQ7IYcxTFDtoECepZH4371Sr395VpfpEwq5
Rzw1ZYLoNTDJRfEmDbMN4VFdfdPJfVkujsCQRK2RsyG0BBoeb+hWFhYPeDbpYipt/JDnmAfiOJ24
AlKfHCrbRtfT3C/wvWc1wruDXRZPNibO1+u9VHJ1QanBquNjATxb5Ar2Y19HEXW3dvGh15zIOh7h
QFh/ajLKmkxGYyZPuj9thdT3l3WTR55ZDA2IIML+a6LDoO+cBgvvTIWmCL5+dEgr2XAtxqEvgLFl
FPBQklUptm287nFOFyw9qEhU4rz0BwRZkxSBrl3MhtgR4j5fXBVHmdHfe5Vgkmrkd1zCDMePRo+c
wyevcr8rnQqE/dH6KwMm9uIpyzShJBFu9nuAMXhOXswvMErBTnEW/yNnYB6l4/GhUzP9hikEO3WM
pMnGtofRHrwJbo4IH2BX7hQGBaSNVzKbVcuNkBuwbsFWHwifg7j4GpnYgE9n6EAmC+s3Be3oQj0T
Dqk0Ofuzxai0hRCW/64/98zBkzNMs+j68wXfCpnIzdWPpVRDdBUPp9lAZ/VqNIQVAIrUueozr3AA
d/QpRnlcPCA1StGMxfA/bKzuVf2yZZ2QnQ+sD5PqNAAUjH2SBZVgWDjuiKnFHrGDlXX/XDv04rBE
speCnPLngWXA8BLKzJlNX+RyDJz899mIq9Lb0E/y7X25UVKgW2baXdABw63+mL6j5k153bC4ALVU
FqR9NntYjg57urOXqOEvKXC3DvuFeUZYMC+KjmCHhr6CrK+ZuTenjAmx2uKvBrf1pC/kKDu3MQWY
+H+9DoMQ5NZMnyDGeyW8DorqzMTBE4zxS1G6EYJCgZP6a1m+z2RkZSHB5UdQNvlFYmOC6NOXiv09
Pay5e3cdxrPuQZBNkkIyD3/1yKIwYIjQeZp7HH70hQLTjtt1VJhWIbLTSfGjj4vdRq9FfZAFKVxb
7VJJ4TNWgrHjtGqdC474LULOwdOZAvFDMO2UglgErrgBZrqhaPrBSU7eibjn5tcWvuK2rNjoc91P
xhtWiDcCGN3HbYc+PuAqMSdPsLom6S6pHmY7Oc6vcpCx9E14L5u4mNg/nPqj5qlKqZVvFD9g+gEv
fzCnAuSW7BOPSuz3ZH0npwOrEMVi56lJJ7ZYLfIaGINFjgR3EackB+4tWSkwTrWR6ecS3XBAmkQB
T016fqu8l7CED0Njl1RWvIal/F9OIrY0v9/tR1xB4IT8lFaeCxGSSMyE6T4chvPZRito+R+nv5pH
4i8hY2v502+sNTro4zFGOWkjMcB22Afwtqt5i8Ieys89hYv6fTFvQULe9sbHF7fSCYA7p4JDg8bR
huTlt44wtljy/BGPNLL9Lu6LYyL4wRQt4D4o35L6EwdSPYgrYSqxrd+TSu9cvQAHoIEGYNrSm6fJ
tltgevjamfDAevIrDVPgJbyjXPTkIKy1XjSYJc4SpiCcQRzCW+BUR6hIqwOmp7La1UgkyIfuSoSA
aH1ErtWel7D0fHlv7KjdcRVOp7uionvP73LCOGFOBMkOv4Kk0UHTtBFvICRIdSTyqg0m3XkGXrK/
MdiCHkPDV6dAv7dv8TwtD9cbOfKNEsq5TvgOorD4sj2VEGKWO5iFUCWBGmxjctJTXecHDy6IprLm
w2it37EnF/Xq8CgixMxZ6I2rFvguuz6KtO+Ev+OwcApksCjZOpzOHF/o6T8UrnJr+2dMyl42lbIg
9gOfVo+frW4Y+uAUEyvtCnuqDbXq0xQJ5Hv1Vnv7gm5hTnydm1KPZC5YR1Jf77scAtbAnZsh+YVa
xOyZ9vUSGQd8cXnQpnmxmkAkQn95KTi7DUD5fSAxgtvQ87HJsPDe1W/vBOhXwG961/+5a1us69Dm
ePZC//k+UXRZRrAHa/cVpDe8X7QDlCxwXI7hV89VhvShuVbjFvF7vDWixkwZ0u0pIEJST0ZffZqv
8MgNffWlFxn/w3xkeuKhZTBxXgKCu9dIdW7w5cwcISnOfESfJLsDoCTLxz8pgd14d/0Vj08T4sL6
GAhqTNad7L4In3FLm5MuMzqqa+pJrCdHwglKJiOb52YrsteJfGG9p8Ofu8SIc/MVPv6eq6E3u/xN
z10mojO8rkIwQ/KrWaaI0wslQLJ7zyMThLRTVmUlQnJDRSzhU0UqwdHM4WHdCnDH1DZcM94aqNaq
5BtA3bK8d7HCV3YxdzC04R6IIsEaOE2IEmWPCdVLtOaBmQOe8YaFRKs5pBzyT6C5aH3MISczkTov
lFc6iCkko8janH/Tof+x05Wa8eBdu3Ip/tIYyjGLIybt7UBElEgi5gFmPV+lWAIGctZSE4o43GeS
NnRwIueTDFTwjLX5twAe8pTtAw/8sICGO4a69veZenH1tkehtJT2d1zpQIINnuunYwFYOLCIZQ/l
55qRlK8Dmp9j3yIGXXAspMcUXMN40cH2+xBAc2Go43q5yJKYSRDHvovkpcpawiNrBHWPdxGK6TMW
+iqXLYIhiJCHcyi8Xgos1S8ahjs54+rg7BtLQ5xMPz/3hCTohVYuMWIgJaowu8HxxJ6ywYIGQjK1
32GzMWCoD4vUTJS+7FrLQlvM4u3ky2a2F/Ad5ozcvS50SeRp0VVKVVkkbn3xl/wYXAQ1rJvh3sBc
cSdBE5mKk+CdUE01fZD60LtyezLXtISJJiGxd3mDnSxrHAS1o0ofUwjA2mJekHMomA/3jJ+fuC5P
qBXci40Yar3tiO4WdAzofDXkTc6nCBBgJp79ttS5su2246vaP9m/V54DTQkErr4Dor13GBDq4qro
vT+mbfhaNLCqpwNZmt+UYYPBUWoYguldMSG6obDr+5VxD8qek17fnHygJNyDSgdjiNiuXLdKYywt
uW874rmVkAiOrJVzNPoO0HkgfDkvT4s4N9L45cJyWSYlqVGhh8uy9JJqDcCGdTKWxmwAXSh+vJRd
/PuCaN2rlnRnVUmN/x1y6fPC8Eh+4N05E4vrEjbu8FxxbBHI06S2IiFM9f66m4wNuXSyJxeQX2wq
nGSdw7Yeln22Wxt2n/z2UwbQ/ghzjV7Lo7ilm573nsepF4zZpiyKaknPbgBvJqoWnqI9zFb7atLN
AVx+iccBefr5lGLUfLKWcJTsE3kGEc0zyHQce9FPk/jywqPUmiTOr2KQCpxyYFEIAmesd/IccOd+
Z0MLT4T0pDBm8662tVLfdGYfp9V+4IG2nP9FbyMghxbnCbMbJ4SxP/tVDuiPQbhEEt9IZo7Z+IkA
fDu0dX/MvDGetNMyTo1pSV+B8nun8v3Gunbn2M1xkKK5TZ2nt477AURyFrCwy4mjhYiiwbtTzV5g
bai0kk6colLhC0xL6blgZrmJylaKQa31WI+TNr8isLN6A20Jde6j5FXTTXDEiZ6k6eYavcjIntDv
iNtqJiph3SklP7hWW1NhbQuRWOo8gKxvkyycmecNy4q4+yja49C71kYUnmuxstqLfiQiYQnMamYG
wnCjqzrosbxEz/4KbNbCcQ21X1av3Oi1nn+2LOVvrIV3My89TO40ijGzAtLdBy8qO27jJ8TJbPNW
Ecw+OCVDPYKK5I2D/6mxj6+WTi/L1iMIgazB84c08CHd8wvGoN89VJI+04A1iecLxtwFNyjVPJQf
1FxeJUA6c+2fSVu6CZ069SDNOzTLvAmLhp9kpVwi9bwDed3LTjAv4y1bEXlg3em2dDOJNmwpopJe
UGxOwk9BR5Kw3XLPN74LLJUXrwnrcwl7hOCDg1w8ih+ZL8cpHAAYqDugtCbWBz1hYDS2Xae9/gZk
gEz2F4gZdIJQX6OsrAucQzRAf9IB774scaJJaCAet7hhknDZY3zG9XrJDMumoiIMwI0cyuJPqLk7
AR2hryTcsaaM4m6F/tinCUBNJhZ4JlJC52ageYC2TLZOW4nkT3Mrdg0hlgIEhuXUDlzL6tb+46wW
hhQ22B7nQUsZhYlaqKpo+MpKbF52xP/DZs0IqTZ9Cj0G7cS4d+DlcuPoZS0BUNiHAdGdAcAXe3HG
Xl5UI6xxnE5iVMohc5vLk/Gz4gxx8r1I7w5IMmhmaAN87qGT6qe1q8RL0XQOJhsrPlZtNrixU+T1
aeGPyl+RgPqK4jAYGzTkMuxmiWtbVxvEdIa8bmu0CW4srvaFZNcOIAMqHoLJ4sYjmnN2GHSHZflH
pFkU2p4B7v5tTxmuUsMJSyfeE9vhLgBhMspP5RcckblpqI76RQNrxuSY++Ye7Y+FtP05IzIgWbSV
IPgXZ7sumren+aXgTyjMCyhJergNxo/Gb0XOnZcY7DJ9R3e/A/OzP7rcvI2b3g+XL9EK3m2Mbw7x
VBSJ6x5aS+rhtWaXcUWntP9zdwXty1dvDqgLF7NzgV4/9K+JbrTgeeuKwE+3vt2IqKb9kAD/mnz3
nPUE23T4WAyPDlMR/d8amnIORLTCrTtOg7rEzIeHktiiQ4cyrrInj58Chd4Cp8yjEF6Aqrvu9gRE
5wNJyNjpJgTnSXKA5l4t2xakgIvFazrkTUpaRtc/3n7re6+qhb1f6tpRtCeLRfnAvrBPTFwyHeRr
32D1MUAXQW0hvTiPGrRguT16SPPT9uVgJ6Do0YhrkwHmAI6WZ3M/9RO3rMrzKv7nzyZ3TaA0Xf3Q
aNJazycm/LI4X3xgpGBeBqiA+PAlyMWUmGd5cVYot+Qjd86fEOELV3Vz9ihrYcOLcIuHVS3vdtQy
gB0Ftf8p0ddUuTbqDpEQI5jJR7359HgIECee0l7+gJspDlh4jrNsz5g0MT+ICEKMnjlQKLvvhosp
Noo3c8PJrNokFMrPlMjUVT1rRgmlbFUuZm4I/drxnVNS8ET7L6obUoIHISRwDI5FJAUPAc9gQrUn
NlFQryvzpsVH7aoHF/K6LVPZyWQOmFw4SXzCIHOd1sHMw4ZF/F7jFdaAqp3KyH2CzeyRHYMqgNg3
IX1+r/UIBLyXCNG1Tl63UhaTulmvcPbhvyx+vGB+FVcj/a45fWyDWjjUZF3YinSQWAIRJxdW8wKW
XI/IlpKpBX7IDcvEyr4Pm2yySgxc9MjYnufCjcF4N8wi8pybmIGj4mgKF02MBCWDGKFN5HBJryxj
VD3UPCWc9HcCkTUgswUIE2BsMD5QLZUaOhSsJn0w7GFpBJQ4ZZyxx7jfqGv3on9dkseT4W0w/Uz5
4T2EiQcowONGC/CGl7s2zeQitK9KZ6K72JRKt5zST7U9MiQj907MdDhG9eTeaEYWbhI/v7VgNXz4
MMUiF4/cjMwHyA4EZrw8xeRxiCh8zWxYnX104e5gOGMT6QputS8B88mmnnDEXN4PA9nfFkgSX13C
r3wuSAXmNyshMokkcnChlUqdZ426yfjmfeVBF6V0B0tseqoO2q0Ymf+8rtTJvasj89DvshRw5+YC
Mul8TDxS0Qkyp3AmOAbPezY6q+3PXMjCeeb46bfTrpzDz2kTo4VRqeUnZY87GG6KL376yaTSj6iU
1aHk7wnaurJ2sRrQRBon4PiR0NE2ikD0w8+2CV1HDuKYovF7ejMdsjCt3HXQsef3IsawHUSoS0lU
ohif7q/qlOvc3S+Cgq1DTzlnPEJLyEY6t2MToFRCJOzrGt1y5TpxnyQt6KyG9wJ1vCySNmz73RzA
eC5lv+CItdUvsL8B146h8jaWFyAXfaq2I/wzEgEixDPSmCpFtQl0V8nW0e1nu6cZ55SU70dsXixF
WVsmKHXNECtwuHzRjSxa8HtYFLOKCC801s+jp6a0LRNaG+ui1/tNN4HsCnE3AJmmMPhokAc5rYVT
5JLe0bDkmM5LcwY0Ryu4IvFAUCj9pprHJh4uRuEMBZEDmmGpTdFdaLoeIz+Ziim3II2yMF41ECcl
dwNNF/dPb+CtLEpEs9yiwLJUufUumOPDP9Hzp/65kHzRO0gYZoveQLxnaVGYstdQiVhcOx1PGgnN
O1jCYEs7FZMFf7hpdm705I0OtdZgqCMjTegKZo31S9H6WVvcGkL708jiMEIL8l9YLDXaMQC670Hn
UMvuikG5pwbH+vT5Mb1pocSP2KsVpXGqG7a9tMhbVL3bXAPlOOK8lD7vAede/v5tajMyMOeSUH47
CdnIAv9bDRYIx2nirf1XMskDEQJi4hoVPpymEDgkXtvbL5KqDEQMJm4dARy6PTWKsoFFKGWItRaL
kYVQyrhSersYHKndcNIsnoE4bYdagrnh8rUxut9omxzRXImS0DL6f0E/CkSVRfCKAQAO+beHYC0Y
mBHxCaHgQcHAvXHdEcptnyxsKyygulqBL2khjgbB/3v1Rb57qNqUpqHKQxYsfVerH1kzt/TQ1iZe
G8IVlV0nGcyO9OnieID7digDO7scd/FRJeopGNt+qRolsBW3HgFtkLKoGVoAMkSkHa2rmvyODo2L
ao882I20L4G9q2j39xl2IpitgDIRo2eihP58LEtOUVECoHfNlmbCtvK06rzX+hgaPFvHs0+VYiSS
H6u64nS062duOHTyO2KzEljtzsidNVW6XiqD0OZhsiCqHlCOddGLtLygv0rA+FJbVRZ0CwQv5V7R
1BcjKXasQMX2v0k1qxkX/3YWoWJCTpqZeaqXLUWnVBKKwQNbvv2fvpWzeKM1SOpyAHjI7pj+qZoa
Yi/fFNbU0Sb+lPumbnyok95xgcf55WH3SbRdSBEmUK/38ugkkJt0oK+NjdDYZt/mMFOH/P1lwzTE
DpAcIsa6q4RsdZLhCuMoyXUk/uxmYOUfOJrRmNYO1ghWjHP64Jbv1I3xP4W3dq6VrFD4d/TUpRxD
gqbD3z+1CxXVrei6TW5f5d3Pef9DRta8fpapnVOt/+1XL1guBnLKq6WuMzRUCmSfZirwWaCQcG5w
Rlofc9ajEAkuDRkQIjXbAS+yFpC84aUY8pzsSjoFaDfvmCHWr+7kORT+3mT1TJIsD1Xe0CnshzrP
oF1h0T+++8XgUMS3wLDo7ZkGpNeBUP1po+OSK+MeAknnUVQdGF8hl5FItF566cnbljQhVILbCksZ
vWj8hfM5/twzkfuehRYgBe7qCh5zWv1SQcRHgGuO7v1/9AXk2YxAR9HodpZWuFCbsqS+EvLCbiHk
r3fS8iXc2V0IDBFqUBN+OmlFU+fYMuPr7SUWYo4WW+94RUW+UdFVdOnnJCC0Z1MJEcQPGuklb+ZX
ykjQL/6MwE+fUinbeefAsowoDLUfxJIXMOgwePqc12XjEprqX+FccWZv8X1MONkrOJ91l/Y2x0Gr
GNRCS5j5tzijjpZJq4xoQX3wWbwsnN2RP6F5yP0ufLSuXw+eHYhUDDOCYV6WteRW3892pL82SzOZ
Lz8XWLGWdA5yJqBr9b5i9J5N5qFbQxR9EDuMODO8XJ/Ma7wfiA8asG+lRhBTqXIdpFlqwvGu+Maz
A2Mt3WKw4rsj8I0WFJi7L3SGbt9S3qZD9o63XFytjziznmMxJyqA3FdsNNV+2burXcwe/A5Dv0zs
l7nWb4Pfx6+6Ns1BvvUaI6CVK5D7O411zZBeDIOcnJG/JLXl7V594n/ealqt3b8ZWAqtafLOmLtx
hPGUXDLl86m5dkEYi6Mwe+21gWizz7YDXNPrx3pUmVo5l6pa6fYgtWNa6xVOLjAWeQThBLYD3Nkv
S1z7vcJ6rJAWCyshYUM/onD9M5GLAXOiZ7cMOlVhs3iCQ3WrnRcrX4oc2brZO7gFy/vuep0/T5mF
WkRH7hSBLzVsSjgu2CpIRZgWqB/30ekL/9QkJuKgx5CODkSobzQQeSUv6TP84tgaxYxU+6R9o6TE
Esz9cjIC/QHCsm/9eFUTN08u1fvanwwYA2QqYpAO+6lZeM1QTg6G45o7OJG4EsMlMc+AwvwzHtCb
sZGSQM8XpROQVcdVG52sHx6/a083O3Bpidfh5g4gPlKDpI9cHJuwhyPMtYAQgrYsMErmOIpg4exx
8VA9Z/FZAlC6BaPs7NhvDRUaUWtEDtiBKge5jXddIw7OcyJbRhDXfODfEL4Qn+BtZT/NwEsf5Lup
23vZ7ugp8CDORbNNZVsNUnC3Y3IqrWfonKFxJ+ovNChQK9Y0vDpgYA5kS3TAwkP9Tav+aU6kx/6g
/HVc9FTy7Y097NqvIKcFgnpsGY+lD6TytPaK54Cxxuu1HJiXk+qc8xrYTmfU62PuIKtkmcS+4btc
6D/1QBKtiV7ztqukgtwZQcFM2ZmUCI+/6D7Ml/oYl0rSdHeSsMgqM42MbzCcRc9/EOeHgGil+oK4
7pH7TW8dwfi6t2s9DurnPuQNKl/hgz2Ic21foSC/bSQnKfpGih2AOhFa//Cn66MeIIwUAVlS9kGR
EiU3ofRgPl5KFzD+Cx0MZkw2DtZ1fJMeCH6eo2KOAG+DlIrV62SP1oPYxEDt4wezvqq9O2LUc4GS
bB3U9yJEdG/LNhSlv/VPIA7N85l8r2u1VdPOWYiR+AiyTDlc626rcvPcyAnHeES3ZkNHoZVDJCrw
mZ2dp0x1U7bvSc0N4SxTl4LeCPkpPKEkhBzggfGsREx+zR7D6pauZllMFzZqt/RLr7yenA24CCj9
K2+fRf8TpuY1F1g51ngBu7VZZ9JYD6sob/rWJLDeFbJPB4TJY9HS4yLKnGaixu8GspLQQop7cNRY
ljLgVlzwZYlakro8mYgUg4w+8ESmb5vrmU1UlXdUVP2zuCr7KvczWyNfm5DHgxsa0akZX3gPv95A
SDfDufBAvqExrdAzq2lxc47sDiq7GALNuTNhYLfYrHCWkkv64ZYyO3iLmg4jXK02alm3XbXC1Rkz
6wCZTsfV8KoMLP9R4si2duqq36V2qf6iYMvoNBsFbasLUrS2LAHjE1CIbWoyXucW5HpocPX5sbpY
vFCfsYCmzH3E5xAY4AES7D0kYqv0Iqjq2HMXPhJCUxu6i/fFatgl9S788l09af/L//c0tUJJv+Kv
tuQIy1KFoj0T2LJ4NXwWiysKEysCGCqgleHdQAdS0ay9ASGWxeCVBnkObdGcblrhUe9N0xQuSUUI
z4CLHzDrbxCePdLlpGAi80mo6e5r4SgX2us1TA3AEV/nGetV+5PI8O9E6QHUjHYOdFdkYdEsGu6M
V6JUKPzixS1W5j9TaDuZ408zKLSy/jclwqzpshwpJmsfUXSBMxfmuh0vk1ZmSw6//WxA7sMISQE/
WRwAFPgZXI9nFbEvdk8KjDOg4dNG5BK+8UrdlQuoLQqUkotx0NRIN2s9LFI6fGIwesM44m1JpYiY
dLikjsc7HBbr1IKloEzBnN2+K29SDb9H4h8A8pv6CRnHgL1kyko8nHdxyh6OfuqAOynw2cc3oj3t
EIG38BQ5KJVgtmDXgOeeTIyQGjrFPMJiwV1bSUs+5FEUQxlXBSxezFf4KHrk76hx/0swSzv1lT6d
XcVHBeo7R/1Oub6KNstz1Jxt4m9mohM1GsfBk27lX9oNOY4hLtK+pcU2n14dq9zcS6fKWM+IZTsz
+tLJBfA0pB1fibNXA8xm/1HeIuJ+qI+PYqBdkEEbCim0OUx4nLuGiIouEVZ+ZaA4BQU3B0MxovXt
4pKDgTAk3TB2Ig3wz39VDjqWNbHL789ockmFvK5vsLUHLN1Kb8z/LOWbgP7PkmbYCnUFIP0UKVrD
6QujiKuM2FD/E2/PLqzoCNjBuRDNZVyWW8KO4aXbOypSgjcpp8M0cN60vdsPN/eXObhVuW5L317U
dZE/a3u+zNUpLLGYGfrBt4H5P+rkCKUX7Pnez+ssRwaBmiRDOHPvDTEnLOCsEXk7gMD7U+C7ctCt
DeRtvgEgC7F6e9rwSWMKteFjoXgMoMBrXlxN7dHtNf14o6S16N91zrZ3w8DoMcr2JWG1L0B3Yfsu
f+8pF/NSPnl+NYTUuJLaxgWrtTxFk4FWyqCFwDno2Oq4AhTMYSau8OsX4+jnMGBSmCV7rIkcvx80
XAAUjwP6dbAAloRPGbJaOwC4rZzY5PDOyI22sFFVsDbdlvlqVp+vIdFJo4FSDOOl8A6v2ADvFf5A
5h5oFBDODeeWgt3TrNUUtV1UaeU2OZscDHPjTo6PeiCxHD6Jn2BB3DItgDWIjR9ld/hOeyJ+1fze
ZYMenUWvKPvh/m2d+4tsbqHsyXEaOUo6L8hIDD3MnDHNZhmeFOvzjAtlxrMmTPSSmu96hZ0MaCOC
QYN53YuQngnH08FkYJtuwnf0AQ5ZF7VuZG6wVOQbsJDKG2+8VwlIraJrH0GxjcK7jOcaz5NHcUrY
pEk3W4aqxFr8zbDC1EjyTESlm/Y68ibcYKo4GkHrNnrdh3zkYaooJjdCzz2OlxwLT/sUKQHl23Mw
9aolCtbRcbrE4Pj6RQs0vI9rhgryC294MeM/8SEVRWit0JGqNz5vlEnqijjb+83mKqUZ3gRymLK2
fME9OVKIKqDi392PvqtSQurxjqfF4znLJfIXwV8Eoc3U89Mf1o+NrwTA6YFWGble3+U1TUpdBxvB
bQGaHm6Kd6fR+YYqQqLi9bMGg70UEWSI0FS41X/uEfrYTPYndk45zI1b+MwwD/F8MuBRft1YDJc7
nQKJTUafF8fr1P2nyitMOjYX1hxr6nuA1kLn/XZXhnYQeFmwAzh5hmvgQ84SyHcNky3/PF/TilfV
sNe0k3sQEXOAMOmO1c1O+Wf875YVvrMVNIzIMRqG3jp3rJH/4hE2qCPnXbK9MTX0g6IKP3Bi7pzO
vjsAnZTR5ZK1UQKkEtZ3K6ZLrIIetvRmYdMWdyLXjdC7Btg2jDh82QHH8PevwZBEtIWN7AUnOKP7
vA3s2rjjNZKS8Ud6EPPiB+qri6BzPE5L1Hm3Wp6JRNOfnykZP3pcU1MRfPxPmSdi82NppxJtewa6
Tgu4uIgiZNI8Hsu8LXN0uosAQ7z+6M5PHqrOMBsPFJ69gh2AgF2Q9qNYt+fvWwhI1p00ZSDB5ZmV
ZSTCcCIwWWVxu5xn14OYGsPmE8/F9p4TPgEFRTCzU08PTsOX+LKINNuY4hBkraCG5HPtMG1VCuAN
SiasGVjydu2Jki1U9QmfqvF2U8y8YY7i6jUeJsUrfIa6zg2BbmmaI8khWoT6KGsVXDLAtlM8iTJ0
79L2paZs9ewBSNN+VjkejvazIOLOdUJE3Sxje+2hq+rpx9cHaQf5n7ItgrXm7u39cH/9prd2F0HZ
GAxPUxoLW/eUOVX0Q3UsuPG5GJN1jPknIpNeO/k9aFNAAtMz9Cwdu1nSOrNbXYKlY7Q7nsK0+fei
3/x7D0uGCyPWEIlKZwSKNTwsi3aI9hehRoExA3NEtuWnV+6oAL4VAk6Xm8BYIQ8v+XTfcOnVj0F6
8oV/pgPZTVC0d5mnxHxjvPQfe8870XghAkf9ilsLWDhx/kvFE38olH0KTUqVEoA3E34zaqxqAOyw
P2rXXqaTW/DzDsKZWHg7Jq+j0XhSq3n9PnDd1t+9sCE/k3fqFEwwRAAQIOUz7G7ChhFWacbeSVw4
aePOhzAue8k/klIuhZHK+izUwdVKm19gci6gE+TfnSX16ngrcEBulvuyPs6Lo2dOFLP0xWwqm/e6
8+umTiSoXZkkJ+ilJwjr1rTKbIOF4cYcpAznWTSAfeBg7PoDQPAULgCTvof7bpINSoR/dQOt0WoP
WhZnnG0mGlUBB+PvEcg+06JQGsCScYCUxa3X3rGPi8x1GUL8cIH6R743I3e/F9Um4neSDJGhdTom
fbXA9rt3Wv4dfHOnyBxZiXlu4rT+no637il66hFNqshNVrJdC1wxviU2cqJXGGDJAd/HP9B68kVo
mZVtu/YDqti+3Eff92C5nrzZTlplrCCVBAcSQ9/fAumFH0KKdponDpSjIOdjF0knI8z7PiO5g0+4
Ja3ArtL/Q2gw6uMAjCP+3C7FxL8lpuDMzvAHkpY6i2eLcXIhp1sC+i7b6hag4x810y/72YgeiQ23
nV2PD2TkBkkMurBVKmZNYxkNX42ZiB4AEuC3CWVS+gzlfWLBcrJw9Aq4pnmZ68by7Gwq/zP+7l88
gtArul5JZwpAE+UaKLDETy653TmzBoCQ3J0GCWGnaKN4/yTo+SFxOdnRn9wv1xlmWehLRSnNeJe+
WzauxOj6i+QFe5mitNDVMXQKW7CyoMXsQCwgGXbYgI8GHDNJI9XmdxMzG2z2Q2wWWMudyDgIZ7s3
K41V1+1lavd8nK3509cLxRgbRY9NC0UeHLZhR3slzTri1RckG4gdd6QRnBuMrmbqOYjhOuquH944
t0UPol7bF1qvoahA+mtnphTickdOhmxcojvUiVXnlvj5vPCGXIt6Wo1zUSuQA92L2xX6F8wuwcmb
tiO/VBaUYvaeTvktpTovNHhmVQ7Nns1WpkHSi5jUTB/bnQkA95gWKnkYd+TZrQC3SFCcAZuj4imW
Dgc9FivZOiCeEkTZUj2MjbeQfjxfWuPjq+CA6PEqFp8O30duPWguUxz7GUqYEvr+aAJFHdWfbS1y
+ffwendK35GQ0xSnycv7KSGjBiLCyvqMDJciR7ElVImo7dOHVyZTGyoCxYGLF+NwyYFc7Di3b/4A
1L/TKAEBhGHbzs0Tx34Txt9o9oyued9FqlMy+oyfDdVs5wFdTszWV6cduaw0sUDn/tevrj7JHLmH
yKGW9NBFplVLCNSNNkQ4Wi2T/gfwJjvsiNrTaGiBrSdOXnEy+gdh7qRT1GVRfZZEqI6DgGX29kKh
r7Wk8p6Hyjmhzzg7JFhVc9GXvWZ/kzEIUAx0i60PH7l4dEOSokfaYF9MjWyz+2dWOK5ANM+BW+pI
j2LyefR2tJvK5ecWahX2tiKAI8oOLeHrutqHZKAHkbXzZ63JugchJTSlysd/ADPESt24Wabnk8xn
aERCDFAP6bKK26/w7HrkF9L+tI+uzMafnp5qayweSk6ylY++ZlLvyJV7Mbgb2IIxDxy8xQ1/m+RY
J00ChVwYDbDloZ9uvW0exV7e0c77rwT7YjI1OK5lA+/LsmoLQPjrqtd5oDKIGFS7cb2nGEAeHd3+
Xv03s75MkOUfPpN7SDms0HHqFdM+HfmMVhiE63Q1E3abxmOguIFQCMMW8wEkL7GJF8IF/nasYkDK
1aRSSFX1ARAS0mlXimf4XH4jez4+eWWYqx0hGVZKwrkeIusUd1RYnaTRfQnJWiZSF4bS9uG5AUsk
+bILXDxLWIXk6yUCXoTyMU5Pqfjp/NS+ELw2kN5FwX/JdfOPiEh9HOToKw08+34WAeQAEWP7DPC4
4B1HUL/ozBXrPcgYRhuRdlYpNvbx3rmI0zdbA1JzPhdtAO/5smHKzCZJivzfpKQiydAjqf0j+VHS
UaTVQLS9s1Y8fqEHMLUnGZwn0orFhwsLBEaEZX/61Z9ZNHIhCVquW1f0ww7qNCNcdsl10s6J9mx6
RfiXCbZGdUoreqr79c54wctheEeAz6ZZZkjWaX7VPlMAmzCY8nqMASmpBQE7ima3YRCNyAg7S8aT
HyYoteEo5lGVNSJyeRYgEdk4VlO4gdumGm1HH87niU+jdXUwNeSNvIl9/P9xx277Or6fnLQYJ0CC
Wc2U7VdilYgkLSpldaJ4kBuhzDz8sgNg/UULJOWThkuMOmIo+4YkYq5A5QJgXbxn64I7LXlq3JTN
LJ86TKcs6ZdX9f9gCK8f6TKcDFEeO7Yicje9s2qteBtYaY+HfwA7de0zDPnduPviLfN+veZdPL61
PgiJhQOZbxwjRNAiWDmC+AkiRF80Fy0ZxMxEVkRGaQYSY5nXhNB5vUvuGIe89mOIcdeDapqseVdj
B1pQCum+Szpc1Ti65KreNCi9u3ehyksygSKQp7IRcft3lve221tIsGbraKB7pUOEChQVnv8tXjT2
6/XMApzXwx7jn8A3dgWHTev4WHkjkVEwoB726J7aA6CLSzMe0emVPou0vGKeXWXR0E7P6o7rJrYN
1IJ1GQ5mYcGKdDtWibazzv+A+IytwONzzwROK1SVDq/E60J7FQ0mN4Tk+EJslee2+zhVs+aSSuvi
rBoRyl4ovF96Gdb4aFPKn+Vp2mCZEGzOrIdF8+k1OgW0jNilK2V7g5Zs1XjOeFpTuJeVE84NUChh
8K1EYn/lMnp/FtceyaJRT008qNrH0PDZMbz8nTld/3KXdVG5JdcQFcyX+PK0gFHzfHa6cWEqA1YK
NzSUUHjbUtL5JoNQjsE5N58GUhjwzx9K8NLxIUyaRvDPVPYy98CTDEQcewxekWHB9bXup1VJQkHV
FICd1prM6zRA+H5WwCuONKAgHo2ldfUfSU5Ezn8OKhydQu5V1Rtpa881MkDj9kQM9i4tp+p+UBTK
Nm6+L2tsGEV0YfxmMCrOqjUpfKt/0Eh8fxYhUHT5LM4MDACCnBZR2M18ut0FOGtNPUWNyHFn6iEg
AFiTqpvgdHclQBktnLhRR048ikPM6R1rPWKtSsuR1Rfjb1CRTa86zHZWRLuVHDI5ajjc3xDVC4J9
IPEeOXODnMaRQI17JP9hCVjvITABMICbexeqJj/cRITEAnweUeDCCFNB50lergkVS8gCiyuVS2/n
4T55uD35L0zN13wum/vUtwffZdfhT2dfdv4m2NIRc44zWdR6as/YOiysYeOqpI9fA915Qtyv2cxp
kUV4/pU6KgyybWNxqk2a/0lx7qToVq2hZfrknlYckxLaeXWtUeNkqkdJLK6iqKMrUSxgHCgJFKu1
l32uXWHa142kho7ZKhWf58brHReCqY2b6m5t+qc5p5sNNp1BHt8WXgoFxLanEw+Z9kahJqcDIReg
VVMfoI8SahZM3Oo2Cro20eLjtufX+ikARBR8DXemuGPC7Zqg2W7IBEC+GDbHJJtUDxw7BnwS434g
fkNycJIH8gMalypEjpeysgiLqlDDs6OC0+zC2J8QWP4KIL9tgGUNaN3vxnM/WeaOvgQzB6m6/Na7
CycGuFIVImOOMQQkJJTF+SwPw/phlwtaD2FD7AYvmTrZLcQ8My/2/dKyqVTSZCV32pJnG7HEPMZn
RxoCWZO6CZmhvT1LjG/3RPZJC8XfLpusxbwgVHursiXCwr+c3MvqelvpIOJlIm7cg8d35ukM0zV9
VmPzlBxfHYntJ9cwZNCFb7GFLfNK+bM7HK3GQZY5wSKNvM0Akl0xq6N6sOwBFcW5mY6fPBhfS72L
oT+bjE0lSqYKsCbMk+w1pMTPL9DC87AQCqla1PnZH5F3/3ldER9fjTJUfOfq421GOc/2iyK5hw4Q
BNj7paDfOTs+X/ImZJypnQIkk2h6idaVC8y4ArX8R0CX+/SI6Xtm8/oB1bvikvRH9JzRVqIa7gHP
Spm0MLZ+HMpwQFXOAAvpWKSRt0NI9wiOUVx5EHJaqsqRQfLbgZQpTNkBIrwcEy82/tdOiT17d0AE
iMds1Rwmxz4TKZKAPEWyESQV21QuFMXlvE4wehgs8Alf3ZWkYq0V2cW2iRqoUxjcMib4sJD62UGW
BP5y8mASRVTE+Wv0boKwnA0Ve3/ukadTi8EChCDKZmR8f1lHdMDrb2H7gdoqY8Ojb31/85OPLdQ2
yY2rDx21dT6xF+qSioYpSrpUrWvVfeGP+GqKsvh2Nc89JSJC71NLL6qRi8GJXYYNbL0kIskzxIYO
XzHCxnWsxlBG7+gci/8DNvaHaMv1R+Tr6tdpDe0Pr9IOMSwweqCJyPP3KCPYJT9OofN2n+knsBMM
jq/Q4fapvzfpyh0fnQzs7DlKDnT4CdyPcGtj0houjOSi7l0xxM2gHLoNMQ1Rkdiy4wlrCLREge1S
Um9LRbsVh/LFw3Ch/HAy0xUx8iK7yF71L4eYUH6ZOAAke6xTSYSxu9j7dUiwUqT0Fhg45vfwq7UT
eRPYoXD9M/I4bErAIdFJGp8fQFGBLnsVA99pStwOohonHHaUAayP2Vx7qHx0O1IIGkH+yrHlnOOA
1MPsKHbNdJI8UlptAUxRRw4OwGgdSIcRzDyGzTYFOX71UOCPVJwC0OVbIykldoXGTZIL8JXngHVM
qZSrLGHt8sBO9CJKK7efFyENvU0G2FZmwIS/hzDxdL6OD6TDk4Q8AhwWGAQedLninS7Nu4qlZJlF
Ysi4QBs/5i+PO0CclQ1Ve4aaNal9oCBycj+cZAoXrOBLQkoVbFbj4HiEMZjQrSEf9GlG7X1n5hwZ
AgS0DhvLXHEyTt8fZmmb5F0EfMpPx49x38rq/8T5qM8WfGVj9vAWU8wfAAjWS6xe26w3MO9ZDYR/
AoPSdPqZlOsTmAvMYUdqfedSQ+RYsoJOeidJDAmh2AOF8yEBfoH06EfYIHEFp06pRf3rckh7im+v
XMd06bZF4f58rV2/YbOXQO0K0RxMiKrHoVE48+DmU4KSJWwpBeI3FbP/Yks0cZSwUFXZd+iOpYt3
nGWHAMA8EI8WWIMxa/YUKbseEIYAVQ8kd0uI/yue4tGr3SEzdZ9IcZb5afE2Kbeiu9k0UYIUScO/
WqWUMcStxaCSxgthomc70Tk8SyG8cfKcJs/A3Z2s2y53h39IAgGfEqvIZ95st2x3KSXEO1sswH2P
aMVm5x7NIlazGz4V7fxkKMWqOPOI1aXDx3fQs1FlixBrrco5t8DL3CP3ROdH5gnU6ywJ2hMfFGdt
wlZTAKTs+JsENCmB6ffvGGg4n21GfkVJIiOsP037VjZ8IAvg+EbiXHX9fDBui+No+CPXgs8OjO8i
yayrktPvP0EgQCQiSwb4UwXAVG4Ku+6FLawv83woC00MVr4k5mwQe/4KNQAuHJWL2vZPEczzVUZ1
/+wLIgeRuAJf4NVTxqr5HKP1jMLmUw4Ou9C3yDacVOfnK7FGYb1aGRSNgvgNwXbYf22wd3BgB6at
8vRX5/Lu5Z/hPrkidnvEavpM8dxl61Nh8msyR8xvTJJDinhsF9GC14XMSNqFnNyu15WHm1dO5I1P
zd/6P6czI4jDy1eZTreEsy5CzEK0OeLiGEVDMbfNlXQRPl+ZnkOBh7JWq9nN0idFxU80kHwVZ1NV
UWu00x5QQMjbE3NpdNxAqRhvrnzAU4xOnqHYg1/h2XgNDBabN4Wsg2zmLUdJdqAzgqXssislAu03
OdZ/yBkW3cxugbd4mmBc6BnB31LVk9CblQdCp4CLPGyVsxPIbxPbDvhhojHZ8755ItWEbPy673dS
0FSux8Lnq+FKgd/elzkaB0O0bWhXKOSWNisHpDkRx5C3S9mIKP4v6lcD0JId3icj91aUF4NiwlDx
gkkGQBfjIgMHIL2nLw8QOvZn3R4C+wMrLFi7uw2OMKX1UhBR2ckNjp42JmTcf+fBrc4mCcQwenBf
Ln5xYkMqJYkrE4M6ZXuj4wk7+NwrIvmQx8Ht8KESJPwMr8Em8VvXeQNaEE5TNaVoeMmrqxQwrqH9
C0n8mA4D51w8O1LZvVOBKEsQ2r6FJMDmGj/Q7nt2kamsVZYLIJaS4wMaJEn2guwAng5umOVgxFeD
O3f3IUey7ob5j7JKGMDcn/qwhHpV5UXP0p+V2K18qYPqP4L7CorBn8Sr89e3ULEmokka+LyeG/mE
X12u9TPMU38nbhwGrwnIicTgjZKLIM13rA04ko9MPdWWolT1KFyjTb5/AQ4MwnnajszOJ0vKvUAZ
HkAhBXkV9Pvfqrjydms2J9rk5WjckQ96QH2pFxv9x5ssJg9Z+II/d+B/746X7TXspJ1R+sIakQfs
faOBh0vDuBhXKyaKt/Hrq9twotwRBKdV2eVXJQfRrSKUniy5qmh3WWo7/SN9OCdPh8weDmj7Qgke
XI2UZRz5we1R3R2XqRKLpslBIhsj3OPqwLU60QUntMF7QKxTp05jIXJYTzNiosO0fp4fAgvUWV3+
iSNsjJDKjRZA7KwcIh2LXSBxbd1CNqSHkXTxtDibqsAskhoYhVqkIpV+xJ1jtupF84vmhn6MjjvP
v4Z4NFBroco/UEMG9663vAaSlsLEpgDNROEZhS98tIeCT5baMtxjyqPmag/yN33F9xKD9lXpk8CT
S8naGKkBw3zZCV0E7dXsmR0IxiUEM42scLOX4+QqNGp3jlnEgYcBam0blQcdf7LyUm+tTF3sO5gb
kzIk5gNYUO42XZE6YqCtr3TzR/DXuyRXdPUFptbPnWY2nRvwxMJ16L4qIWL5uZNJgYs6CItHhKb2
02PtEQ+mWLoYfnyvnDaWAYoeq9oOTmZ8Rkuec5phAlAZHzMJmz2UEsBwcE4AiD2zAbslkxtjYrxM
2lVFm70I5pvfo6z+Ibw/9GZeNPi/+lKQHfZrWo4ZgXed5v+8Fv/zt+tajflxcQYmJMnBCsoxY+uK
LmnHMOGBnC2Vc+GEFlXuhn1IOVX3vsRxHvQHBh7LoxBw+ysDVyYcdLeigANHXa1OTsrmiH15x9aL
QRrKcXGTRWYFyIeZSjPtef6ABmW8IC9k8+jBXJfcwx/5+gEdK9lrzB/kS+gmyk5FyKJ3GFwX/unZ
xFy322jHdkc6UD0lQgMgH78uSI4lqbfUo905x4aUdpa1cwy542nSYeGhGjLLYFA5xipbflKO38YQ
QpCuYmwwzEqTQuz6/uyE2vJD4yEenzb0R67wlQz3/59V37FBo7p/RegPS0GU+79gq0IxBxupiub8
cpatH3U4xYw8jN2yF8QKr13Cm6WNn8jgOfnml7DY730bTksrWrJmkfPzxtKt13mNc34RTcODGXsA
UzT64zWDJ/32U0ctShSjFcFaW+LXLsHmy4ghTPI/KfyIuqx4Nlx/HKB4WxKGnHFLykROMY55HEfd
tBcmiI9QcjseClBbgLV0fqiukJlogjAazLd6ppeA5bcimlQt5h36nRgNu25WE3nieQf0OXz/qCBd
hjWriXxRhjoAe/3v1/Dfs6cSVOJqVehEgaxIqyqURYCHxcqlagEOJenSF+m1w7P7TmSYkNNatryv
ntuHIYcadFIIBSeKsxT94mLQfdV0ILHjDAgBTGdFjV7pcLv0yMQlxRGbm2OeP0oeXnCqPVC/btWK
3LH6nQvoM1Pe7H5kZ/JcosUMU07II3XtmoHt6jHGPtD8MSHUCAWwR7BPcOKkNdiTMIoEfHK1Htyk
j6gnshzWqg4a7hXni8YbjEXtpGMiheOPw1iiOZfyH9QUNrQJiicq6gWhWGalREizPQDySKtyhAxS
8oUf8c4TNuAHb2wzcl4y1wk8cSVoxaicH42NN59brH6luJQwpawRPr5DzxvFLzgMAkmFeCxy3H5y
k8kGWoQOOQP0ANUFGDMR/8uGP53cYSu1zK3lWGRSn745YR2EhX4etebvkz+Ui7+H68n5Z7iXxwe4
FGU0gZyF8R9bpGvetK1Gf02hSZidGaOCj16Aiz3Rt1teGePUyYvvZNatFMnCzHIajgE/k5vAtgL8
RIlFIxxF6ynLjVwKyM/o3cZw9sSuOlM1l2KRIy5XQWdoHaCVR3kTeuXW8o1jummoC1iaXz6l8MPW
ku6Tl4nzn4jil3F5LM91yXyKvgtCQzkhZrmrgMpd53gf6OSiS/Wu/veisUANmQpeSKiM6hngkSpe
Jo2RYlnSFpSG9fxahbRP49YjrWABBzjs6QEZGzwAx5RUoyzaHFy64cS9NnbtIF93FaCiliCvAAPa
AzgvanrSVJizkFK4JkGnZSpbw6IZkeXxYwzuIQg5LGuBd57gP7JCjWYwzomFfxzB5HCxQeDZrrju
BwRFfhtoM9JmkVF7XaYsCoOrZAObsvXkqmPsHeweMNnb7EenBSUGJ7/lTbzHjXAaC9WHQ72YySpA
EptqiewofKJYx7jMN5wnVkIMuY7QVOrJB23h2OOewqk1zaZYI8Bd32h7AD6XlfntWagbedklmr5w
HF92LHzgJusHuaP7aNHD+jGrHTIsyWq2HuwEgcbNv46d/ZGG2HR9eojkDo+0T6uFDv1e1Xgcja05
N4QxAGKUDTAc50usYbjc9pU3go7DWVmjEGbu0eO7lGJa0u6OmK//3ncBx0WROLOyBxORS+3N+IXr
0DfpNA84CDv6Vptkmh5rTVugCGAVDsHoDDvGVfhL+4TQDqoipiIi43+m8lIaUWciqHej3RrA8msK
JfEmRY/pfjBpfRkygoxDhBIjpRhB6luR6hxxkiDn8dMOlZ6c0aCXqMffD3z/lQN7hLF1CkpDaD2I
OjA/kf794LJfeCRIpmGcuPqcQCWNAonitxNIMd3Hba+BVzJRft64eRqnnmktRzADMGZubmONTDg5
eRVy0t4xeTRmvv6GKoKk3CaLRz5LFM6ai9Wa7+lO4yzBkas2D9Sw3UJpyS4hqWaLNDVPvbzuGORq
ev2cGZ5vRi4vC3mCqESDXGNiMTa+EjaM6Z03THe5fhGlo+e4VcWZpcisSP0CbyOEhYlKhyMYDsLZ
9FDCCVYIHrCDz6xHn71/pSdp/IYnffgUlzX9RAh7UDjXdZ6JmlHHzUNE2CaO592kc7G3SpoksAQ2
XtoMYpyTBOGvRo5eWLLM1eSM+3WJC6atN1FudYOZA4nWu1qpKHOnPum3eTFWRlMygxZe+Muwg9po
GdGkZe1jbOYvHro1256pqJ+kXQy3vIET24jTIFwrUWYJPEfmA0VEA447+YAqcwph5bOw130nuAz5
b55TLcZ8gaGR0KBBrBFeA957FEI8CuQj5uD9pgR2v77RJW+bg74IY/zwaYOAFjffU3VuGzDg1MqH
xc86UmPQnjbj+looh+RWRpFBdKH1kjlcA/NVZUp4APEqPpOBuDo1GDZqnAtdzHyjhCP/Ize+X+Ia
FDZPje3+vQmaQvg8QDeZW6Veimux7t7BSSaQrDj60Tu4xlr/qCbUl/HOd7R8GVqJVgrXlixLJ41R
NaODJvxCY+dhz9750QgZ/PiamAN7uoQhCFwNS8Mb1vBaoqnfPUmxfAfQpAcuEKN7oBX9VamyUMF/
CZWF/3hagc3Ql9pLlBHdaLkzbE5go1CXYfJG1DCP79o+gj08WQhg9LTcnNYTWAurg3rVXVY5gZxW
6TIy31VCFP3Wb2VeagMBFAYwgRdRjAwh2cbr4xcmh6/MGuPnRxTQqR2fTZfRacTCks7pgphHZ/bG
21kNXywyLo2fkE3ENIbzx8eZQLIXVZOQCQ9GjIZ1cCHD253YoS1iC5JggQ6Pg92TrAXwLW/LLo52
Y1UAnQFpimI/2e64bGO78t1/A94bgvcR9v94GCIfq/1EhDqZ0FnA8Ektgxjs5MuihOO50GkGv669
mQyDiu3jLEofojjUOyFgYwxcNEG/4KDECBl0X/HQmN4vEMTFm7+ZPbBO8xel3I8Z5ijXVWiDOvGa
cOtaQeefwPQgnl/MpRP5P5vFxE4nbl9x+cC/FIrVJL4SqaxtLepxbJvfUUKNeuW8Sv5BsW9rbpKF
CGrmYMMOH5ZYxCVM9wULlJ9g5hCL0EL6yXZBe8x7QO45au7hqJAjqJxNDoyolzzSBzVrpf31b6bV
qy0/Bjk1In4cPELTYRzWsKAUHMJC8I6kLBM70mu2ax6t/UKQb4k6Oy4kSkvnfwQcpesF0YnOVzYU
uS49XNSDDqfAi1m6FZgNCejDdTPDHfYSaDQVO6h0X7vdczq/8zFwkGaJ8YLzus8L9JqSG28rciJ+
zUcDn3PoJuiep7OuSLLlDkvLkykbPg5IaPA6yB5UM3SWXw2lhzRSHGe/dPgSyEYjXqiaUzDT83Te
7OsVdMtfEPlPTcifNt6UwSyA7F9QcEpVNkyBjpgoTbi0Xul7rykMH8/GXIWpY07/eVAMNRLVaY0Z
dlcw4JHdMvzOdamWSydZy3c9hwizTGZpoHhVIGTwtFiKIFrBrNapocWs0FtyGhjZLO7a24vMISIf
mhJvQbWZNBFKS7uqckFc2bAm4Ar3E/nzw/23WHRTYT2RiEdC11oGSzNKEn5qEdQgEB1qIWU9/aBE
vUJ4YB5hg2t6mO6mJkKB7nVOkOR/hgP06zPG+AaUN5L79LKg22PGWJKxU3VHnqqCSoZUIAlWRkMR
Ac9Xi6RRlfCZhBDhRg0TVolw7KX6nGIaWSVS1WY+3jd3td3VoHfDqeY8m+exDDfReOJnDWGbBzVd
7iAJLgeUcNN0c3G6GR5YtTz84Nwy/Wv989J5kEFpqdD/f2gUSYJfZjEwD/8oR7AVV6qEpiVoTeWW
AnUHJzwExUfhNTpkqMZBLXauHW525imam2ImFa0vsoULq5VSq7MV5wH4sH3OYZk0jmmCKegLH2LJ
kS+LadDhGI0myetxsmlx8ZC0OcNKzLYb4yiKfC11lMwEEIbXlEytanoKssIaiMPv1kbXjO9lanDo
YJuUjZ7HEZ4LFl/RE3yX33LAe1l2Hyqa7RkOHzPpnTqEfY+rpjl1bOsAnzxVO8szLWfoNZZt6vUG
UPSnRTPckby0NHSzYmyMyRxmAg3ZCj6igFI5iS3lRgs3ujEUNHuq+amqEl2r9ef0ZXVlaVvCbI2x
oXipy8guJmvaSwpOlqnCSqC1G1NfOyLbtDvTwe8FT1/DYxGLntNmitSn0jMcodKVkdIrTPY9RLSY
CsNyV8dtZkX+SExEvAo4iQuvSBG5JolxyfOYLcCcMSxMoxwGTpYmiuqtMJwbMCMCuC1KN9RNJWxS
R6Fupw1Aj/hz+gdCyTujevPYDYw005XlFp2K8kQgbHBueu2AyqF9CiROI1uTAfRH5B32X2x55PgP
I0m26h90S4k+insJxy/co923xTIhJ1Tb2VKdxBCj9bNzOVlhYpgwSlb8BFR/0AgXH2J/J6Cx0eDg
+KnoNUb/InFnqwHIZ8ozPSyhJeN8aENFASZtdLTaK0q8GXHp/N9fqUOFAgnTjZLXR6GneL36VFBC
J227ybZWJQ1L8Eqaa8pv7n9tXeAKObxmJZOBdlhg2Smn+44W50DOoGcGyLbAR9RsPXAEvxFgOo91
GufsVAecDDN3xs9TFmEp6NMvfQX6TZhoPWdpXNVhKa0ITlfPju2or2SDUnq/ZgZCvem9qTNxDAov
3JrnP4ldP0Z+3iD7tV3MGy87Cv4OFBdJD6wox7ulVVwsuR7cXOda92hsnd5JCLpS01SqBDHnOCVX
+OYF9ydkmNPsBG/tp9d7KG1nEYpX8bxPP/7FOJUuGTEqiCLwEEfdRCoXL6zM+kPkHcReCaQTnd5I
Cnoz+XJ44sfqhq6cgF5Wbj+/A91IIZ0vuocGYOyVv7oVWPLsCGSh6J3hq2RxDAwFLF1tYT6eI19x
+5pLxSvsq2Y3yUO0BhloOTTGuN19unm0+Sybwkb1OR+KvIUFuIZ3BZzpfK3G1gyfNCeiJZV6LNY7
2bujliMbWlI9h6ejsavZ6/Q5bk2paFWHW/V2b5W+rkNFdRyyAo6SLP8ZYVUI6Q5nPKSmfzdQOD0k
L6jV3e35lF2v58BEb3BBP33lH/CPe28nhTlSYBLi0zrk6vX4uRDirBFpFMTCwq5l/WQasZpckiO9
zYX3wJKTnHN8pfKJeKG5xq+fvONJjdTRKOuTu8uFc9qi0MtQFqLNVmjsCP/QqG2FxVtJO1nztJNd
ig5XZg/WMlFiYSLYN7IxCzxnvqG1y693yTfF9tXG4lK/y1Xxml8Ftl9u2KIOy6jriupmk7pC6gFc
w/PEj4VhgdCr7zBDUmMuyLPB2PI0j4qe9zTk1dIn55WNMXY79LKYw7VUeXNvSQMFeUcVh0gVfsEB
xelaajd3+ANKh9HtXBORqOYwKI+vVUeoFFwkav7qfwIeZMusuna7nGRMvorE/wZ+5Bphkj/3arwi
l3sYWQT7mYRjsihWjoRMJqhffnH0SLNrbC2a8ra4w8dvODKIw7efn8MM+94nv7j3mQxizLizY5Lt
KSuTyfPoeeyLXI5vYjJUc0P7OTt7yMJwwBUIXfGoyZ2//DhlINDldnSByvvUeXZq8vZs9d4qT4af
z40SpsHOOIc8r4tsP9cbicHTYNFiqi+RWpbRRhyRO6aJaxm9Ecs2r+hp8roeSj89jPRM5StDPHgX
BKHTQDyxJqLKtOIYJsCgU8bVlgJkKXa3pwWddCKgmrki8J0Rv1Y4nMicn8xGgSFWWNv0xDP9wQJ7
uxbzl/RFWzHIzg5OvkfSMehTmTgf2L/up25G4x8S5dI3JHl+YtMUzbfrkeA+Jx0cI2eFcTQp01hD
veaQTR35MA1Af+oBRvLV28wtde/ax6abRnOsgFCDm4+T/6EIBUP0ktNf6VBDlcLo+5m70st5xyAM
64DG/k4W+lO7sr1/mOyhBO0IdH99rIYeHymJxMeTaM3wY61IZg2A2FnNHCO3CUGj3zJCK2YV7rMa
Ek0tVr0DLPML0vEzHrhQXwqAjz2EsGlA6syT0qCZx6L5PXnYRgW4SiXj3o+0xya+NXDeRWCVFgKd
VwM+o2CBD7ycsfWyRmU0CmqD5mkbhvOb07KLEKB2OnVEx0I/TLzdRlK+Pm8IgiJoqybNsrfGOIch
/RbVUCz3LCb8c3R+d2YCXLs9QhvS1yVa2pAwXQqaZSJUGHc76tYsFFaXw6tNSw8TMR4rCaDY5BFL
+dm47k1ZnhAX/9nXJUodXtQt+w5hoTcGuPn9HONF5CmGB6kswiMt53lChqNSkHlgdcyrL4Qnfnvb
mPkD9kLiovdzkPW3PRm9soTMyinmQRBwgQdPvfpcP3fYIeMe+BzKULf0h9oD8ce784uF0ulYCA6O
tc/Y/WlwnXPRnuJ6mFsdREiUYYH3LBA8VsXNMoJJuIFgfehUsrjZLrOs+DJsWzrdHdgsG5WRDWWO
C6qAPV4Ot3D02saqLHplc87fzThMv1+rZnkrVFQHOxHF+C79li2yTawLMgK8I3WIeBvNkpfn2wMl
9eb/NwWNyddq5mivv1+A+j+RGFR7D99ohrIM8Rdb6767RUR4FyF6QFpELc1EnBX4qvT4cuQX9ktH
hLphUZ/nBhntXeSHnUnREVRnlhRvjFJTrpeLDsLW3uMRUSDRTz/McgmMMgkbU3IeP5k/9zAEiSaI
Uq1jzeU92/ZF+s1ZHM+YQNB2aCXgVlmOA1JUSNvrQCfdncxfw+4/cUbxIE5ozC0j6E+7p/2Qr/C+
DCPRTSVLrryUWEEyCqLQf92aJVgcgbnDm55XAbwG/TIU0i18eIQ4ZXHQf8UeVVOzGH1wotJ5SCuz
06jmEi8btDR3p4kzxZ06Pa5drR/Z2ApXfoZpUvP2mO3GUfqr8MUayw8aBxsSJeSDf+v6J4Yqk/AC
XDPjnNhQYoIcFoYIObip9IRX2wYpC02SRv57IplaWPzLn7oROavu62vwPudRPb1LHlUlxEyUimjI
8laQL1Qez1RcBVRYDBPsTUedfvDqZw0O6YE+FLEf4tCzfx6wanvQtPS1aNpcyKf0awFwW42LktLN
7z7ErbIohzXEcAwN99H92gJ8wSaFri7jZ3ek8r2EdJdFhE7KGzvMyI4oq6LWce7vI2QhDviQY4eW
LQa3iEE6Dty2hp0hf1hUgIeJ2ydLwT3powLL3l0lqYUNaBJGoTyvtGQRfclptkm1otzPEbDdQdd3
Nq+LMfrpKxm41MYTl8qMy7/hTcLScKRIjDi0NAx7ffZOqXhaNrfhOeI6+G4fUJ5N3MRJyfxh8mAE
7OHKA7G24T4i+ywWk+t+uBy+lFr4tdiXsMQSYYDKmtx9vjhaFTrraXkLGN/frl2GlF8r9YVa5GqO
ostTDKWaj/wY2HgChE/+q4Ct3I1ypcWdkfZxx3bpmg65KRu7xKNSu2Mxrs7EQg/K0hZrS0WxA0sx
hVjS5Yo0B6B4g704PkpPDkcfb93m/uCZQKeZZH4QSuOyI7lHlb0582rbZC5m+7T3eh8bS8BgcSWB
0+9nrKK02K2zxY1IUIUJ/YH7IGRJqU2q7Us/EJw9sy6KDr31TPu1ywvkI143Htudm+4Ky4na5JZD
3jOw0thH9XMwuO+hKzSq2j3DmMAOZM/Wmfg3/v3c5P/LukyGN7L1YjH5HydPlvTBBJWCyCMc8vL/
YmFZFkcqKXjYlnkP4U644q02Resu7KElMn8bG0hdi7uYMu3wDeuIZ7YgudBIJK73lqP8lfaEWyH2
JhTYjzxUSUnxWAM6cmV9ZwMmSZcOzCGIzoWVxm6j8L5ISC8O7c01EY+83h1m8Zb9dbeq3khOSiIY
28RPKo169r1N7GUy6yy/r8A6H/9ex2yU0bqHK/S7aZYardE2dnsM8Q4QYq2zUUWICN9c0n+UN4xU
ukaN1GfyVz2CRbHa6q0uiAh7DH+fFLbuN6UlSgB7v/GorapNan5nQQibd92OzXK2Q0X9UYKWpABz
s83k6nECPWYS+ljLVzrEABV10Jb1oaNoH0xCh778KqC3l83E4+1fqzFGDpvydpEy1NDlnk4jDDgr
cXs5aLbMhw/NuGiUDKJrVFJoDT8m7x57Usp+P0/9aXRqpdW4k8KbPMWbNIm5jajBdeVW2BHyrcyf
SGIO6oUlNDgxVX7FzEpQNa0cn+GxvahWSRZBBxyZ3foQgSxs+Y4fB3E6cSoSpXff0oK8e4pe5wZZ
cg7dV1FrpPg3FndGCYh2WS08Cmwfu6YhYyxhllvoWh8q+mlWv8Qy+5OYPjTAOKpLlnZTjAzj9fNt
JfUj91YGWSBRQ8Tvm4tdyGa0QEuDjfTklosv8r5DHF6ci+9ycopHbBOZkYzmf0rf7ZytsDC8Wi16
hONfxNMfjFQ8P6FaYRz1jfkiShvrr/ScFKTP19vhXtmVfu6qjZIatMQVUXM2PYjki6xO/VNDXtzo
sj0qnM9srPUBFLUkc2jTJG7E1IRkhe/qhFQ5dxPUObQGuJwAZgNsQprlgLdfFM0O6e+hzkdK8kPj
30TIN8DS84zvcMVjggPivqCaf/jzwujm1G13x40tRiAS8wEtVfFvL0enOzqjrU4z9m3rPMqGF3S4
VC4tWoB6+sOFllFpvTVMBy4utJEsG+VSZn92G3S9vFHKLxAlKAr8qJQs4HiDiQ5MYxWnvyaY9Qwc
gVpEmDQdlnlBciKQnXXpfsJyCQrw5Vc0VRd05q1J5SD8IFszWxNPrpSQK+8FY+ZcjXVZ4B38lShr
5wic+n6KBZLWcAC27D7m6hacnAOXKTB0XD0YTqTaxpYc9jubVVHDeFvMHl12gGpGTu8qAZcR5jit
U406k8RjNRB4umNSg2Ax3fkSOMaKXABeX6oY9obi+u28Y+FPba1KiOYEWGOm6foLPZ3mcWol1ysj
Ykyk28QGlCEtC6hahGiiNoA04mIDsJbe1OmFgp90rEXyIZpNmWZSWOju7mUBKI7bw5Or3w5I7Lny
Dl5yfy6tx9mMVIFYLfjukONzOOzBOH3s//uyESjYi8DSxsyfVwG/RO7/VCXTbm5fNPN5uCtC4L/k
mCPyxu3+DzU550W/APfOlC6BxMugd0m5XMzhXD1hO84SEx6ZdZdcqkwCGrfHkk8CBto9yulj+oqY
8DDxAM+ou0rNkdATR5r41Hoj6RoRBOVAZnrrSr/MSJg1/uAvBYWuifmhc+dd8M8Y45XkgiEW5/LC
woOmPcLv/YUeQE1NnUkWOaVeYVf9gNFj4EXWwz+9BzzAN6iq86HjDlQF7siIqHgt+phx4TpED1bs
ivaMedk+ZWLl+J7iQmiFbPR/R0Vw+9PseYMfCjMvB9XBSuVaxxDb6EzEK3yLa+f1Pf/0k9bXGJNP
MkPpb+bBGidrwE40SUej6k6ibbSBVdy/ZDgaKiEB4dSXkcLa+vNjwTgrxGLcLQkzGJk+N/+jmerj
fVYKsPol0GSRYw9FjSsPHpB7p+GHkFEGLuEQ8gN7CXQbIYbHAXv1UK4cl6V4pDdHXb85+SN8I43V
XIUtcP+dSgTExhK7FUVsCzorV18WQwC04oMav/qwRJWmFFaKLRsyBCWmctEmhyNPICFcs6RSRJoe
onKgMR8Jkn8QJl3Ctp8cvisUt22p7KW1Q+RLJRKBidYJ/R8pRVaHWk8ZQPERAEzB/Kuxpl8Desn6
ioE+hfIJhlltciAD+cIShlMW+EwQqYsd+ozd8ncI1zIFm7MP9cK6gdebOpsMHFkreC3Hr3cjJU0M
PnpGXI7KOkh+VaBTPi24kshIbcLOdb9u76VfNQQ497Ng7cHGQICqX3SzzQ+00XRvra2Jd1KRxJco
i7KTfLWLXeOpyKioZF0ivO4vDkxoQTfByITxRna5E7fb/5/E5CqgxWNQQ8wxJqXLwQUsY95+7WE2
qUTx/3IKQPpn7kI3oBtCB3Y0VDtqdNnfjv82ndKgh+PbrjjQfDRYVFwmxCSaJ4sGuztI9BVuWtKl
YKdVRlTJ3e2bXWIhGgSXkga1EqiinK025RY/s/dMu7mOj/RlXRc/hHvyMG/gs/ThMyCnNYdZBJUa
IrHyTc1unpCSyh9dTSbUQrfLMwrXZJhh1Stjc49+bWZURlpl1+GomBPFypUEvigb0DAHO7bxYGfs
fqmoHgZnHenRWvfvoO9uecMAFfspxHfiYPFE/rNQel184ZcxE3Hrcy6+cgR0Yd0jxfT/9VVVDjrV
b4kh/gSiuBdDnJ7WsfbJPa3fOcORZxiS/gCbPLNnIbtc2lpAIxr0SVqAf84xbXRLIWdMrUQkpWKO
wjVHnNvEOKAliNm6Opwiw7KnFadeZHa7fOC8yB02jgXVW1rvErlY9S1IGepJPQqaytEQsw1qIKJR
ppFEbDYbWnGhFrbHlmgjZOfQdLuSPJ0uhiKqv3SZQW2jgsc8P7HzIKXISmuEI79KVAlLyYNU/bIp
ACWuGoo2EYk51mDe2SVGvJ9D/OwlQiOtRkotbRttIQnrbin6/Rnwk6BQ6pxZ7GvSLRRz+iLGrwzM
m/D1s8f2WcBR5SlgBmFWTUxI4IFaU/CEfUyGg4B+O7xobIhwfdXQCwkvrngNFrSkojSIaKMtsLBi
IW4ey8P9OZTinFTIOcymTCJliCD5aChBWS6UJnKmkLmd8aa77t8OPwMRs4BlgiCsSVCl0tpa4DT6
a7Ws3gVT3sDkO+DV73Zg5GlQ3CtCD29a5AlpPHIqbEev9rlpLDAM0L1TxbfNWeFL6goAI291b6Eg
HzhfG1hptUqGjJqysDtLvgAeVpPbEDnUoDLhotFJPQ4VEajB6kyf3JWCpXoVPhAzEM9lmLah7d0j
oMxfLeldaFYpJDdMWouK2Y3D7XIzWwyVOCWqNiNFLE6sG6W5HCe/XQ+69CFVMd2yiL5CEkTps4yc
xy7d9r1dsPCFKTDFNSqDXtvaEJtVXFcRskdvlTNyObIcGMWP6+7M5eyXB81YW5WmvCRnjc8wO5lr
Fxc+tgYkzQrucryI0j7Wgdq9iU9jqc3+2A25P97OC6vttkTwLQoEy8P6o458usnMg2fXqY6APv9B
4ID6TUN1dTirqyXAOVrStkcz2+YYkcTlCsQS535RGf3K3atM2iSWjIHgQWFNqNJDBj/pmt0kh0BF
/1ANTvL58t3jGjg9YimkQQGPkdl9kMIE2/D5fBLXGcC9tbVpFMQoN/2X3MiX/r7hfOch+PNGrZnw
s+bERuRNi4tsL36aIt5jOkhLnwr4TKkMCzxaiB1ehE15N514akQ7sdvjhrfcb/PqmTU1//+OlYwc
HFSrhOJXqG6Juj7eCHKRo+mkynIRmqmi/pwoa639QNCyhs5W6UUtaCN+iIvKk8xn33qcC4m/hy9N
6hO/PTDeLFTR4S+l9iayuZdwUjI3wf13ppHjREc0U+nFkeqerQFh5qaN3V55nwDXY2hYHLF/DEfn
uqdADRvCI9DoaN0lK/6GrJJW3lUJ+qW5ssgmBtdMTkMjvKFfKACjMMyxYehntfvPF+U/E/Nb5v9D
8JeONRNfV2/Dw6jfEftTcBQKMku6X2mHp+xiDvK0/BQjQhisN0DXU/+Y4smfUaGVXpgzSjDBVJ1N
JgrzQHsAaEQNJCfWMVVeav6wPZfD9XoDwM9V+lE1be3uNVIWEFhlZH+WP0n7DQGBhv0xSCWZLTQx
rAOQhyD0quOaObsTqu+xPwj2xEiqOjYb0pKjBnZzA/xH0v3IxqPDSwa95A6Fg6d+LDbyjZ9qw2Ug
wld3v5eWH4EIQsdgep2VW0IDbmJptL8qx9WzRUHBbnOvcnY9W0R1lwzVYgwfJPNZgrgepOQJ6Sl5
5ULo/wydakrz6GaDULsCtj4ekzTaBBU7+zuoiPY+H666pFT+BoVBjh/aSwzEwurPcCDALAIS0FTD
P/sw1lTxTLbc9NkCs+O95rGRFUKbN/ii0UwSn7JF6oOG5iwxCWedBF0MxE8UC3YtJqZ+YmNsFx2x
UZ+7Lj8xhgTE7QlgB4JuZ4IxMAauHDxR36SRaLHQHTOx8pJL7TtdTa6US/DWc5ejCA/3S3q4H5ID
rSPO/A+ult3o05JXXmnyH/3ZgLsBC3rWanEAZYYUSKvjAZKr5ekMfV7JX3DsGBjoRLqw8f/ffjQE
P/U+EWHB+mqZiiHVwRVq51p6800MZLXF1xrsLVXMjGxUlAOSTCAbf314Pzcqw1T4OY9udcmUOwBE
XQHMSqvippGsGyzASIxdkTKSGrSzHaa13v3oVSpCQdQcMKa/EnBUQRE9QYwcddxQnsXnk2e342t5
1x5pxKDjhuTMMAVFPSP9u1A19kxG74ozssdpKV9grCTjUY7RUuqbdEWpcF6uXi/xKMXabpBoBmQF
teMDUuVJqB2Odiapuh4ym3UiQwGljkbGOXEEPMWCNhgoQFXHt7qkwEzFHzKwNzR+EOEaNsba72HW
kRhsCd1YwzVcEfDYPL/26fKPLcNygaQ4nrYU/QBNsya0jlEr+NG8MQsP1LIPwmaSHncDMtmYJDDl
BcBy2NBl9WocbUTOZYxT+QneRkIe+4OQ9AC29bpGkyC5Xd2iOjN7B6+Eymi+i9OtPXcORM67xnnX
OexOJ45OWGxTD6Xvj/aJgHF4+M50A+6/HFxAt0910t8P2vudJfdIMIhe6WnxgTPj4VzKNgzbQYnD
j1gXeuQNSG3Vc4YPNTQMt+oBRavdRCJiz/UPjfNmA+988BD3nI0KN0APUPVtTv5+fqzxW+dm+y+Z
KUmC2uhLFnAujYOA3lCePUoJ0Jg94PX4ZEn17SDFy8W5H3z0AJDOP+0mMSxL6AZMykxxg9VDbfo8
AW785fT/MojgnVAlhBDU63LM+/XvLYROqbSldB/LD1SpXY+lIhbG3I4wzV/XjiPCp1V3qGfywSNW
hUP+yi/f9Eu//QwGJjo1pdCZEoJqCC6ryDlkLwt5TdV/Y0E7d/eVoRYRbHN3UQ8DI9VJTP24ZkYd
vvL+CL7rP8GxeVg2+VA4gT0RMSoK39Xuq7Jju1Rae61OYIXd8J8URcAI94G53RBFl5341i616pNf
7OQsC1sJ5uRct3dhnp6Nfdy/SbmjYIeb3vifB0eIaqBRPQ1H9PgW6SRd0eF9RIpChz56yQrbGdke
dajPgXd7xKNop90xQq2QvpF4cvqHAbuxdBq7SL14B0Q+CJ8501Hpdpe1nzwVDHYe3dkGrg+n5rVY
EII61oof4ZLbeW6ufE6yUymLK3xyGqd+ycFFwt5pHbXF8spanr0sSh141LfPQ4ro9iEjH4k0ZpEY
CTGL/PjwoR6Eqm/u9fOqLGJXmHAV/wRRTG8uT7Xrz2SQeTfppN2ZkercK/PqozPW3u5bVKSEsFo+
vQXX83f/HXLsX6o93tazCuoKS3m5qa75IN3mwGAaQEU61THEzuwyDPneYj38FXdEgN1ua2CloDOm
xIRZUaq5No5kqwEOkQz0QwjDuJEKZzeyboKVwS+AOF2ZqP7W0Co8pMEJ3Y5iEO6+YqJf+qrZfFcw
PymrX8IU13E5MQEJUj2AYDgSks6++I4tHqsNbeVpVR6U2vkwnAqgoGIO2QdXFZC/uXPi3Gh/oC6w
7fc1yxn29dsZ9Fu5oHnEzRVThpicbI8l9+kyiBwQpPl16k1SCSVZQSDaYwoeryatsnFLTeoKvDW+
Ino+N1b/yZFkU82QLZezPsjSI0DpTAIUWGUMPVDjgQbJ4NR1FeulAiQWi6lHGg+bUh8WpMNr86ea
DLQIBROHu9pYlal87yhua+OAIYN3aYVwr0oCAfdQgkTmsss4zMudUJzM7E0RzvVliSVtaaCn67Dq
gecv57xZk0krhFlNPNbXTyOZp5VVKcyOQhd9KlCzVCxHmot7e3h08SuMngaewJVtGk9RFDBbRhF6
fuxD4xIVahd7r98r4jEnDWOsjHRxDPpmZisBfYihc6RmBoXTnQ/BAoxGXc/7T81mrglPJ3wV/zrt
s2BqLU5JPSipPtaLOdUB9fgeMOecPqDlPQIpIo91ep+VZmdC2Ahl+zWa53ZYM1y78pgI3XX9MFNm
L35bJkZC9C/ZeP2Yku2Dnq/7Lyx084lK50CZGGa1n2kX4dCYX1rJvb4i3YAjvmdWooSe0jeLDhft
ttwmIqAg7gc8vvx7FypgopAXNi0sr1DuFkl9anr7pfd3bn/n9VHUitRsUtH/IlzsoWj6btp8D/QH
EFJTA6gBRuHeqIWHGgm2lfeNkJzMKkpwoaTERgTIxF7kK8Uej54CSDb29PsJkeBg+52SfMJ1PAKx
A2F2Lc1tROTmYqvUXjufobd31oqN1soYIgR0ws60wUALuHMhnImmxBgwWcgyUrFqpFPmgP7YUs7U
E8GydyraGpWnrp6vBwndThPVW9F1NEsb4Dt6zI2By5m6N/TFV2t+Eph2U+/56DbUlBiSH/QVqtrS
eYNTpLelV8y3M3qJ8MHeXaXjIVUy7dtzPg37Z68rv4SisXprTjxqYW89y/Eh62THghNUHomlcjfc
Dh1PhkY07WKwadepvGtXXoKrtFq1b6QVp3GGIOhfjxlrwIBkySdcQzx03SNWSSJS3hfdwgUebFXI
vqI9zRzELn76/N+Zjf0RDK514OTvVXJNrTDdBIfqPtGtmQXTSJ7DAo9vZ3UvsVLLPAy4BkajCymA
pPcY8OST2pMopBM9VQ4lfYg7qPhvtn/XftZirV+ew3Q0xDGc1eoaCrIIxkYeo2VHnoq/zd/uRgLg
0F1B+z+FHh6/RpckVW/hm25B5PJTXrBt8jrQ2ORAZG9y4Sy1hskjAsZdyAR6+K1KSdFBhM7tID6G
MnfS0ddb28OMQmmHa1zDzwYV1ITYSnP18SC7rU5yQX+0PwJB7JjC1Q1G4mgZTeHFgu54kKcAGVAj
OCXJUJi4v80ZiW+CNtOa+Vl/U/knNlY+GMC9jwShBPWiSEqOOR9Cqu4weUtI1pPR5cv2EnLoSNLl
LRp4csUHwArPZZAM0lCnZuwj4ENIXb2lCVcArK8n2U4B4orUT66UWyYkl5QvNZrQy5oQ8dwMKstp
IXP62Q1OqN9oTj6BovksLkVl/a4EjG+0YzjwJ6WIoYG6KQ9snfhxkLRYjoEKovbt5FV2RYV6nZrE
YM7uwlqxuq8KSoD3EH29X053tAUZjntynU8Qo0RYmdwjIKoAy0NC6Trq4VTBR+IUAYaFX5FzoTnS
Eg1KzWI0wxDnSyokw2Z5rYelPcLVeFAFzebhk1cwWELAcg2ONd0BhLbkx179ZmrwNaqN4wRANWQ2
vepGlslW2VvGbRKiM4/0PhALr1IjVfMHUfqAHjtBnxl0MYISl1II67aq4GmM9lNnekhfmmdBtTwI
k3q+0x3J6qh9FRDqg4zSo9ofuMQwBbDSUwHo0tIEziQmEv2a8gC8Z5bBDC1jDPMkXwHVCRyY0c2d
3/cmQTBfmzWe8MAset2qZcJTUIzPqsQxY5P9x6kPMJ6fTAKoGh15HUm1My9QWBlvKyPb6dCWwA6v
AYKC7XVZY3WxBjtSKNP4JUiDcj08FyVspzfLGtGykFSv8TEG8LGD9dc8S2LFEc4vTJSZsN1kczpq
8YglIlC506c4ESlLKnoq1FHwISLtd681XolcyPnV1RgYrvVzVPFqtdIRqZ3Bd0YQwNZA+m9v/C/A
u9lDUpYyz1EIlx9X654z+mrVrnqwX7CjwCAGN98eiai8W96qprBw/W4+l3LU4WE+KNywj8an6Tve
P/JMGucMubvI0fMzVChKZq12kLTBlZv0E9YFTMkMT0Vlp4NmcCpw1evZIqspJrveKIAnIiPmoPE8
GqG8yIU28a/SKwQWmp7EevkEGCzdm85rQoiumrMF8nuxvEtpa50NmbYkaVHIj66Q1ievlMfVKukq
289ZiWXjzRDLJIdofjXEy2+omjN5pztOz0m/YY0wVa3b9Uqi+7kVlqeHuvHcH1oW6spcAfHW8Nsh
sWxXEpWTeycQE1AqrabLOpgpx18OEmpey9MBpueN5QcPBn631b3tVa5Q/ALi2YFR/l/LwSN8xLdP
s5rUQpx5mEF40q26wck4aVwmKAegOB3d29SX6h310ONLl9bNockF3+VvUPHDV9XXJm72wCSNlN2n
YsZRHpTkS5g37HtXpcvJ8KQvHIfjLGLLD6P752AnmC0lfBmdo8LMwIJy+QHNWXkJD12muXiwimXN
CMwXN9Iq8kAuhZjfBXNloKHbNaYtIu92AVsry/NAwyUNVNn2xOhSV0Otts5tiQpnRKJySxrU4Y2f
FNe6xFX52dmSamyLwLrLMkG7v9E3nME5SkxVES9UDkpyyBiXpnoEoqgk3zbWzhhDK/+gnBnXzibK
wBOnE9WPn0QqKK0wkjhNYiWV506pMrz/PZc8CvI6AP9YRoNUfXR4R2ObnmQe77cLa/CY+7604sSx
LAJVtUsQjJ6/KBM0lGc6pr1RH1hlPJZFWiZx58R66Fk8VqSxshvIo7NjRBk1/uRYWmGTTuByRSBw
b7zpSkTRGWp3cr2NnJmmTNqqnvw08fMoNG1eqlTLI63wm/M0n1161T+vzzEy6iaV/0WDIQRlvaEe
AHA3LMSgBiqDUbue7CCE5CxCb872UIwHFl1Q9dFNcV9QMAzdt2qJfKeLdt9hZSn37MkWdsJgedn8
KGGCs35ysAN3yU3213QVdELzio2Y54WIJs2kJbV3nmZ0SB1Np9J8xeXaEFPIHY6CukSGsIkAH502
KOrtNULjsvf3vnttgi7g7Q5N6GxJi1iE5ZhTrAjlebNMVTz6CbuG2K3XwmQqx8xBWaqvavGiHtJM
K9qu/CnNAuTgf7CditSxqIgHB5y9r1mEoDvSR1couGexZAUbIZ1os8EssNii5zz0UCjCNRepug/x
2jTz8ROkpfEOVdfOFXw8DxVUt/VmoLlXEJ+NV6RR22zoIEwbJ0D1fHclcSWwyKGwlq0f9w+ntcV1
KjIHRkygcWrxdfWdoAi83MNC63UqGE/2R3hF3a6d4CTAdZeYKQ2Hue1+okApbhyxhWr3K+rRC9kR
dqv1ZBRj80nrWoMcGr9fJfeJ3f2w6ceTFg3ky5TPUUzw1oMzEDrdR87wu8juW2ZsCjE4079Xlndx
afi55THht2FmH0mHX/KoDRoChuFIDt1s/V/x6IhkwGnP2Ieyh0e3ANwj5npkG9OE5ZGeIgmXjTlu
Rw71mnWSxRu4fp2/hVXgPuBaG07E/XkN5eATrfpBjz75t9CUxojlT8DVn8iUN0afz6IFpoE/BnBO
FMU7Wn7KC29lb5lwex4IJpov064Epovk6eA+sLD7MC7alftQeeIeofQ/tM09zehgSHsF2elXi80Q
nVikGGD4Q7KimY6MJOFohRXb+QAmypF6bQPF60iM8xZ0WgmTiGbbH3Tr3vcn8Eo0WOWvtA7FIUuP
4MXurR7qxtpNnTMuggeKXeAA7th7n15ieHiQHZ3DLr4kJcgIidbLEKdadQhYRar5oQ+i9QY9L+xJ
Q4k+GgnYbKez71eQ9pfFHHsQgAzEKeQqTclpkS2N12KER2/QhNXqQ0X3VO79Vu5e8IeXSD5DWxMs
BZbARJcLeTC2RKEJQiDIJwODnMXrZm4j2oJHp/Z6LsZ3l1p1T5nn+vsiCnl8r9MuQAgCNRGEBaCL
oRtApvbWsmXvLihTn4SZxAv5ziX8tWmtXztf0ok/iQg7v+jd52h2zaS9H0paIyI4jiAivh9dJmFq
2uGlHztK45I1zQgfTYbR/H1wafocnDyiVD+BYNbDw22VRhp2QkkSFSYFpC0dLk/HTe0Gz4lA7T0S
meXGAgpLdb/ouMO4btHzNMEVVWQJYOhNtxdUFyHu6YmX/t89lho7/XLmROVbocwSg6X9kXKJCIF+
wGSDKUIucZfs4ux3DsdezNMWeK8W0sMskE01a5qOJiL5VXExW4PmuysdZw14Mtf8f15i/JrNkTdn
W0iukKWV0nRBVVUQabgpqKK+jlBR2TiK/VWE0/t8Qzx/h1YlSLuCBDdYvvMZvpptl5lUJWwbg/d0
0vOFNq3gSYVUSZBqv8h3TPTbIgJBCPHIibJVyGacKoZZJojkz+P1RjQ0YllVt3vxfSPYRsOm9CoD
SYNy3U5Mw6sKdQOR6569zm6Gnel87flN8F/CqXVzraD55S/75UOrrpPs8CByHRgnMAjKlWGOBsIG
WRDdUzyAMhbmEOguyLMrIDTHxoHHvGXu5PWg/q5ry5T+woiHV4FSQhQMNQPnuvGFJ1aUhgOFFdbG
UaBVAlqe1EjjfGeGNPswxL8q/4rTrlmWUbbhCu95dS503QKIgZAFY3x4FPoC7yrQtix0O3eY1W79
nM3fMaGzjAYJi0psBviU7DNRH9CQeFGF7oFnhgTYPaW1KnUX0LzNYVuKjEJ6NNN/EEBCSyMert2d
mh3geNO+h7pMRSryjWFiJ0JaCClsaUUYRitLUa18GDHJrPLW07ZS8HM8RY60nRxs6X7NUl5zpSpt
6ppkrd2M3/XNNlvi0n8/CMxzoeP0F6et7ms7GtTUk6vxwNT8vyz6+gZqUVjGzLVY70Pqby3+eDsW
HcR79EWvOq7GdVcn9pn3GpmcsAjEP9uwijG339ddT0N1TTI2wwavyvcOGeQB72zYm2iD4esXzOI6
XYQI3mKunJVD0QDIIr21PDFQUfL+WBzluTyBU9Pfu9GJME9B5aWq+cFzhpjGvrSoy9I9nBWZBhjw
vkAgGul+RJ2M9zH/XBWPElfVUfpCIQNRbLTJj4DpnytxU38hXb5+E72dOTZOOQRWGe841lMINj/g
khDeLZtV+cU/VfG4c2Gn164Wf0lPqQitsIXiFQ4KI6b8Vai35U5rqC705JFZJgvGmgYpvlV+fOVt
Sfo+tJ+ojxwkX+0dNKbPzi/z6CXYD3ZzUxU+3r2wlgCv33+39x27r9/NsHt3IXGk+pOQH7iN2yrS
AOXK9IOQAePQfbRvjnPmzRS+TbDPEaQImLAQ0lBaewYmr+22hQJ6tHzyA6voCvmb9fIyHYqlPpUl
8TBFq3wR191p0BT4WDj5c/VHKwo6R4m3jAROXnt1gdwu6ry3qx0FNt8yiU601rpzDixeJr50fuBT
3zXzR7VhnleApTgpGzQyxrjHLCYrkLXHV73WclfIF6lsA4ZIm0Np4nCEAplADw+YGhULopaPwME3
GXBenY4tyO9GDugzOzb3w7+oNWBtkaXiSbFRDKGuQo/FWeTBYT6lGZAQzK1aTPo2JzcZ5oPsUOLt
DwKmoTriMQ6u5Sf2VVXcbvO7eQ9g9uvsTnMYrWCDgrzwMRK6XL5Rex+jk8HSL19Vo6OwpBcWIFBg
NWO/BqtBYFIWgILRuIvjUIR92KxTV4D/CrljnHrfx0WwFKMlHHkMboF44j1YngK4B76ctGGZzOjs
sadFQP/RM2XfA1jZm4Ycft4jX/S+iOwr2ayMGBzVMfdmVCvJwvCfRf4nCPYBiw8zNn97/gSYXmQ/
Ngpkvt2JKg4RPAgJARWrPsz1Y2ncTTymo8r1kJMbU1/e7zkiCSQa0u6heuNksQ5MT9eKWHRrjjJN
58A5SpPrLYpQb3lgGDzmi5cnZBLUhdZZc1IPvYEdTigGmIpDPSGdlloT3qcwVzAR8AK2DK8Yaljp
2zRR+afbdLEwknjlfNn7s9iFpMG6tHPaOGvelMNtBZ8cvCZNCeaVP12avIt/FR3SNRtooo0Yp8tD
/fO/IHjCQrQnDTLA+K1ex0MYUmUJc0YdUl/VQc12kriJ7zbKKPfH/KVKerkUMxFOLuXJHDWWQ9TB
key9M3cpiMtLqs44b16ivP97tzVTrGQic/oyNy96fEZCQ0zz9lXSro3e59a2HJCVtZ4OpzQUJZfh
gF7AIgg8+WiKkX+FXt3pL48+oNkAA2clIAJ2x2YXdhccoJ/9K+J9vt5sSfZE0kZbjpX5vn7jx0LX
tEZtBnroMUcgQCARPhcQOSnaUA0xlOAYMxRQC2HTyvVQV6Sh2E2EEx0qSrGd29dz+Wc4K798N2Fj
to8IKsupvpiXrzEXdpIZj5p5qH8dnPDUBV6Zs91jz1qgjt3ip5l5Y1xZxjp/f9794ikQo/jveGaO
qn4kF2HpsZ41QCG12pzAKHYqsEEFMKqWBdatC4NAWqlkxSL4YcZ5tllC5fMgLNivEmt3yJeObcrR
L5z9YfWf/TTtbUwDESUA2GsQZbp0rwOhzSg+t9khp79z9U7ey8ftLubkiuA/X7DLEMfqXXF9tsyy
niH88lcj30fYz9CigcwrkXXkqZGd4jJ8hEjz7Q523lgAXp+qv8HrnHP0EhInSii+INxMpbb6IuUl
A3QelHdVIry5n6C/koqPKRlwiS+b1b+u4+7CFQFm68CO8XmXWFBO2kkPtYpnlCVYFyZjWuzLF8CU
geI0q8LJhnVeHdcwITtr7gnhWRHm9LGlzybrtm+KRi1Jn1bmKub3zFm0o/3E4f5NO8Upex1PaggO
XULF+PvhIXxDOVhgFlCpwSVFpIX84H02eX6TknVtLYXnZTectBVzyWQvO5ARa6w38a+r46KmetRX
VQKGIEVikRj5y6nqXqcwfMDJQiPNFtvz67AGM/uunxYvyWqsWE7sRbYvn6cQwlLJX8ewvQvgFbM4
ZPP804ejZp5SEX9R88PoM/SzhYSojhxj8L3KHe+n9//8r4tnI9NQgkUNyttxAsoB+CdBcwvGyaFd
UcmAFSVy29AQ2v1YAcg+NgUCqeQN/vtRhu4LXnuLvCX0QUCBAjqcR52ghU8K0VEe241Dkif733tQ
T/YftbExh6MRbdf2qdZG/lh0LfRb1BsTGSU3x/G0072Myn/1vj7c17bVM9c0f181yMv6Yb8DAjvu
0mvAED9KCRbQuXow6k2EcD5nvRn8VP2xDFj8nW0yF/bJy+bZe1oWkoo7VPWtLKlXRQ8MGvA81Mub
u+C8A3C1bl+bd+r8LBwaG7lqeMiD3al3qI90ddgkhieay8Z3HcQdfQuNM5aeSufZZOsKX7kn6br1
VK48L86ZSd/IO9xzFKfeVMiqSE/n0QwMtV6IOnKagKHrfcnwxuqnC1KxE7DF3uj5CveqfGwKZuVa
/q+8k5V6lIQzfawBPm2eW3f7qG+TwGnbRp2Noz6PtUED1MJD5FVQM2a9kGDq4W4hycvwEX2POPZM
NWxvFxsDjMykcN+jBqb/nST4cJ2wGOWoxavciV8zkd6L7TphnD0YMiUXsoRC8Byid1fW+jpcPV3B
9bLG2ogAFJz4CGjvGX/YD09lrFDNSn2hMxMyBWSpph6qaib3W55oLEP+f/UoV8NR9uWIIvFQUzNv
uO4Cxu5OVMB+6Pvs6bxKl58JcSSgorSo4QP5S4b9Qwi3/ikJGnJHWKfZZ7o/60u+0Tln64/O+prD
9munEyxwioJnNklVuuAdEEE/UqfGi1yK6dlTT0+HpwCwsQivDcqcBse6/4d77pIvAEUfy8vaDEs+
qLouqaPRDyEM3Sf6qs7cv7DitNKur1WfGiSk2kBcGXXnHWNVoVjdhSP3QIKB43Y/LSIFgyHyLm4h
IbX6QDaDvXVB+o04ZajtQ3BufabnIHYJQpB0kBBbOkqK9eCaY/5j0DLY1B/AFSGL6scFAS4CNH74
cmCNKb1F9Hg4TicOKf4oKo2MHNfHll+zzCnsbktEKpx/fnx8nfCW1+cBbnhuhjVmMOuMN521I0Tk
U9fs53CSUzj8uJrRqUHiKSREvc5QqzhJOMYaDUf1unp4yJHb6sts9PNwDeLLOuGG2HJm7xzsGyh5
c8zq1fPE14y/FDzQ0zqWuxgeD1B4FN0teoCPzXoSYZgOw9c9ndpV2NX/jWEkNgS+ewd79QdIoWVY
QSG6qylHSY8JGYDGO3pZPDkbIkNMvMtrbhaKaWvC4yycva8rf5irOQe9HzcvWSg0DN/aCfxUPgeP
YXV8Ho+cNNm0ZBI8r4BARldsa2Npli9cFw4qEV2CkaWB8Xy+pMnZE9vWyOokfqYtB8+t9Mn2wmpV
fs8Q75trkx298h9DQz7KMwtxat3B2KSDkjI93vtFl76G6zam4V2oFm0D+mApiTl62AZ0TQy+fnNM
qR77dwt17d4xj5v+/KLMB924d5j66MZugxLQsDXzihwJTYhwSB0n4xEb702UmNiYkIi2jxf7c1ol
Hj+4wayZtI6uz4/edLOcnbI97n+dXXvW0zeEzedvRZg8edCg0xyHjBKf3s9fdkK9wB6NCF5ZB4sp
6dOD9FzOrMLQqhG1A/NXIAp/BHGxnqG7jTiVlqUgJQN1WXjhBK/pFse5G008bq8CqoDObPfn4Uyz
jq8zR+j0YZ3YlCen0+KTSj3qQOE+BHCREVwS63GGSDqHA9cb/2L70htbhKRdGWRjGF2ZGCVImnbM
QncvQ74SKBnEiz0xHLCzHqqSQIzGv1Y5A3k3KqP8ZPAczOxKHXUd5zsEGKRWH8KDzig9vNgbI1Wb
4QIu1KPfgTrv69AhqW/CqMyZfPWUCZZgA4PA+RlfZNZUAyfrvaw9JLoo1AWdcEK4t3nwMyHOXHLQ
D4ANdx6pouuU8OvNtAgioUq6gzp3XhpebPR5a5gMB3QihFIBIXrcPwHNv9gIawxZNt4dGomAPjp1
VCurY3pDpR4aD0ojTWIBEcXwEkJDrPpqjfNFz3VtK6HaJtZzqaVXvuO5w3cyn3nZtgrGIYHGTniO
TH97J0N2Sty7tT3wJ6mlSzCQfjXStCptuP6yrYpeCKJEf7kRPDdZKmrjdTY/Nn+3S8J1qLKAAVdW
ZsKxyQDp7wt0BOa0p+1WPZ4Nc5kOa3XI9LWsqzC4up5CABu6CS142sr7mQUBYt75F760vYvJ0Sc9
8l6DkPcNy7IwW9WwUoA9jVUtSFByCqADhh3Fz5mnx5lyuvzjB4JNWS4GKlHt+D4RO5t9zKNA8WPu
br1J8bXGm9tO6AEyEdXy+n0/ddusDkGIcs7PSXoCZks+01+XWzsmXI9Y/ZVdD9en8nSU79or4OWF
l0JyOIDZxAwFtzxt0sewyn9nqgpPqTCbaIMMQqj3XjKjN+LE1QzIWBv+aSxoElHJEgV4BzHXdUNR
KHUtpinwq6VVDX9UXMfWkVvfEGkVepsG6+ds0D/sIodlm7zbSsJUnE2DqwxqYi/lyW3pSV0EW3i/
pTJcQaSLkuApvYZi7MuUhvMkwf98C9/Bmk+cui3+uqBbFAqnY2QJ7wIjQ4yVgR5MqMDX00UA9yvs
/JiBWs4o5rqtS4bf9e134ST0ice7cI47X4RHWJLDG453KHJpJ8OqlbLlzYR+C67qAC1PH3F2xdcf
Z3rWgrY8UzDhIOOahyaT97eWB0GVBa8FrsZkClgSHrALqFpEKy582vU30302sVLFLcnpboGSkibM
xo09DgkDU890CxjgQdRcSaU4sgwtwdKrccsPQDKBFrbz9zvM+hyh9eb9EmHmkj9/fUaVjy5FdQr/
DCARYDOo18kCQC+zeVW/9PMY96Pirvu6cQib2n7VoP/i8NOHAdLXFZh8k6CvpXhQs15N0mMzsSLw
9afnjzvin9w6lcSa5IoxduLkvArfSro7omm1U3Fq4ymtJ22QVWgh+cyvaYTgqV/P/pEWvX2TLy+0
jeFd4OtHxxD3Z18Iu979TBOEi2pVjXtvu3upC9sUsdN/wCtoxHCeSXwZI5XLI1nlxbDef1K5XgU9
Es9OFkHS42c0DeJ2yCg8vh12y+G06lTm3NtzHJ1rX9gCyTEbs1GTqi24CKZYredB4KqCodNsWTDE
HxslTGwaQ8zWOId5F3EOtVxR6awTNdL99mPMriKgZskI6qCV+ZBqgycmDHDL63lfq2c+dIOxF2uS
elcg8QtfFFQpHlsJ8xnBMcAuopEeS7SypCHSsWiX1P8+G2tXoaY5u09bFKDnpudZSkxvuk3/bERF
dmmSVmx56OmnobTpNV6sI6vZ8HJm7TLm/W3vvwPFtImfjtcEA2l21Xtu2aynnM3lnTRvY/gbnY2d
qzwWMcNZXElPZ4XNKA1OWMK0NHQN1pbXCc4Fwq5ZwHRMfWxdr5wTkEEokB7qP8fC0E4azUYN0yIs
30/nBi4v/R3usDjP6NTWupPlzjbg3jyIpgBFB55GvTMz8VKoBGo7fZeJvKrvYPckS7lpb1+ITXu+
mHtVhUyqxOMlzhkz0q9VP5lbtw5XQqdeULa67dWdJBw5otAs7WSoCQJOTGVoa2n8V19HDA3RwAod
DwYd0pNTXmebOBC5rzHtu3oq+VgdSZBT4zG/W2mx/Xh4NmYl1Qn0zmBtdgSLuwiYdkcvZDlCb5Vv
zmIUSFlv44C/YBbcHsaU3GBb3A28yxUEjbm5baQmTkr2SbarPMGVqqn/vtM82UbED27ksAQ+xnsP
X7dBh4Z6WO+ORGfoKpUXhJ4ykHOXy5O0CxXguE+IKX0ttYS88NCN7sTLZP/YT2pdAmq6sP6bPdRK
ZxUWnLYJHAwZbnK1r2Ktl/IqcbvQdsmGRE+wq+Yln7YpVgwHfH3DJOxJOAfZHhwbH5DUpxyNiaHt
WqxVmqVfLrwfE2iBiGx0/JdYyw2xhh8CqFusmKb2TthqNUCItT7y1RTLmWuvbYgVPsxh4OJqan0w
cVbbsx1BH0DlOFDzQvA0ENyJsPCDcx3UTiBJX4EMSH2PyTA3gurJDE4RfOxQVaXyGv1vV4m66VXo
g5gLB1avuNZgOh4IHvt+yQTmIuOtCbMPgOcc7n9+isQDschk6u8PWhk4W2xm3xRLnkYVzZJjp4Cc
wsUWDcSH8Gz0cba8b2TtsjRxBRKSEGPzqlt5cWjT5u8hRwFmPtRlbu9Qr8fhcrNnL6KtXII6ceNy
jCxctY8EMfls83ZeoLTEXg2NIjdNKtYfG6hsV02D3mgfEC5rUjjWM4/ae/4JGHchC7L/0WZ5jlPh
zVTatQgFbkdHIcOG5Rqm+GaJSpQfPWfOr7e6ocNrgW6Ox6PUcfc9Fv0y2QfkzB6K0/zpgfcngzkF
S+DMlXuVAi2kWgqg9dg/29EKSh/B24KouO6H1yrTeAnqrAXjzMa7Val27QQGjqLADK3pfSkxQvqt
48PVyjPdOVtFSIzLvZI3/X5gBE5ubbzfLmrOYrXExBFgluCFyuKNfS/ggC/m60EDk6kzHeTfbrui
pXaHWImOt2QS1JOxfykPWoEdPfXeN82hPIsHHwsWCDyilqD81TJFEoy0R4dHNS/amucn91f7mbGD
bbttu59nue7aey56vv6dn9AeFsBecEh7+kRRIK3Djxhc7YKOrN4psodaqq7z1SFNAoLY/1hXp2vh
cGjwTcR3VUDVguJ+1lnAo0BMK8HKaNJTCR92xUfdZkuD2qKlwXCUjULh25j2Xi+2aM+SxKJCJ+5Q
HglXJ+mlc+K6DfR7R8B8QBluIoP9UFm84KMQBWEUrT3yZKpCGcgIkdvaZCPn1hdx/kMYpz0fqPsu
slMdh0LFJD56cai8obW3tB5pIlA3U0ZSBwI1a7l47YYuZvIxnlIhz9sMJLsIf/71atM27jzU3nTh
MSh6220K82BB8ueTgONCFm+qjdtJi5zJOerRUDIDvLNY+rs2miHb04/9uBpeA5vP7qy4x4T7gQjt
xauZJs8vt0IC0WsVvquV8pzQgkDizAWGZFdHJzCeYUAXMU2IPqx2+SBKouiK5DDTrZvz6n5jre+l
M4d0IDeWo4VW6psQcl3rkNDRAhtzq6JsGJuNNAwJGCX1ppAR9OMHZx/KK2yHuksT5UpO1aUVWuoS
Ebx2aA5UovdsHWojpwLmAhwOtnPpIn3xLw3pmpvCibqskFwOMgvm7pXBiD+Ckeplaf8Jc7j78arr
p2yXGWY+R/gdMaRhmiJoUdu7AvDR8qlTqUDetiM2HY8LAyd2hiLseCsZYJRG0SAV7NH53dqkvzV4
UA1XdY7IXyfQvTMb64CIURnbaQ4b8YKW5LVb2USeoLcE0c9B56E//ngjvq8O1QzMpDlngi8HZSVz
VsNRSR0YLkSbHwLRLERFTLwfdEeq3Q8n0mkW/TNcMljMLRhfvMhh/jOKnNEB4Fp9yStCKDuOGjEI
TwEVFDZLOB5DAoqFS7ESGKvSoYRE/p+U7ldoh7jmkXklRlpfHTnfXr2eB8wuPlokATr3siYDUGt6
YxhOFvhlfYr56EWDodgKLULvEBrim4jokbIWhLlhvdNmOZLqDGr0NgqjeAIjtO75FJrnMnzinAwP
YHmtuP/wSc1pzg1T+MgQZOECZulATa7tlSADtphXOvfjQmEz7hQE/p2w7KKPiTc+jv3mxEKOdQ0U
S8OhTEsEl20vA2Qkw6i19QaBklOFmDRPJILxn9Xzi91ZJMVhV4HN/KOii+tx0cHzNhUpa+zaHbQq
P9yGMfPyUr/7PZ3LzWOqGqCquTbNnbUwjYwl7uMCP/d8P0cpIHEZvwtg/1BFZqSfNrK3sBuC8drd
o8GTk2IZoecPOT5eUazLW2hZ3GtRB/vZ2zlr+a1Oru+q44e+1UsQPqcI4wlif5eIvAzRKWJg1u5Z
dt58Y6RMzubHU2k0J66VdHfDpQdRCFw8KqriRNiZ0fH7BXCaVrEh+LUOyseXpfJ/JxtkDaNNUGjs
jHpFgi4dXCIG5X3e6Ry+dNsaAAUiZ30aDH7D9edbenNIzBdPV/745VftejbrqFOuFSvRsTmPZ3ae
eQ9Wp9EAiyJPG3M9zhafAV8+v3FAiT/lKtZ+mjiZGnGb7HPOiC5zGsMYummz1bdTRwBWZubSOOZm
3OrWGwIiq50VZlmXcFeh0iGDizzDM+jSDTJqJUlTDq8XJythQDsz5yvpge7SJLDgfxVYKCnlT8AL
BAABDzbOUHmEZgykV2BcrWKeEkxaxAhrOczF2IEi7V8ik03Z37XctcOwrVQWMFDznCy9ENO0Ota5
CadZIrAwQQA1T/Kivd6bSPIEOWaUar0gsvAVRtv6yD7FzbDLpPYuBd74qQLpmaleUwgjeJn8wTwv
zDEkQB1jG4pytjAzHXin/tyaS8Pry4G72OkwLfCXaWJRrf9DKUJuw2bOn1x/ZFaeyQbef8+iMjry
uvYF9wgR5Mvmm1L+ub+/pmmphJ4GZZKuGuWg9ouQa/QIhPVsAc92aVAcVhwpu50tWVbr1FQgoeQD
w00GXBOpdQUByJjV+EjQlkOEIsc/dXBbu9PwdWJd9g3PyOSbLcO7BvWWN5UiEs0CWDxMgQYJh8pC
UTwUqXBMyoDQL6bv218zKTQIsA5eM1wvwZ8YO6QtRjMP+Wh4mDhxXOl30DXh6tLCTz4LlhwB1l6d
ZzU2mOjmS9hX+ofXciFj2MeVC71nXdV0aSFa7wE08sUrEwKBTnOaAULLqoAeoMey6MsVfkBMBpnq
Va0z/riDumZYNQVtVrjiJVOXuymYGcCGY05zHeGQJy9tyGynU8UB1PFJL/eJIIkDAhTBDFSAcK8t
XRl6akw+/YHKRkmSaCgejf+0PLdrhXddrXcGZIwGp//eTalAPQhD5BhsIFAVJc/N55U++CNq3z6C
VhB4MDiNjxxOB+j6yKCzH027NFT4+q2US77vZVgN9l69p/YE4bNoXrOPLEPUicodU79kZz0cK6Y4
jHy3H7LPiIz5c2+ZdRfpa/Hrs4dER1zwoPd3j4J89EwkgEdyaLOOpba5RwVMJBJ+QxaGnDlUAlVK
CKiMxkQmHSHxmPaw8zaaRVzgO9kzyUhPMpil9PvwjuheGkR3oHRYyd7kzKtLvFJphxN/qLJBg1yx
B0PkxhHkVmQ+R9a2DeP1QPTfyN2PGVftOghDPQ3ss5MF1vnehtc/y6iICY4829dFdfwFtJl0aNGt
FwGT8mjcsevxJ/GdcA6Iy90rvsC229hlTuchuoepvpPiaFNrifoQJlre4zbmKFlE0YhBRXNByIKq
vYPoCDMTuNcaXri3QTxdW9b4a2ZzU0vkqamFyHzCZi8/CmG/hDW08obExhSJt4TFM1kaqTq8TP6z
QqfBK0Hg/27W4GoJmmKWoQKi+LsVcJNHfd5y5ZhJUY7kWwHwvsAlIuNxVLXTDUO6y6cHI2HB+Ejk
/xVH7kD4yLHFO5tp+Zdf+R6zAdb3kHtKOm5ghJ1jzW447/+LQrGRnEu4pIeYtKav9FmKqcevmOe5
5ZtNJsQuyipD9Fuq3MbiEiwvRnMnu5YbJnolVHgJ7nAQzLF9U48EitpvitEY9BaP2X8NFryzoaCH
x77KmuxFlcxIbGQzzx+M94EETLozoipkLLGZ7g4DFIcfUT6+z5i8A+Em7S5PV6QH4q1N36QsADrU
c/AXTbLPGaLfePJR4Jt/2vW0BX3k46EjXtLxSthd8hl5GWpykFcdvOGiDNHfGQpvB1rVDUBH6xNn
HkJFY+KK6Tqn9gJNecC0gJ9t0kLCGVF4WXDQNZ46NISFnXvmax1oW1X1jZIz6MLEI9JzR3TVNueH
gAtTz3KOpQy6fyO+mppIL9cKK15HyNFzCggysW4IC7Nv76wJwUKjeQekxdYIKEUFRLdw6BqBJPvC
9e0hxi862EcFXhOh23yD1gSy9N/UymYWnXW8ym4be+mb6HQVGXmisw/rfLCnP39qo6h9Gnvd+tot
UDI57T+4rkcygp8S8kNUP2uooFP4g76clCUAnq9dncFo1bJyFCEcRMIVqXhTAL+evZ9wtKro2yBw
s4Zy7hDCciZBLtiUg21QnCDrCMrNa6X4J2+sTSFT0P9U8JZGm7s/Yyo7AN1bVE8sFQf+3lZZQ9x7
e10u+86bZaNIjMm7Og4A9b6svedFCyq/yCaG0nf4M3xlHr8YHXbZFoCIIv6u++3KLt1kKNESYYCM
n5RC7rNebBN2j+EnxN+gKnNHB6IKx+4PvHq+aJqVjPsZGte+TGITExqrv+jD55N0xLp3PbnM3hD+
Ag/iG4Bd/2RbVpCsp7YaPNeRM9/EabwLikyxComqvyY44gIFjtFiGvN621qzoQIQsNZ7grcX4rdq
FT3Uh6IuyHzASd1472eChNzkt/FF3kBC+/aPicbIIYM2PYG+P22SyNchDYrzvOoQi6OsaGFuocHb
Fl0k4Ksf8jl/xGMy94BU47/0Z0hEYmcCJA1u24dE3vTNoURdUPisEeg3nxyOPcclwvmjwZ16qQT6
gOIbRRf67zphoHwmIwiO56N6vnr1oPMDI4Y4TrOckeSqOTabmCQ90IsaA75W0Rj8aOE1FUmOhY7e
lLfn/z/RhDx4HS6qIGV7+KrntdUucUd+VJjh+EsSb+oGqiRJNoFvH9RC95Bg+el3S9Hm31n2PN9S
3cs2aVrUNi009LitzDMeEZJGGHpU2xTMVamf2oXrIQnxOtO7HmX51VzlfpDUTA/46Nuudws58JId
PhPWvrxrwAvMHi6hcbHvJHRjHne/Pkhl7tV1lSqq4k4rmsve0ifOKCa3/mU4gtUz1OGmRP/qvzvd
liniC5A6cCA3e8zRRQAHhMmXufpTH5BWw015AtM6CN9yN9yexd5vBck5TsQVpbwrJCZFWAjh4m33
zU5ZRa4aZy5kzLk5Br2ri26VUAkxO43r7j4wnhPGlTZr0fmPXH2pMlLhgWSnSpz8G4t42GfPfrBR
kJM+EirR+tkwEwi5uQ6iO8g8tnN+UHQVeSAW8vzaByQ76YvaWk63C+rqVxWk/GGT9XzAIPFzBC5O
8Eqrcf9u3H0k7oS65cXFdrzlnpj//lu+XftGRFJrC3WSGawKdhl7WwnypY2xHi7J3CKpuJmIeN+Z
Nq4cSjEv07T+WUIYSzz1UMGnI8fy1HsvCOjuwRbXe1QtLijO5dhVVaf5l+Qeil+QlOXZYOalOMqe
6/hKdOLVlEqLds1LBRioI/+aI2sHF4ccQaLzeQror6LTfgQRqRbzoz8i5CNEucmEnRd6lF6lLt+y
lLg9JA7k2JikMSaH+35pPe17wLUWZq3k6pHN8LRdveoG5ukfalSmGoh+HSbYOF9XkMmQuGdf/+ZP
t4TSIkhGFkD6k/NAvnMoDA9nAqMtJBVJKuGH67BUpPm10z2Y26LdWjNBUMprYmMZ3LJBwHN+nnUp
zvpiyzt/9p2jXz6JVVkT9S3r0hRhMWcguC477kf2nodkY+6WZkVjqfYMkKG7/W6qWhlwbLjzBlnN
kxkINkINhAc54HyuIv47xI9II/5EbMBhACSTLsk/+vItF6MHyvd4md7cQvncpr3D6+dZl87QtwE8
vQScLLpvuyz8IO7robelEfmSonuURZWqbZc0FDl2Feyjs/HCdOjGiRn5T4lvkx8cxpcSbMrVVhYn
VhOOGdEkzFFibPyfta3o4mTZZehgrqoiZU0Lm99elP68fVo6QY9CNBLKSP42EWGEHj7PRHkg7jqc
PpH2zUENLyVWFGso1RKTr0ohdHdERjndiR5eJnO6lsX0ZkiGFqVX16LMTWq8qc6yK/2YbHmvBVzN
Bj+QUTSxT3qc9k96p+DA3o2JvuiLhHVwx0bTbwJ8A4FhAET7na33vrEp28apfzs+qg4WRcRRnOHh
3SYsFWuF/yqIGxzvO9AfW5Qsqb+NUZr8i7KKcTeh0AnOz/39jVs7sy+VYpsM28Db6c7VD3BNQPUn
DJP0WiP9rTa4io+A4SMzAuE5L3L+4XpeiODYnMSCjyKvwQLQgw/fWShJZEA86w7kQHQCUkwFPpoD
DTggepvuK0NeSWQ+EIGZX4PxA7MIbBhTaqd2YC/ebucXW/U0DX0WM3b0M8yr8jq+cAozXVo/bfpB
IEPptd5T5HbKrk9IrFQCatnmx4OMyUbuRGUKd1/G1sqisLnQ2Imb9014rKXV/VBiVJvtm8QBcizu
TVi84z7+EzpS52WKfOJ3quxIwbb+WVCf/6A/stMmvFaywsn/Ia/PmO7TGWyqQ1X2tG9bBoiMAkWa
jcrYe+yALIioZJ5Bavj1OHQ+ZcnQXtAPsl4CoP+C56gWcR+T4a8lmviCNoPObXmqK1IzLS0NbXMa
gD6RRgJw5yzqiO1qrJUU0Ddkuxu1r3SWIC3PaMyWopBPSTeVTQDP3f3oV6edR/yCZ+6x+Pt5JVKp
VZApj1q+4PUUpgzkK7MK1r28aTcqGEyiVY6A21dWmuQWUTDkUGkYeM9+YK900Papy28ZxabCkepF
JVXmHBE7xOBGjkLzaAUDZ/L2uZc+aHIOmxwbkDbsIlTz20gFWSfMJKkB4zhbn3zUnWCXO4ZpqRlP
EF/dy25F8QyIA7P8ZQKTkOF86F7mV5TRCWoToU/xGgQjlaONIwQIHJxP1msiDP5lVtGswcdxH3mZ
ZmwzSFF9sraN2r6Okc6c4FCXww4flkJ/SSWuiF0bafA5uSuoVmtCOnHXEmJBor1t/8wmvEY4mh/B
nUaSEk6HReCWn3ovL/E2lQv1LVFO3VC2076ES7B3wXECg2L8RzgzNQIcARmuuiJu7dh6kauSHtaC
rMlNJXSlaSnM6cghs7hxTZblcff6o+EHEkV7wdl7h5AwEg5wN75DiSwKnp6XnOHcRscUD4kckQrJ
QJk+ADmpWsCPQYV97BEm4Rh2cx0Fw/5WKcXz/kvCTfgekf420WlYsGeOE8/sFp/JcrxvaabFSHDM
9WMOsb4MmYmn4qZnZ1DYTLJ1vbyP/CMjnMg7X30xSvpk0XVoXpANBF2r7GQOLVvCpgYzrvEFluAp
KqKN8UNUlrLCteyTxhYk+iu5ilZFiBpHEVGO0XVduU9VDSLYW0PPqXswtUnWwnfdVoYdAP7D+c4i
UtmKATI8vbNBAmyLWVj8J30PeH8Y8cc4jeSis6uDK3Fdi/zxkg3cg2rt2cuM7w36rwfyo6OFIHN1
x0Kk4uC+flHnnDPodrvcU0ulwpTI35u7Zc2h/aPQwBMtiMa1JBMShMf3cR+T3FY17uon4NxfGUlh
K/1w483Yge9/Mbly0rEGeRt9h/Y8t8G9i50AXESYO2iNo+z3vfJZgCqFQnENvRkc5dRsph2rcGXh
ZLzPo/QqlBW+MVWtIm+6LqZQQe3hrfpZOsm55cIqh3ZKP6tNjXLs0bBmPS3MXPg2PYJiUvWBj8hO
4xfLXTDEaDPPF6lOSRdRbDh2aIb3PYnJdXfFZWls5lSKtUNyG1PsCU7KmjSvLZSrPv5NW+oQJq6Q
MSgJiVVF0v8CnbLiiRtf7GsgtsZQFhqaChYjnNCCjosnFjVauXoH54U29vgPpMdXRnig8EbL+dzG
QAyOtqDpqt9WcxhrWtEv49sex2Zg8J92qHV8J1iCu9LkVVrLM4F9Xs8f4lia4PE0u84OL9gKLNw/
mQuqRs5HRkHmsClAk2EUmfYPuMIMvJwLPGjdN8R83Pms4azqf8ISrFC4TD44PhAAoNYSfcOEBC+b
e9OTgpsb33/ctI+tqR1kBZbuCTmD0gvO1iWn9G6gtp9keXn9CktlWqUvL4IxVya3GIO+vBe6aPSC
62pdHx3+qw+bQla5fts72ZspSM0H1KuT1kVjN9T7CQ6zLnniqwLgsMEWG6GrLzGAoAxOokkDFA4v
kVTGXOaTJLP9Y1SSSpkFHDiCP5NBWoEoRDwdB7FlKPGiSteri35l8qka8bbfp+dpBreh2BizlLXN
EN7whAPmlLJn2FaiN4H0uOxjdmv3I/GZXdGmxgUKZJE0AU9H0MD/3lJvALsVuoymERarsaqHfHyv
9eLI74HYWJFnlu/i/MAQRe9c3znDbUuupYhOHFsJpbHjvj0EHuys96TBGHIUFTWJmxsprom7iRI+
ASWw7CE1Seuk8C/8M1U82xTU6j6AXWN+V7Kg+8vwuDIbfS6xzjKcWLcbG5jlflNYRHG7CS+UeWUo
rAkdoHcOLkdXkxVDQY3uuHx9EwHS8lPJPr9WnjPTDP/ZNuOCEWJQxgpp6D8LDMIxAtev8k7idEVr
cdBvBVm/tuuDefJCoicpAY1o2COnOjqMeHZOeUlT57N7RkC5Dub+g6vY6ExTLcptYymmlYeq9YL/
G57RCuRsmijztMkgWMrta954kJwZcuEgN2pQHZf6sjnyqyFhurX8nHWkPb81I0dEqXvyqhd+Y5lt
+paN2JjLjIKKS0csQ70yViQw7b0aojTGfZ4xCTnp/Z4LF0NakNfJbAZYgmreHkYS1XQseVsQOJ5V
tFwdqUOHHadnZq/eYz+z0Gqc6aUKmZo837aS/Hj8YJoXRbbPNfokQUxuucH2YMahnanu+x5dKPea
mEYqjGDaJvFdhFs9XiX9xBFaM6pB0HEKrfN4Rm4L35Mcd3kGy2fuR92sjlbRSjPCCz5h1B83/xp6
hkMrZR24JlpsOX/j1a/l6KATtOwwGRLAJ5v44oL5PJ3K/kkJ7vZQOILC3SYyqxcoGD0Rs/QKE9FT
MyXK9wCqv3t8veJAofRlEkVLkpP61i5M8/HDCEZ+Uh+1OZUcggTlUTks9qnyvUdxP86BOR4HQWjl
0/LTJ0pF2sn452htPCa1t86pkGB0S4Uf4zrcdZ1LfNW35fn0Oz0kCWixbLqqd7I4yBMw68JSfIp0
Rq6Re3LJvSCJ+BBhokbSf+upyP9xCbZqnY1Wb5D8ioatt09hixN47IDISpiR9QgAApGDJlwUa3C6
bY57STwiLGkAXIyv6aHb+kpVrxhF3rs9mZc3yEAAMMjLZAETHgpMfd45p+QOaLbpaGK2bI2BdO4e
1jqfFc89MBuIPl6SXcLZlc3lYDdti6nMiOVrN4M3o2Uj7NNyr+biIqkbty5Dq0BD90RZ1jJa8MUn
BRe8GRLjx4PVaAxKBDZCsoQzKaZJrAuw48rQDWhLVVFcijvDBQ6ndJ2kl+FRkhHeDFYNN0KafR+0
yWRmFnkZpZ9Jenc1eLzrtZfzjXyEYBFJ19MiqrxkXMddJLFweAC2LhWjA5zQv9KLjY/SEG4Pr7Em
yxnxCOQPJb757n8Sq9WdIN7FD9nzmDQcYTSS2gTVSY2+63JWwSFJOUuPBbrnkytISy00qGbch2NE
CTJAR5/P13T/u7HLeYxxDpopSdjjvlKV9vF3i5XyjZQIwod81bsn7ovyJUNr2kRWnyFAikA9D4tE
FUMwAEDv8+hbPwcnGpl+I4hR40iPesx9Z2T4SbEdsWxW+kJKiV2zoBnlaSzV7oo6wEFaHEgBYwod
qx2Xq59PZnTzgGJMkhIqeAb80q0mIu3pHcJn7mrrdiCKZcsiE8KSNdfXhs6nGnP5+Y0PL1z6DwBg
UqBIErV93mBo9+ykPx0C1+1cRk5lia09QHuRslgOP4fHCTnhpu7biD2OJZdDd2OLyuDVcoL1fRl2
ccjUlzusXhUYQUP+ONGj2y1Wu8+ckGH+6EkzHjNRo/XnvFyI0ooH0OJnUDG3B9BKnTfW2Xi0Po4+
YfhcD7Bvs2KaDzJBq/luIggx/7c5qcanBz2cWN9jyyCiAQa6M8vEg8BYv5uiky/c67k89dCwwQs/
DGfakFAgMuZwmjMzGBsQKZOJx/9/9o4c1V1jbXAjzoA0QDJhk865ZQ/HSzLcP5X+wK1s380hyjE1
nxjQEpnHiiPLzbrki1j7iUKNtHJYkE6RAUWJZKFHuSGrcNYQAsoTd93pRFLvW8JB+IRCVe6T0bKa
48ERKnPt1D1z8T5vFgETgCyoJafNKFPQUIRVUOcGdrjl71ApKTRIHnSInSgKLtWR/6p/mDlFQG3z
EgRQEiBx3r8Fb8uGqyqcg0TatpxPYw/+Y8+kTLZltmcfhwD07oxTp/96MQCiczQ6/LupP2BSkgdH
eCUN/Mjeb1vjL9LtNx/Vtr9LLZb556iB0S7MDVo5/1K0eKRaJOuCfIWtJa2FCyrYc5BRqgAOKrHD
ozBJ5QygcIFHpnC9KBV3r6y2MoMZHiOKSJjI7qDjwmKF04JS8stUKrFoJsJyuXeXh5MyaXJ9DqOv
/eNDIThPu8ijnBnhNBZAN8z4Tz///8PzXZCQL57wkwfzoSseSBithxCNwc9ToAjGUCvqOe/8qeO8
EygXhtO3px4kfLQraB+zYO11e+yvaxEHtilPn0QYvAR17vmz4bw/zk+NhuVKFQhveyYewaIAyv4T
1SeoPZDtME2ZnpEDBecjiXitTG7q4Eeafzixx8RFhfFuzUcSlbNKsgn5ocM/N52OxmmMaMxANwIe
5uLWo7jfy3ONVHqgSNhMH4ToXVY4kianBVo7wgiln6e/HQqqS+O0cLxH0BA56aJ7YG3m+2UKD/hA
Xho1+wy6o84wMTBveS3yGMaeaV5DCliiSm7KslY7F/KODxvF2O1b8cHkIJw/dn7nQ1FftQqp/B/i
dBsqn/hGAl1OvQorbxQGOck5LxfAvnZQZypVZ4KFIZpLhG2rkzmn4GYjtxW7RZRWQ84dfX9AVXQW
X7h3A79UOzXirGkYzDxSI0Z32hIcGdGS+wyM7sFkXKEA4x9X5TxnzVSWZ0Tu0pXgnJ5uME8uqDGI
uz1DZPnMVhUX7ci00CaKhZgCglQeaKjsAIAu0uovI/lIeP0ONCrkJhi7v49I35t5xct4hT2K+jyv
5I768FioavGmkcrrqRnvfeytQKDltygRPVejjvJWNlpyCNgsvh8kOgcPKiYs3qrS6Evb0jt21f3D
4dlEx6RaM3MHnuQ+LnXZo5SIJnecBlfja+YfYh2KnUv2/mLQFa+Rx+FwQCmeHiphEBojblHZbXIq
aPS2T82Rya/o15eHFMukuNtE7hvW05i3kCZrf/I12h4DA1qPphSP9xHZBzH0LcIAxPrinbQP3pL7
XogCBjBtZ66jsMnii9Ilz7pxeE7ahAAUV7C37XWinOmDM5M5fSKK/wTOaswT6vfN7iWCkcJjw7EW
QJCoAunUiO4Q895fiCmLCkLCDAicLD6C5A9zSEtY6ilRNHE1/Hol08JIe5+OTzecS9b3pmUvjlIr
G04e1Fz456X/YYGX3JcNyVEaaTvxWxu1Pg/Id/4g7+2D/3F6kUuscyvdqhfkafoATVqUpPtiBR7R
SoA9JXzz9aBfYXmqNqC41DDim3/Xb2M2JU9uYj0GV+utXHuILDjLz6CPSYdkNQtHILK2XHEauLYZ
J1mu37HqVslCduLQAy+XVt1bdrhIQimdIIbNowSxNF2W89mKKB+lR2JowvF5hAJElq9oJC5YISqw
JEEZ0EikwbC/6MoBT2evb5VT6CSIt8Q+7S8GoGOHhEXHAZTF3OKw1BR1m0X2FBsDclhr3oZZcAG6
4eWNYyTiPHxumW+XOCylxYOwE7cET6vSvd1DDvoksXXkB/CypSdgMY23nkNOvaFicynFeRzf92Xa
FMAlcFJqibM3qGGpq1Krf2styp/GShSiGWzJjzeiWTDj2G6jZsZy0RhZN1eF0M8kv2X9f3E16nGw
EONMWVEuMl5UKOElf3Na3M2d6IlKMVNa9vZNn9HGQ1LLiPTO/gyT+0yAn2SWOCaDYeJoivsSCYoU
ibPot7wkbCIKHocMfBYYnUy1OmFGTAzUgSGLT8LkCN98T5RsDuuuMc37eutEH0w2yjY9zTkyXKAg
qtuGylBgNV55EtXW4CuutPB5faeBYJswlGJviPTtDJfrS+1UJNTGiL41+JjDDAX51cjyH5kM6e/O
uqVkuDhrk9XAjVMCVUVqhQRfHJgaRvczaiMR6aGir//aJEQ3UBe2HequCcRXL5bOm9+ZpKpui/f1
uw1eGj4DLV4UbGKqzG3n1/SnJ19p+9oOrvXqJMrPHi5ZJsYv2SuaO5CaZ4vxKiAaf1U+mksC6eJ2
UNyPbW5NL8/WCAvM9rZXMYisOyskT4QPyCG9cDbSRDIMpSitaKhsUl4rTbiMMPI7DIPzn5pY8HBS
nI4FWuY2XxRxVl8mbeMZPzbvcO1tmQ15C3+icRVqaKE/Aq+m04O3iSO3MKarRsRulmWzEU7Rpkjv
rcNVVsmfx6rJiCKxW0prpxuYdix15YG37VWPncf7Gytx15Ui1Kl5N6J6VKFxVN4+u1d6uhPqdxbW
HX4Dl1WPn+ltAkTdFIKtC6Z4UyZ4+LdwXD6Jm0MhZWYqV0cc25Z4l9zNvDRwNV4uVCOdFSeryKgT
Gga2MzX6reseifxKQO5bYL+5U9d5ELB7YAbRq3jZU0K1qAzmsDwOFymrr8SjlycOp7Kz62XsZ19f
Qei44ow9QxM3Wxr31UFgTwKE1ooprmWt7MvQhTFC4nCflUxRIRt2RVz87IZnHHdl8JLzGWPkBlG2
HIeOScg0nDW8SDiZaBrq+gDM50+ZTG0EUPfWthyysbRtnWJR0pXOmlDsa8lnNcI0Jdyf9YEcsZcd
Nyk/a4X2LdyqqW39Po8ghKqkueU+x+qHZRD9Ez9yP2kAI4FXLQzf/gN/VP8WQDS9Pwy/GgJc/yrI
UIPn4eWd2T0jPhxQzQD6Oxxk+GhhF+uEA3X7l8WtYjsoAn+NdyvFkvMwP4jJgbT6xyjMaU6yl8Nf
uI4/IiHIZT+bEYFZzPD33j3Xu8VDO+1p3tDGjeK7bR5KIipmdUio9aRISXZtvYnqz1+0WX2GwgDz
+Uf9gbp56d5tXDMC2oWbWWQn5XLJTSfW1oa/Xw6vDGippTCis72wSiwrV68cwJQUrmm1YZzcgmdD
W40O7u8/NVzRYvyrqHgMHSmbTu2L10an+Fr7HpDBsHXeBtvBnzrdkSbTSe/0b+0o09xfrSBaMey1
WRfj9XBlF3FvQyisyZ06IhRJLkqSDvL0SEZP82AQ/QYGaT7ptD3sNPug7Uc2PgGeMUxblr64dzdd
VcYkAsgEyS2pFNp65ngI0jzvLanrY6Fcm5tuEZo7pl4BFIoCrIym23LNbxNBTPNhKv+Y0RzYX7AA
Wzd5J2tgansPvOTCLjAoWaIkGJllBaAyJ9QiMwXoesu2o74hyorOntoVZGlLSP0YyyGIXYXmdcEy
qRT3mEe6PfN0UrjFP6RiY7dCzq2fuiV9HY8QaYOw+68bc9vQNe3+jtrdyq1jFcmrhvU+SBgSZOTG
u0NimxRivBKUQTjV2hDMTW6wGnFS5qnwj9jPicrhsA3DocugmcVpFcKAEuj1+l2Ulr6SnNnWVTLs
qFEWbRhJ5oMCAgOOb4XpKpk8qLfy161BKho9harK/qiOGLyiAnv20LY70dSKvM9vzYv6Lvkon4qa
nZ6XzE1AtSQ4weAthaV1Ky29vILL+2xZ9FOIOGU0jNcfWJ6D9gceBBtKfvV6ltR+6xs7xFq+5vmt
AAWxWGHWGM4Jyaeqlz54fiaBvauX8/aNedL5QsxSgb08DWu96nT5hwCWErLG6z1NY9yMPt/3VI7z
1k5HAIqyPFjo5WW2LRTTH568UQjCsnFEgvftGtlXz9dyhjsWFUOrg7SSYF2Mgm93nmFd94Nvic/z
+lEt5nFL3wLbpRliRXkjueElVQ7Ml+iOc6WqxGP9BQyAaIYTB66aaWskrRPSlbIFVVtu9rkMszpr
SdyficyOXUCIDzQd4FcfD6GRZoTCEtNO7GnAbRkqOv4+VUB8yKtzqgPN/CBnYLnR396OE4Jncmzp
WS9gmq9HQ30bN4HKEuq3ZZv2JNDoRTSSgd5GvYLgbVT7OxaRbJ3snC/sBtcB+h7GEnlOtmd0Kt5q
5ZLRb9Q1UAv4mi0cYVlTelAeqX7pQ0VgZmRtshpLkW/0DHuqpQ9RRdOXsg23D6GZKO9PtcaMofjv
Wu2W2Br3GRFGWAvW79tHYmEvQXDOsrNjnGNDEFKRTTDyjRHslZDz8H3QEHW4FJfxWo9zyA3xzdds
PDmDYh1caAfmHCVGWWh2HaJ5XJymBhbTqyBB70X+fNoHBMWoDkNNtYEwPveNVjFbe1s3L/cZ/0OQ
mt1/iTWDym4kMLzpy/hXeu6aHaVqSZh+mxsUhI4jT1H8yMp10llxpmqphXUnx0XfAj+kot76l46u
w5NS5REHBg9xlVVJ1wM+YAsylB252SWCiNDxOJ/G1K7skw7OG37TQI4yBP3pm7iSrdNPkmUc5l5P
wEzaPobj9CcGpA/UKmEHCzrAF34fKnw9o3yfZjuVRo2Nn6FfV97zyOQxYRzJox43PfvxE7JxvNeM
gtyQ85XiU6XkfFM6Q2aW7nDINb8D2z+z+MpjgGyTbL9HXZLSA6Cj6yrRhG4jhtv206ItL33ALXrH
ca1ZxEabkvqOSzNilbCRacsCzWSHrTx0cJpGb/wFFwOrSZoSOOi90RidQioWPRTv2X7j/sFI6vSN
YkldGzS+lCNVGfJXts1wXkOv11HzWX6fsJsgDV1sz2Bx9JQcQe2FaxnrneAONdHjG9/d4BCFYHGy
PoOsBzO8CZB8mkFWLTujxOEN88b1eXVA9uLQ3z1iH20IaVzwcrJH8jK8LcEBgnyS8T4KOKgKJKPQ
XqHr1Gv+6ppfwdkF/rlfuNQPJb4ryx3aDyhqs8fECka18RNLi16QMaUlg3ntjXc5YpoIiy+hm7Yz
yoMOqmkmUv6PGbhZ4wTvPzTAnoGDj3l1pf59yL3GnQa3TWcJzvSjG9aePGQ6NcNgKb9JiVL6uwCj
bmgz/gZI3iTlqutymwP4pVQoG77Pt5IQtRIq5iTk7ZqvJnft6aRPw1aT0hLzMcAHu8u0tmizQd6B
L+2DvI09nDo18PqMm++UZm4aU+Z51/G2PfntTD9aOJbMxbwDDhUKsbdkiNfT3rRJQN/3Oc6tvvF0
ALkLDzUADYouspcVPO1H+q43UPuBN97Efigt0y96Qcu9oBjCM50SGKqzxzVSwTRJ4eCvymjLvVaD
MPJCBoKgXsuC44qc46g+4LC/wzDF1Cmn7SGMGpfxaP/lyDbE9sADEWorZL6aJxHwnYj/Hy2F36AT
Y+/ekcNLNvWXfFGilo9G0gk/2+HqOwd5GYKxyiPIwj99QvKOq1JGqGClp4VUmkrehTNwiLsYYCP+
Wyr7QMqCBhB0r3H6iZbeAaCjuOLcCTSfAeo3O7w9XV5jy9yQ3Z8TjxSZ9NuRMocE0mi3PV2lBiJy
K43cQmRSAbwkPXAbcdaL4cibwpiWayp20zvMotZi28jm/Mt2JXxsPh7GfEsVX8Hu5s9hHz3OcERJ
nQegQu4VUN5caHiSM4CAd0/pBbA9Os7kgAONEelmmlDDifF0TGbssQ7eEUeFgRL6i1yduF7gJYsE
ZqyFV19BSIGj321E14x3CUcUCgWsHb0zmcsSNMbRJcHIB+8o07xfGNG4x3/cl9tSx2DYYwTn5t31
s2J0q93hAYyuCRPhLxRlu6xeXDTPV6FtsCUc4bdd4eoeA1lMVZPKDSjXqC5fIZVCEGhodVZVEmjg
JfbXyIzB1s7q38PQ+ORlNp56RmODqQUvCbAO64TEKzOPcDthn4YB3bB+mpyJJknkRz3V5OvBJiCm
ulZXbQnsonwZODc8QmijGvqXwhdCYiV2Abioxe1Ffr+MMbGEZyh5eblGBelqUlGGTeVIc0a5CHdm
DFBPkXEZcsyII3N4AVOOz1A=
`protect end_protected

